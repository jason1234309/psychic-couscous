module top(
  input LIOB33_SING_X0Y0_IOB_X0Y0_IPAD,
  input LIOB33_SING_X0Y149_IOB_X0Y149_IPAD,
  input LIOB33_SING_X0Y150_IOB_X0Y150_IPAD,
  input LIOB33_SING_X0Y199_IOB_X0Y199_IPAD,
  input LIOB33_SING_X0Y200_IOB_X0Y200_IPAD,
  input LIOB33_SING_X0Y249_IOB_X0Y249_IPAD,
  input LIOB33_SING_X0Y50_IOB_X0Y50_IPAD,
  input LIOB33_SING_X0Y99_IOB_X0Y99_IPAD,
  input LIOB33_X0Y101_IOB_X0Y101_IPAD,
  input LIOB33_X0Y101_IOB_X0Y102_IPAD,
  input LIOB33_X0Y103_IOB_X0Y103_IPAD,
  input LIOB33_X0Y103_IOB_X0Y104_IPAD,
  input LIOB33_X0Y105_IOB_X0Y105_IPAD,
  input LIOB33_X0Y105_IOB_X0Y106_IPAD,
  input LIOB33_X0Y107_IOB_X0Y107_IPAD,
  input LIOB33_X0Y107_IOB_X0Y108_IPAD,
  input LIOB33_X0Y109_IOB_X0Y109_IPAD,
  input LIOB33_X0Y109_IOB_X0Y110_IPAD,
  input LIOB33_X0Y111_IOB_X0Y111_IPAD,
  input LIOB33_X0Y111_IOB_X0Y112_IPAD,
  input LIOB33_X0Y113_IOB_X0Y113_IPAD,
  input LIOB33_X0Y113_IOB_X0Y114_IPAD,
  input LIOB33_X0Y115_IOB_X0Y115_IPAD,
  input LIOB33_X0Y115_IOB_X0Y116_IPAD,
  input LIOB33_X0Y117_IOB_X0Y117_IPAD,
  input LIOB33_X0Y117_IOB_X0Y118_IPAD,
  input LIOB33_X0Y119_IOB_X0Y119_IPAD,
  input LIOB33_X0Y119_IOB_X0Y120_IPAD,
  input LIOB33_X0Y11_IOB_X0Y11_IPAD,
  input LIOB33_X0Y11_IOB_X0Y12_IPAD,
  input LIOB33_X0Y121_IOB_X0Y121_IPAD,
  input LIOB33_X0Y121_IOB_X0Y122_IPAD,
  input LIOB33_X0Y123_IOB_X0Y123_IPAD,
  input LIOB33_X0Y123_IOB_X0Y124_IPAD,
  input LIOB33_X0Y125_IOB_X0Y125_IPAD,
  input LIOB33_X0Y125_IOB_X0Y126_IPAD,
  input LIOB33_X0Y127_IOB_X0Y127_IPAD,
  input LIOB33_X0Y127_IOB_X0Y128_IPAD,
  input LIOB33_X0Y129_IOB_X0Y129_IPAD,
  input LIOB33_X0Y129_IOB_X0Y130_IPAD,
  input LIOB33_X0Y131_IOB_X0Y131_IPAD,
  input LIOB33_X0Y131_IOB_X0Y132_IPAD,
  input LIOB33_X0Y133_IOB_X0Y133_IPAD,
  input LIOB33_X0Y133_IOB_X0Y134_IPAD,
  input LIOB33_X0Y135_IOB_X0Y135_IPAD,
  input LIOB33_X0Y135_IOB_X0Y136_IPAD,
  input LIOB33_X0Y137_IOB_X0Y137_IPAD,
  input LIOB33_X0Y137_IOB_X0Y138_IPAD,
  input LIOB33_X0Y139_IOB_X0Y139_IPAD,
  input LIOB33_X0Y139_IOB_X0Y140_IPAD,
  input LIOB33_X0Y13_IOB_X0Y13_IPAD,
  input LIOB33_X0Y13_IOB_X0Y14_IPAD,
  input LIOB33_X0Y141_IOB_X0Y141_IPAD,
  input LIOB33_X0Y141_IOB_X0Y142_IPAD,
  input LIOB33_X0Y143_IOB_X0Y143_IPAD,
  input LIOB33_X0Y145_IOB_X0Y145_IPAD,
  input LIOB33_X0Y145_IOB_X0Y146_IPAD,
  input LIOB33_X0Y147_IOB_X0Y147_IPAD,
  input LIOB33_X0Y147_IOB_X0Y148_IPAD,
  input LIOB33_X0Y151_IOB_X0Y151_IPAD,
  input LIOB33_X0Y151_IOB_X0Y152_IPAD,
  input LIOB33_X0Y153_IOB_X0Y153_IPAD,
  input LIOB33_X0Y153_IOB_X0Y154_IPAD,
  input LIOB33_X0Y155_IOB_X0Y155_IPAD,
  input LIOB33_X0Y155_IOB_X0Y156_IPAD,
  input LIOB33_X0Y157_IOB_X0Y157_IPAD,
  input LIOB33_X0Y157_IOB_X0Y158_IPAD,
  input LIOB33_X0Y159_IOB_X0Y159_IPAD,
  input LIOB33_X0Y159_IOB_X0Y160_IPAD,
  input LIOB33_X0Y15_IOB_X0Y15_IPAD,
  input LIOB33_X0Y15_IOB_X0Y16_IPAD,
  input LIOB33_X0Y161_IOB_X0Y161_IPAD,
  input LIOB33_X0Y161_IOB_X0Y162_IPAD,
  input LIOB33_X0Y163_IOB_X0Y163_IPAD,
  input LIOB33_X0Y163_IOB_X0Y164_IPAD,
  input LIOB33_X0Y165_IOB_X0Y165_IPAD,
  input LIOB33_X0Y165_IOB_X0Y166_IPAD,
  input LIOB33_X0Y167_IOB_X0Y167_IPAD,
  input LIOB33_X0Y167_IOB_X0Y168_IPAD,
  input LIOB33_X0Y169_IOB_X0Y169_IPAD,
  input LIOB33_X0Y169_IOB_X0Y170_IPAD,
  input LIOB33_X0Y171_IOB_X0Y171_IPAD,
  input LIOB33_X0Y171_IOB_X0Y172_IPAD,
  input LIOB33_X0Y173_IOB_X0Y173_IPAD,
  input LIOB33_X0Y173_IOB_X0Y174_IPAD,
  input LIOB33_X0Y175_IOB_X0Y175_IPAD,
  input LIOB33_X0Y175_IOB_X0Y176_IPAD,
  input LIOB33_X0Y177_IOB_X0Y177_IPAD,
  input LIOB33_X0Y177_IOB_X0Y178_IPAD,
  input LIOB33_X0Y179_IOB_X0Y179_IPAD,
  input LIOB33_X0Y179_IOB_X0Y180_IPAD,
  input LIOB33_X0Y17_IOB_X0Y17_IPAD,
  input LIOB33_X0Y17_IOB_X0Y18_IPAD,
  input LIOB33_X0Y181_IOB_X0Y181_IPAD,
  input LIOB33_X0Y181_IOB_X0Y182_IPAD,
  input LIOB33_X0Y183_IOB_X0Y183_IPAD,
  input LIOB33_X0Y183_IOB_X0Y184_IPAD,
  input LIOB33_X0Y185_IOB_X0Y185_IPAD,
  input LIOB33_X0Y185_IOB_X0Y186_IPAD,
  input LIOB33_X0Y187_IOB_X0Y187_IPAD,
  input LIOB33_X0Y187_IOB_X0Y188_IPAD,
  input LIOB33_X0Y189_IOB_X0Y189_IPAD,
  input LIOB33_X0Y189_IOB_X0Y190_IPAD,
  input LIOB33_X0Y191_IOB_X0Y191_IPAD,
  input LIOB33_X0Y191_IOB_X0Y192_IPAD,
  input LIOB33_X0Y193_IOB_X0Y193_IPAD,
  input LIOB33_X0Y193_IOB_X0Y194_IPAD,
  input LIOB33_X0Y195_IOB_X0Y195_IPAD,
  input LIOB33_X0Y195_IOB_X0Y196_IPAD,
  input LIOB33_X0Y197_IOB_X0Y197_IPAD,
  input LIOB33_X0Y197_IOB_X0Y198_IPAD,
  input LIOB33_X0Y19_IOB_X0Y19_IPAD,
  input LIOB33_X0Y19_IOB_X0Y20_IPAD,
  input LIOB33_X0Y1_IOB_X0Y1_IPAD,
  input LIOB33_X0Y1_IOB_X0Y2_IPAD,
  input LIOB33_X0Y201_IOB_X0Y201_IPAD,
  input LIOB33_X0Y201_IOB_X0Y202_IPAD,
  input LIOB33_X0Y203_IOB_X0Y203_IPAD,
  input LIOB33_X0Y203_IOB_X0Y204_IPAD,
  input LIOB33_X0Y205_IOB_X0Y205_IPAD,
  input LIOB33_X0Y205_IOB_X0Y206_IPAD,
  input LIOB33_X0Y207_IOB_X0Y207_IPAD,
  input LIOB33_X0Y207_IOB_X0Y208_IPAD,
  input LIOB33_X0Y209_IOB_X0Y209_IPAD,
  input LIOB33_X0Y209_IOB_X0Y210_IPAD,
  input LIOB33_X0Y211_IOB_X0Y211_IPAD,
  input LIOB33_X0Y211_IOB_X0Y212_IPAD,
  input LIOB33_X0Y213_IOB_X0Y213_IPAD,
  input LIOB33_X0Y213_IOB_X0Y214_IPAD,
  input LIOB33_X0Y215_IOB_X0Y215_IPAD,
  input LIOB33_X0Y215_IOB_X0Y216_IPAD,
  input LIOB33_X0Y217_IOB_X0Y217_IPAD,
  input LIOB33_X0Y217_IOB_X0Y218_IPAD,
  input LIOB33_X0Y219_IOB_X0Y219_IPAD,
  input LIOB33_X0Y219_IOB_X0Y220_IPAD,
  input LIOB33_X0Y21_IOB_X0Y21_IPAD,
  input LIOB33_X0Y21_IOB_X0Y22_IPAD,
  input LIOB33_X0Y221_IOB_X0Y221_IPAD,
  input LIOB33_X0Y221_IOB_X0Y222_IPAD,
  input LIOB33_X0Y223_IOB_X0Y223_IPAD,
  input LIOB33_X0Y223_IOB_X0Y224_IPAD,
  input LIOB33_X0Y225_IOB_X0Y225_IPAD,
  input LIOB33_X0Y225_IOB_X0Y226_IPAD,
  input LIOB33_X0Y227_IOB_X0Y227_IPAD,
  input LIOB33_X0Y227_IOB_X0Y228_IPAD,
  input LIOB33_X0Y229_IOB_X0Y229_IPAD,
  input LIOB33_X0Y229_IOB_X0Y230_IPAD,
  input LIOB33_X0Y231_IOB_X0Y231_IPAD,
  input LIOB33_X0Y231_IOB_X0Y232_IPAD,
  input LIOB33_X0Y233_IOB_X0Y233_IPAD,
  input LIOB33_X0Y233_IOB_X0Y234_IPAD,
  input LIOB33_X0Y235_IOB_X0Y235_IPAD,
  input LIOB33_X0Y235_IOB_X0Y236_IPAD,
  input LIOB33_X0Y237_IOB_X0Y237_IPAD,
  input LIOB33_X0Y237_IOB_X0Y238_IPAD,
  input LIOB33_X0Y239_IOB_X0Y239_IPAD,
  input LIOB33_X0Y239_IOB_X0Y240_IPAD,
  input LIOB33_X0Y23_IOB_X0Y23_IPAD,
  input LIOB33_X0Y23_IOB_X0Y24_IPAD,
  input LIOB33_X0Y241_IOB_X0Y241_IPAD,
  input LIOB33_X0Y241_IOB_X0Y242_IPAD,
  input LIOB33_X0Y243_IOB_X0Y243_IPAD,
  input LIOB33_X0Y243_IOB_X0Y244_IPAD,
  input LIOB33_X0Y245_IOB_X0Y245_IPAD,
  input LIOB33_X0Y245_IOB_X0Y246_IPAD,
  input LIOB33_X0Y247_IOB_X0Y247_IPAD,
  input LIOB33_X0Y247_IOB_X0Y248_IPAD,
  input LIOB33_X0Y25_IOB_X0Y25_IPAD,
  input LIOB33_X0Y25_IOB_X0Y26_IPAD,
  input LIOB33_X0Y27_IOB_X0Y27_IPAD,
  input LIOB33_X0Y27_IOB_X0Y28_IPAD,
  input LIOB33_X0Y29_IOB_X0Y29_IPAD,
  input LIOB33_X0Y29_IOB_X0Y30_IPAD,
  input LIOB33_X0Y31_IOB_X0Y31_IPAD,
  input LIOB33_X0Y3_IOB_X0Y3_IPAD,
  input LIOB33_X0Y3_IOB_X0Y4_IPAD,
  input LIOB33_X0Y51_IOB_X0Y51_IPAD,
  input LIOB33_X0Y51_IOB_X0Y52_IPAD,
  input LIOB33_X0Y53_IOB_X0Y53_IPAD,
  input LIOB33_X0Y53_IOB_X0Y54_IPAD,
  input LIOB33_X0Y55_IOB_X0Y55_IPAD,
  input LIOB33_X0Y55_IOB_X0Y56_IPAD,
  input LIOB33_X0Y57_IOB_X0Y57_IPAD,
  input LIOB33_X0Y57_IOB_X0Y58_IPAD,
  input LIOB33_X0Y59_IOB_X0Y59_IPAD,
  input LIOB33_X0Y59_IOB_X0Y60_IPAD,
  input LIOB33_X0Y5_IOB_X0Y5_IPAD,
  input LIOB33_X0Y5_IOB_X0Y6_IPAD,
  input LIOB33_X0Y61_IOB_X0Y61_IPAD,
  input LIOB33_X0Y61_IOB_X0Y62_IPAD,
  input LIOB33_X0Y63_IOB_X0Y63_IPAD,
  input LIOB33_X0Y63_IOB_X0Y64_IPAD,
  input LIOB33_X0Y65_IOB_X0Y65_IPAD,
  input LIOB33_X0Y65_IOB_X0Y66_IPAD,
  input LIOB33_X0Y67_IOB_X0Y67_IPAD,
  input LIOB33_X0Y67_IOB_X0Y68_IPAD,
  input LIOB33_X0Y69_IOB_X0Y69_IPAD,
  input LIOB33_X0Y69_IOB_X0Y70_IPAD,
  input LIOB33_X0Y71_IOB_X0Y71_IPAD,
  input LIOB33_X0Y71_IOB_X0Y72_IPAD,
  input LIOB33_X0Y73_IOB_X0Y73_IPAD,
  input LIOB33_X0Y73_IOB_X0Y74_IPAD,
  input LIOB33_X0Y75_IOB_X0Y75_IPAD,
  input LIOB33_X0Y75_IOB_X0Y76_IPAD,
  input LIOB33_X0Y77_IOB_X0Y77_IPAD,
  input LIOB33_X0Y77_IOB_X0Y78_IPAD,
  input LIOB33_X0Y79_IOB_X0Y79_IPAD,
  input LIOB33_X0Y79_IOB_X0Y80_IPAD,
  input LIOB33_X0Y7_IOB_X0Y7_IPAD,
  input LIOB33_X0Y7_IOB_X0Y8_IPAD,
  input LIOB33_X0Y81_IOB_X0Y81_IPAD,
  input LIOB33_X0Y81_IOB_X0Y82_IPAD,
  input LIOB33_X0Y83_IOB_X0Y83_IPAD,
  input LIOB33_X0Y83_IOB_X0Y84_IPAD,
  input LIOB33_X0Y85_IOB_X0Y85_IPAD,
  input LIOB33_X0Y85_IOB_X0Y86_IPAD,
  input LIOB33_X0Y87_IOB_X0Y87_IPAD,
  input LIOB33_X0Y87_IOB_X0Y88_IPAD,
  input LIOB33_X0Y89_IOB_X0Y89_IPAD,
  input LIOB33_X0Y89_IOB_X0Y90_IPAD,
  input LIOB33_X0Y91_IOB_X0Y91_IPAD,
  input LIOB33_X0Y91_IOB_X0Y92_IPAD,
  input LIOB33_X0Y93_IOB_X0Y93_IPAD,
  input LIOB33_X0Y93_IOB_X0Y94_IPAD,
  input LIOB33_X0Y95_IOB_X0Y95_IPAD,
  input LIOB33_X0Y95_IOB_X0Y96_IPAD,
  input LIOB33_X0Y97_IOB_X0Y97_IPAD,
  input LIOB33_X0Y97_IOB_X0Y98_IPAD,
  input LIOB33_X0Y9_IOB_X0Y10_IPAD,
  input LIOB33_X0Y9_IOB_X0Y9_IPAD,
  input RIOB33_SING_X105Y199_IOB_X1Y199_IPAD,
  input RIOB33_SING_X105Y200_IOB_X1Y200_IPAD,
  input RIOB33_X105Y177_IOB_X1Y178_IPAD,
  input RIOB33_X105Y179_IOB_X1Y179_IPAD,
  input RIOB33_X105Y179_IOB_X1Y180_IPAD,
  input RIOB33_X105Y181_IOB_X1Y181_IPAD,
  input RIOB33_X105Y181_IOB_X1Y182_IPAD,
  input RIOB33_X105Y183_IOB_X1Y183_IPAD,
  input RIOB33_X105Y183_IOB_X1Y184_IPAD,
  input RIOB33_X105Y185_IOB_X1Y185_IPAD,
  input RIOB33_X105Y185_IOB_X1Y186_IPAD,
  input RIOB33_X105Y187_IOB_X1Y187_IPAD,
  input RIOB33_X105Y187_IOB_X1Y188_IPAD,
  input RIOB33_X105Y189_IOB_X1Y189_IPAD,
  input RIOB33_X105Y189_IOB_X1Y190_IPAD,
  input RIOB33_X105Y191_IOB_X1Y191_IPAD,
  input RIOB33_X105Y191_IOB_X1Y192_IPAD,
  input RIOB33_X105Y193_IOB_X1Y193_IPAD,
  input RIOB33_X105Y193_IOB_X1Y194_IPAD,
  input RIOB33_X105Y195_IOB_X1Y195_IPAD,
  input RIOB33_X105Y195_IOB_X1Y196_IPAD,
  input RIOB33_X105Y197_IOB_X1Y197_IPAD,
  input RIOB33_X105Y197_IOB_X1Y198_IPAD,
  input RIOB33_X105Y201_IOB_X1Y201_IPAD,
  input RIOB33_X105Y201_IOB_X1Y202_IPAD,
  input RIOB33_X105Y203_IOB_X1Y203_IPAD,
  input RIOB33_X105Y203_IOB_X1Y204_IPAD,
  input RIOB33_X105Y205_IOB_X1Y205_IPAD,
  output LIOB33_SING_X0Y100_IOB_X0Y100_OPAD,
  output RIOB33_SING_X105Y100_IOB_X1Y100_OPAD,
  output RIOB33_SING_X105Y149_IOB_X1Y149_OPAD,
  output RIOB33_SING_X105Y150_IOB_X1Y150_OPAD,
  output RIOB33_SING_X105Y50_IOB_X1Y50_OPAD,
  output RIOB33_SING_X105Y99_IOB_X1Y99_OPAD,
  output RIOB33_X105Y101_IOB_X1Y101_OPAD,
  output RIOB33_X105Y101_IOB_X1Y102_OPAD,
  output RIOB33_X105Y103_IOB_X1Y103_OPAD,
  output RIOB33_X105Y103_IOB_X1Y104_OPAD,
  output RIOB33_X105Y105_IOB_X1Y105_OPAD,
  output RIOB33_X105Y105_IOB_X1Y106_OPAD,
  output RIOB33_X105Y107_IOB_X1Y107_OPAD,
  output RIOB33_X105Y107_IOB_X1Y108_OPAD,
  output RIOB33_X105Y109_IOB_X1Y109_OPAD,
  output RIOB33_X105Y109_IOB_X1Y110_OPAD,
  output RIOB33_X105Y111_IOB_X1Y111_OPAD,
  output RIOB33_X105Y111_IOB_X1Y112_OPAD,
  output RIOB33_X105Y113_IOB_X1Y113_OPAD,
  output RIOB33_X105Y113_IOB_X1Y114_OPAD,
  output RIOB33_X105Y115_IOB_X1Y115_OPAD,
  output RIOB33_X105Y115_IOB_X1Y116_OPAD,
  output RIOB33_X105Y117_IOB_X1Y117_OPAD,
  output RIOB33_X105Y117_IOB_X1Y118_OPAD,
  output RIOB33_X105Y119_IOB_X1Y119_OPAD,
  output RIOB33_X105Y119_IOB_X1Y120_OPAD,
  output RIOB33_X105Y121_IOB_X1Y121_OPAD,
  output RIOB33_X105Y121_IOB_X1Y122_OPAD,
  output RIOB33_X105Y123_IOB_X1Y123_OPAD,
  output RIOB33_X105Y123_IOB_X1Y124_OPAD,
  output RIOB33_X105Y125_IOB_X1Y125_OPAD,
  output RIOB33_X105Y125_IOB_X1Y126_OPAD,
  output RIOB33_X105Y127_IOB_X1Y127_OPAD,
  output RIOB33_X105Y127_IOB_X1Y128_OPAD,
  output RIOB33_X105Y129_IOB_X1Y129_OPAD,
  output RIOB33_X105Y129_IOB_X1Y130_OPAD,
  output RIOB33_X105Y131_IOB_X1Y131_OPAD,
  output RIOB33_X105Y131_IOB_X1Y132_OPAD,
  output RIOB33_X105Y133_IOB_X1Y133_OPAD,
  output RIOB33_X105Y133_IOB_X1Y134_OPAD,
  output RIOB33_X105Y135_IOB_X1Y135_OPAD,
  output RIOB33_X105Y135_IOB_X1Y136_OPAD,
  output RIOB33_X105Y137_IOB_X1Y137_OPAD,
  output RIOB33_X105Y137_IOB_X1Y138_OPAD,
  output RIOB33_X105Y139_IOB_X1Y139_OPAD,
  output RIOB33_X105Y139_IOB_X1Y140_OPAD,
  output RIOB33_X105Y141_IOB_X1Y141_OPAD,
  output RIOB33_X105Y141_IOB_X1Y142_OPAD,
  output RIOB33_X105Y143_IOB_X1Y143_OPAD,
  output RIOB33_X105Y143_IOB_X1Y144_OPAD,
  output RIOB33_X105Y145_IOB_X1Y145_OPAD,
  output RIOB33_X105Y145_IOB_X1Y146_OPAD,
  output RIOB33_X105Y147_IOB_X1Y147_OPAD,
  output RIOB33_X105Y147_IOB_X1Y148_OPAD,
  output RIOB33_X105Y151_IOB_X1Y151_OPAD,
  output RIOB33_X105Y151_IOB_X1Y152_OPAD,
  output RIOB33_X105Y153_IOB_X1Y153_OPAD,
  output RIOB33_X105Y153_IOB_X1Y154_OPAD,
  output RIOB33_X105Y155_IOB_X1Y155_OPAD,
  output RIOB33_X105Y155_IOB_X1Y156_OPAD,
  output RIOB33_X105Y157_IOB_X1Y157_OPAD,
  output RIOB33_X105Y157_IOB_X1Y158_OPAD,
  output RIOB33_X105Y159_IOB_X1Y159_OPAD,
  output RIOB33_X105Y159_IOB_X1Y160_OPAD,
  output RIOB33_X105Y161_IOB_X1Y161_OPAD,
  output RIOB33_X105Y161_IOB_X1Y162_OPAD,
  output RIOB33_X105Y163_IOB_X1Y163_OPAD,
  output RIOB33_X105Y163_IOB_X1Y164_OPAD,
  output RIOB33_X105Y165_IOB_X1Y165_OPAD,
  output RIOB33_X105Y165_IOB_X1Y166_OPAD,
  output RIOB33_X105Y167_IOB_X1Y167_OPAD,
  output RIOB33_X105Y167_IOB_X1Y168_OPAD,
  output RIOB33_X105Y169_IOB_X1Y169_OPAD,
  output RIOB33_X105Y169_IOB_X1Y170_OPAD,
  output RIOB33_X105Y171_IOB_X1Y171_OPAD,
  output RIOB33_X105Y171_IOB_X1Y172_OPAD,
  output RIOB33_X105Y173_IOB_X1Y173_OPAD,
  output RIOB33_X105Y173_IOB_X1Y174_OPAD,
  output RIOB33_X105Y175_IOB_X1Y175_OPAD,
  output RIOB33_X105Y175_IOB_X1Y176_OPAD,
  output RIOB33_X105Y177_IOB_X1Y177_OPAD,
  output RIOB33_X105Y51_IOB_X1Y51_OPAD,
  output RIOB33_X105Y51_IOB_X1Y52_OPAD,
  output RIOB33_X105Y53_IOB_X1Y53_OPAD,
  output RIOB33_X105Y53_IOB_X1Y54_OPAD,
  output RIOB33_X105Y55_IOB_X1Y55_OPAD,
  output RIOB33_X105Y55_IOB_X1Y56_OPAD,
  output RIOB33_X105Y57_IOB_X1Y57_OPAD,
  output RIOB33_X105Y57_IOB_X1Y58_OPAD,
  output RIOB33_X105Y59_IOB_X1Y59_OPAD,
  output RIOB33_X105Y59_IOB_X1Y60_OPAD,
  output RIOB33_X105Y61_IOB_X1Y61_OPAD,
  output RIOB33_X105Y61_IOB_X1Y62_OPAD,
  output RIOB33_X105Y63_IOB_X1Y63_OPAD,
  output RIOB33_X105Y63_IOB_X1Y64_OPAD,
  output RIOB33_X105Y65_IOB_X1Y65_OPAD,
  output RIOB33_X105Y65_IOB_X1Y66_OPAD,
  output RIOB33_X105Y67_IOB_X1Y67_OPAD,
  output RIOB33_X105Y67_IOB_X1Y68_OPAD,
  output RIOB33_X105Y69_IOB_X1Y69_OPAD,
  output RIOB33_X105Y69_IOB_X1Y70_OPAD,
  output RIOB33_X105Y71_IOB_X1Y71_OPAD,
  output RIOB33_X105Y71_IOB_X1Y72_OPAD,
  output RIOB33_X105Y73_IOB_X1Y73_OPAD,
  output RIOB33_X105Y73_IOB_X1Y74_OPAD,
  output RIOB33_X105Y75_IOB_X1Y75_OPAD,
  output RIOB33_X105Y75_IOB_X1Y76_OPAD,
  output RIOB33_X105Y77_IOB_X1Y77_OPAD,
  output RIOB33_X105Y77_IOB_X1Y78_OPAD,
  output RIOB33_X105Y79_IOB_X1Y79_OPAD,
  output RIOB33_X105Y79_IOB_X1Y80_OPAD,
  output RIOB33_X105Y81_IOB_X1Y81_OPAD,
  output RIOB33_X105Y81_IOB_X1Y82_OPAD,
  output RIOB33_X105Y83_IOB_X1Y83_OPAD,
  output RIOB33_X105Y83_IOB_X1Y84_OPAD,
  output RIOB33_X105Y85_IOB_X1Y85_OPAD,
  output RIOB33_X105Y85_IOB_X1Y86_OPAD,
  output RIOB33_X105Y87_IOB_X1Y87_OPAD,
  output RIOB33_X105Y87_IOB_X1Y88_OPAD,
  output RIOB33_X105Y89_IOB_X1Y89_OPAD,
  output RIOB33_X105Y89_IOB_X1Y90_OPAD,
  output RIOB33_X105Y91_IOB_X1Y91_OPAD,
  output RIOB33_X105Y91_IOB_X1Y92_OPAD,
  output RIOB33_X105Y93_IOB_X1Y93_OPAD,
  output RIOB33_X105Y93_IOB_X1Y94_OPAD,
  output RIOB33_X105Y95_IOB_X1Y95_OPAD,
  output RIOB33_X105Y95_IOB_X1Y96_OPAD,
  output RIOB33_X105Y97_IOB_X1Y97_OPAD,
  output RIOB33_X105Y97_IOB_X1Y98_OPAD
  );
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_ADDRARDADDR0;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_ADDRARDADDR1;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_ADDRARDADDR10;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_ADDRARDADDR11;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_ADDRARDADDR12;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_ADDRARDADDR13;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_ADDRARDADDR2;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_ADDRARDADDR3;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_ADDRARDADDR4;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_ADDRARDADDR5;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_ADDRARDADDR6;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_ADDRARDADDR7;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_ADDRARDADDR8;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_ADDRARDADDR9;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_ADDRATIEHIGH0;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_ADDRATIEHIGH1;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_ADDRBTIEHIGH0;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_ADDRBTIEHIGH1;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_ADDRBWRADDR0;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_ADDRBWRADDR1;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_ADDRBWRADDR10;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_ADDRBWRADDR11;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_ADDRBWRADDR12;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_ADDRBWRADDR13;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_ADDRBWRADDR2;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_ADDRBWRADDR3;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_ADDRBWRADDR4;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_ADDRBWRADDR5;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_ADDRBWRADDR6;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_ADDRBWRADDR7;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_ADDRBWRADDR8;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_ADDRBWRADDR9;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DIADI0;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DIADI1;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DIADI10;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DIADI11;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DIADI12;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DIADI13;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DIADI14;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DIADI15;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DIADI2;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DIADI3;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DIADI4;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DIADI5;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DIADI6;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DIADI7;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DIADI8;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DIADI9;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DIBDI0;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DIBDI1;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DIBDI10;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DIBDI11;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DIBDI12;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DIBDI13;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DIBDI14;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DIBDI15;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DIBDI2;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DIBDI3;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DIBDI4;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DIBDI5;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DIBDI6;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DIBDI7;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DIBDI8;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DIBDI9;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DIPADIP0;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DIPADIP1;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DIPBDIP0;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DIPBDIP1;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DO0;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DO1;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DO10;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DO11;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DO12;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DO13;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DO14;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DO15;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DO16;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DO17;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DO18;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DO19;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DO2;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DO20;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DO21;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DO22;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DO23;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DO24;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DO25;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DO26;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DO27;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DO28;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DO29;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DO3;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DO30;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DO31;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DO4;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DO5;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DO6;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DO7;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DO8;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DO9;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DOP0;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DOP1;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DOP2;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_DOP3;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_RDCLK;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_RDEN;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_RDRCLK;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_REGCE;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_REGCEB;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_REGCLKB;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_RST;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_RSTRAMB;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_RSTREG;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_RSTREGB;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_WEA0;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_WEA1;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_WEA2;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_WEA3;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_WEBWE0;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_WEBWE1;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_WEBWE2;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_WEBWE3;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_WEBWE4;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_WEBWE5;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_WEBWE6;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_WEBWE7;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_WRCLK;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y50_WREN;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_ADDRARDADDR0;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_ADDRARDADDR1;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_ADDRARDADDR10;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_ADDRARDADDR11;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_ADDRARDADDR12;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_ADDRARDADDR13;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_ADDRARDADDR2;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_ADDRARDADDR3;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_ADDRARDADDR4;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_ADDRARDADDR5;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_ADDRARDADDR6;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_ADDRARDADDR7;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_ADDRARDADDR8;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_ADDRARDADDR9;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_ADDRATIEHIGH0;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_ADDRATIEHIGH1;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_ADDRBTIEHIGH0;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_ADDRBTIEHIGH1;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_ADDRBWRADDR0;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_ADDRBWRADDR1;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_ADDRBWRADDR10;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_ADDRBWRADDR11;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_ADDRBWRADDR12;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_ADDRBWRADDR13;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_ADDRBWRADDR2;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_ADDRBWRADDR3;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_ADDRBWRADDR4;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_ADDRBWRADDR5;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_ADDRBWRADDR6;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_ADDRBWRADDR7;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_ADDRBWRADDR8;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_ADDRBWRADDR9;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_CLKARDCLK;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_CLKBWRCLK;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DIADI0;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DIADI1;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DIADI10;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DIADI11;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DIADI12;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DIADI13;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DIADI14;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DIADI15;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DIADI2;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DIADI3;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DIADI4;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DIADI5;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DIADI6;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DIADI7;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DIADI8;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DIADI9;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DIBDI0;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DIBDI1;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DIBDI10;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DIBDI11;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DIBDI12;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DIBDI13;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DIBDI14;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DIBDI15;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DIBDI2;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DIBDI3;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DIBDI4;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DIBDI5;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DIBDI6;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DIBDI7;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DIBDI8;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DIBDI9;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DIPADIP0;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DIPADIP1;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DIPBDIP0;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DIPBDIP1;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DOADO0;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DOADO1;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DOADO10;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DOADO11;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DOADO12;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DOADO13;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DOADO14;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DOADO15;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DOADO2;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DOADO3;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DOADO4;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DOADO5;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DOADO6;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DOADO7;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DOADO8;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DOADO9;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO0;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO1;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO10;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO11;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO12;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO13;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO14;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO15;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO2;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO3;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO4;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO5;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO6;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO7;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO8;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO9;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DOPADOP0;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DOPADOP1;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DOPBDOP0;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_DOPBDOP1;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_ENARDEN;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_ENBWREN;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_REGCEAREGCE;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_REGCEB;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_REGCLKARDRCLK;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_REGCLKB;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_RSTRAMARSTRAM;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_RSTRAMB;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_RSTREGARSTREG;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_RSTREGB;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_WEA0;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_WEA1;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_WEA2;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_WEA3;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_WEBWE0;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_WEBWE1;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_WEBWE2;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_WEBWE3;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_WEBWE4;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_WEBWE5;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_WEBWE6;
  wire [0:0] BRAM_L_X6Y125_RAMB18_X0Y51_WEBWE7;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_ADDRARDADDR0;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_ADDRARDADDR1;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_ADDRARDADDR10;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_ADDRARDADDR11;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_ADDRARDADDR12;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_ADDRARDADDR13;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_ADDRARDADDR2;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_ADDRARDADDR3;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_ADDRARDADDR4;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_ADDRARDADDR5;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_ADDRARDADDR6;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_ADDRARDADDR7;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_ADDRARDADDR8;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_ADDRARDADDR9;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_ADDRATIEHIGH0;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_ADDRATIEHIGH1;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_ADDRBTIEHIGH0;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_ADDRBTIEHIGH1;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_ADDRBWRADDR0;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_ADDRBWRADDR1;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_ADDRBWRADDR10;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_ADDRBWRADDR11;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_ADDRBWRADDR12;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_ADDRBWRADDR13;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_ADDRBWRADDR2;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_ADDRBWRADDR3;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_ADDRBWRADDR4;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_ADDRBWRADDR5;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_ADDRBWRADDR6;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_ADDRBWRADDR7;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_ADDRBWRADDR8;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_ADDRBWRADDR9;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DIADI0;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DIADI1;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DIADI10;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DIADI11;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DIADI12;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DIADI13;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DIADI14;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DIADI15;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DIADI2;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DIADI3;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DIADI4;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DIADI5;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DIADI6;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DIADI7;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DIADI8;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DIADI9;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DIBDI0;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DIBDI1;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DIBDI10;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DIBDI11;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DIBDI12;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DIBDI13;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DIBDI14;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DIBDI15;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DIBDI2;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DIBDI3;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DIBDI4;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DIBDI5;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DIBDI6;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DIBDI7;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DIBDI8;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DIBDI9;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DIPADIP0;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DIPADIP1;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DIPBDIP0;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DIPBDIP1;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DO0;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DO1;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DO10;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DO11;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DO12;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DO13;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DO14;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DO15;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DO16;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DO17;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DO18;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DO19;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DO2;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DO20;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DO21;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DO22;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DO23;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DO24;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DO25;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DO26;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DO27;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DO28;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DO29;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DO3;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DO30;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DO31;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DO4;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DO5;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DO6;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DO7;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DO8;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DO9;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DOP0;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DOP1;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DOP2;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_DOP3;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_RDCLK;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_RDEN;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_RDRCLK;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_REGCE;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_REGCEB;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_REGCLKB;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_RST;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_RSTRAMB;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_RSTREG;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_RSTREGB;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_WEA0;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_WEA1;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_WEA2;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_WEA3;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_WEBWE0;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_WEBWE1;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_WEBWE2;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_WEBWE3;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_WEBWE4;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_WEBWE5;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_WEBWE6;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_WEBWE7;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_WRCLK;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y52_WREN;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_ADDRARDADDR0;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_ADDRARDADDR1;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_ADDRARDADDR10;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_ADDRARDADDR11;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_ADDRARDADDR12;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_ADDRARDADDR13;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_ADDRARDADDR2;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_ADDRARDADDR3;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_ADDRARDADDR4;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_ADDRARDADDR5;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_ADDRARDADDR6;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_ADDRARDADDR7;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_ADDRARDADDR8;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_ADDRARDADDR9;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_ADDRATIEHIGH0;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_ADDRATIEHIGH1;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_ADDRBTIEHIGH0;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_ADDRBTIEHIGH1;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_ADDRBWRADDR0;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_ADDRBWRADDR1;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_ADDRBWRADDR10;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_ADDRBWRADDR11;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_ADDRBWRADDR12;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_ADDRBWRADDR13;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_ADDRBWRADDR2;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_ADDRBWRADDR3;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_ADDRBWRADDR4;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_ADDRBWRADDR5;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_ADDRBWRADDR6;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_ADDRBWRADDR7;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_ADDRBWRADDR8;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_ADDRBWRADDR9;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_CLKARDCLK;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_CLKBWRCLK;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DIADI0;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DIADI1;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DIADI10;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DIADI11;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DIADI12;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DIADI13;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DIADI14;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DIADI15;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DIADI2;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DIADI3;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DIADI4;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DIADI5;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DIADI6;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DIADI7;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DIADI8;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DIADI9;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DIBDI0;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DIBDI1;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DIBDI10;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DIBDI11;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DIBDI12;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DIBDI13;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DIBDI14;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DIBDI15;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DIBDI2;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DIBDI3;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DIBDI4;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DIBDI5;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DIBDI6;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DIBDI7;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DIBDI8;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DIBDI9;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DIPADIP0;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DIPADIP1;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DIPBDIP0;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DIPBDIP1;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DOADO0;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DOADO1;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DOADO10;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DOADO11;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DOADO12;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DOADO13;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DOADO14;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DOADO15;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DOADO2;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DOADO3;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DOADO4;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DOADO5;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DOADO6;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DOADO7;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DOADO8;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DOADO9;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO0;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO1;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO10;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO11;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO12;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO13;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO14;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO15;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO2;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO3;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO4;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO5;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO6;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO7;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO8;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO9;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DOPADOP0;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DOPADOP1;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DOPBDOP0;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_DOPBDOP1;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_ENARDEN;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_ENBWREN;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_REGCEAREGCE;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_REGCEB;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_REGCLKARDRCLK;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_REGCLKB;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_RSTRAMARSTRAM;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_RSTRAMB;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_RSTREGARSTREG;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_RSTREGB;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_WEA0;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_WEA1;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_WEA2;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_WEA3;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_WEBWE0;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_WEBWE1;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_WEBWE2;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_WEBWE3;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_WEBWE4;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_WEBWE5;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_WEBWE6;
  wire [0:0] BRAM_L_X6Y130_RAMB18_X0Y53_WEBWE7;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_ADDRARDADDR0;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_ADDRARDADDR1;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_ADDRARDADDR10;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_ADDRARDADDR11;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_ADDRARDADDR12;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_ADDRARDADDR13;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_ADDRARDADDR2;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_ADDRARDADDR3;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_ADDRARDADDR4;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_ADDRARDADDR5;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_ADDRARDADDR6;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_ADDRARDADDR7;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_ADDRARDADDR8;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_ADDRARDADDR9;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_ADDRATIEHIGH0;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_ADDRATIEHIGH1;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_ADDRBTIEHIGH0;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_ADDRBTIEHIGH1;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_ADDRBWRADDR0;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_ADDRBWRADDR1;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_ADDRBWRADDR10;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_ADDRBWRADDR11;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_ADDRBWRADDR12;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_ADDRBWRADDR13;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_ADDRBWRADDR2;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_ADDRBWRADDR3;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_ADDRBWRADDR4;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_ADDRBWRADDR5;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_ADDRBWRADDR6;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_ADDRBWRADDR7;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_ADDRBWRADDR8;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_ADDRBWRADDR9;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DIADI0;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DIADI1;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DIADI10;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DIADI11;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DIADI12;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DIADI13;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DIADI14;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DIADI15;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DIADI2;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DIADI3;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DIADI4;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DIADI5;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DIADI6;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DIADI7;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DIADI8;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DIADI9;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DIBDI0;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DIBDI1;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DIBDI10;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DIBDI11;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DIBDI12;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DIBDI13;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DIBDI14;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DIBDI15;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DIBDI2;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DIBDI3;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DIBDI4;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DIBDI5;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DIBDI6;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DIBDI7;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DIBDI8;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DIBDI9;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DIPADIP0;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DIPADIP1;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DIPBDIP0;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DIPBDIP1;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DO0;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DO1;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DO10;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DO11;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DO12;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DO13;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DO14;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DO15;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DO16;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DO17;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DO18;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DO19;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DO2;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DO20;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DO21;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DO22;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DO23;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DO24;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DO25;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DO26;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DO27;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DO28;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DO29;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DO3;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DO30;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DO31;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DO4;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DO5;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DO6;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DO7;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DO8;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DO9;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DOP0;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DOP1;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DOP2;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_DOP3;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_RDCLK;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_RDEN;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_RDRCLK;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_REGCE;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_REGCEB;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_REGCLKB;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_RST;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_RSTRAMB;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_RSTREG;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_RSTREGB;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_WEA0;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_WEA1;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_WEA2;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_WEA3;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_WEBWE0;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_WEBWE1;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_WEBWE2;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_WEBWE3;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_WEBWE4;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_WEBWE5;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_WEBWE6;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_WEBWE7;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_WRCLK;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y54_WREN;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_ADDRARDADDR0;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_ADDRARDADDR1;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_ADDRARDADDR10;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_ADDRARDADDR11;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_ADDRARDADDR12;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_ADDRARDADDR13;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_ADDRARDADDR2;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_ADDRARDADDR3;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_ADDRARDADDR4;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_ADDRARDADDR5;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_ADDRARDADDR6;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_ADDRARDADDR7;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_ADDRARDADDR8;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_ADDRARDADDR9;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_ADDRATIEHIGH0;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_ADDRATIEHIGH1;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_ADDRBTIEHIGH0;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_ADDRBTIEHIGH1;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_ADDRBWRADDR0;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_ADDRBWRADDR1;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_ADDRBWRADDR10;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_ADDRBWRADDR11;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_ADDRBWRADDR12;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_ADDRBWRADDR13;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_ADDRBWRADDR2;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_ADDRBWRADDR3;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_ADDRBWRADDR4;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_ADDRBWRADDR5;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_ADDRBWRADDR6;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_ADDRBWRADDR7;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_ADDRBWRADDR8;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_ADDRBWRADDR9;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_CLKARDCLK;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_CLKBWRCLK;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DIADI0;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DIADI1;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DIADI10;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DIADI11;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DIADI12;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DIADI13;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DIADI14;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DIADI15;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DIADI2;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DIADI3;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DIADI4;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DIADI5;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DIADI6;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DIADI7;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DIADI8;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DIADI9;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DIBDI0;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DIBDI1;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DIBDI10;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DIBDI11;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DIBDI12;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DIBDI13;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DIBDI14;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DIBDI15;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DIBDI2;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DIBDI3;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DIBDI4;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DIBDI5;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DIBDI6;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DIBDI7;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DIBDI8;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DIBDI9;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DIPADIP0;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DIPADIP1;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DIPBDIP0;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DIPBDIP1;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DOADO0;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DOADO1;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DOADO10;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DOADO11;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DOADO12;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DOADO13;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DOADO14;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DOADO15;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DOADO2;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DOADO3;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DOADO4;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DOADO5;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DOADO6;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DOADO7;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DOADO8;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DOADO9;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO0;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO1;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO10;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO11;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO12;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO13;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO14;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO15;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO2;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO3;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO4;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO5;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO6;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO7;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO8;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO9;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DOPADOP0;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DOPADOP1;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DOPBDOP0;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_DOPBDOP1;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_ENARDEN;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_ENBWREN;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_REGCEAREGCE;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_REGCEB;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_REGCLKARDRCLK;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_REGCLKB;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_RSTRAMARSTRAM;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_RSTRAMB;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_RSTREGARSTREG;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_RSTREGB;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_WEA0;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_WEA1;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_WEA2;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_WEA3;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_WEBWE0;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_WEBWE1;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_WEBWE2;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_WEBWE3;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_WEBWE4;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_WEBWE5;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_WEBWE6;
  wire [0:0] BRAM_L_X6Y135_RAMB18_X0Y55_WEBWE7;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_ADDRARDADDR0;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_ADDRARDADDR1;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_ADDRARDADDR10;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_ADDRARDADDR11;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_ADDRARDADDR12;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_ADDRARDADDR13;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_ADDRARDADDR2;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_ADDRARDADDR3;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_ADDRARDADDR4;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_ADDRARDADDR5;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_ADDRARDADDR6;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_ADDRARDADDR7;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_ADDRARDADDR8;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_ADDRARDADDR9;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_ADDRATIEHIGH0;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_ADDRATIEHIGH1;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_ADDRBTIEHIGH0;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_ADDRBTIEHIGH1;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_ADDRBWRADDR0;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_ADDRBWRADDR1;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_ADDRBWRADDR10;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_ADDRBWRADDR11;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_ADDRBWRADDR12;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_ADDRBWRADDR13;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_ADDRBWRADDR2;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_ADDRBWRADDR3;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_ADDRBWRADDR4;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_ADDRBWRADDR5;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_ADDRBWRADDR6;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_ADDRBWRADDR7;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_ADDRBWRADDR8;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_ADDRBWRADDR9;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DIADI0;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DIADI1;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DIADI10;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DIADI11;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DIADI12;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DIADI13;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DIADI14;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DIADI15;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DIADI2;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DIADI3;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DIADI4;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DIADI5;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DIADI6;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DIADI7;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DIADI8;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DIADI9;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DIBDI0;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DIBDI1;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DIBDI10;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DIBDI11;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DIBDI12;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DIBDI13;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DIBDI14;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DIBDI15;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DIBDI2;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DIBDI3;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DIBDI4;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DIBDI5;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DIBDI6;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DIBDI7;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DIBDI8;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DIBDI9;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DIPADIP0;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DIPADIP1;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DIPBDIP0;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DIPBDIP1;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DO0;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DO1;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DO10;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DO11;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DO12;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DO13;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DO14;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DO15;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DO16;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DO17;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DO18;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DO19;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DO2;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DO20;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DO21;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DO22;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DO23;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DO24;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DO25;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DO26;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DO27;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DO28;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DO29;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DO3;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DO30;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DO31;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DO4;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DO5;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DO6;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DO7;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DO8;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DO9;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DOP0;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DOP1;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DOP2;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_DOP3;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_RDCLK;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_RDEN;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_RDRCLK;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_REGCE;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_REGCEB;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_REGCLKB;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_RST;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_RSTRAMB;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_RSTREG;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_RSTREGB;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_WEA0;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_WEA1;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_WEA2;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_WEA3;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_WEBWE0;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_WEBWE1;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_WEBWE2;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_WEBWE3;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_WEBWE4;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_WEBWE5;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_WEBWE6;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_WEBWE7;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_WRCLK;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y56_WREN;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_ADDRARDADDR0;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_ADDRARDADDR1;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_ADDRARDADDR10;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_ADDRARDADDR11;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_ADDRARDADDR12;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_ADDRARDADDR13;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_ADDRARDADDR2;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_ADDRARDADDR3;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_ADDRARDADDR4;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_ADDRARDADDR5;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_ADDRARDADDR6;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_ADDRARDADDR7;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_ADDRARDADDR8;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_ADDRARDADDR9;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_ADDRATIEHIGH0;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_ADDRATIEHIGH1;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_ADDRBTIEHIGH0;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_ADDRBTIEHIGH1;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_ADDRBWRADDR0;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_ADDRBWRADDR1;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_ADDRBWRADDR10;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_ADDRBWRADDR11;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_ADDRBWRADDR12;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_ADDRBWRADDR13;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_ADDRBWRADDR2;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_ADDRBWRADDR3;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_ADDRBWRADDR4;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_ADDRBWRADDR5;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_ADDRBWRADDR6;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_ADDRBWRADDR7;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_ADDRBWRADDR8;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_ADDRBWRADDR9;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_CLKARDCLK;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_CLKBWRCLK;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DIADI0;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DIADI1;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DIADI10;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DIADI11;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DIADI12;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DIADI13;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DIADI14;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DIADI15;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DIADI2;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DIADI3;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DIADI4;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DIADI5;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DIADI6;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DIADI7;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DIADI8;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DIADI9;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DIBDI0;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DIBDI1;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DIBDI10;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DIBDI11;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DIBDI12;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DIBDI13;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DIBDI14;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DIBDI15;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DIBDI2;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DIBDI3;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DIBDI4;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DIBDI5;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DIBDI6;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DIBDI7;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DIBDI8;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DIBDI9;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DIPADIP0;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DIPADIP1;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DIPBDIP0;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DIPBDIP1;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DOADO0;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DOADO1;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DOADO10;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DOADO11;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DOADO12;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DOADO13;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DOADO14;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DOADO15;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DOADO2;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DOADO3;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DOADO4;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DOADO5;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DOADO6;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DOADO7;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DOADO8;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DOADO9;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO0;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO1;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO10;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO11;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO12;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO13;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO14;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO15;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO2;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO3;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO4;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO5;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO6;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO7;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO8;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO9;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DOPADOP0;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DOPADOP1;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DOPBDOP0;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_DOPBDOP1;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_ENARDEN;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_ENBWREN;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_REGCEAREGCE;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_REGCEB;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_REGCLKARDRCLK;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_REGCLKB;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_RSTRAMARSTRAM;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_RSTRAMB;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_RSTREGARSTREG;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_RSTREGB;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_WEA0;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_WEA1;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_WEA2;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_WEA3;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_WEBWE0;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_WEBWE1;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_WEBWE2;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_WEBWE3;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_WEBWE4;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_WEBWE5;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_WEBWE6;
  wire [0:0] BRAM_L_X6Y140_RAMB18_X0Y57_WEBWE7;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_ADDRARDADDR0;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_ADDRARDADDR1;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_ADDRARDADDR10;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_ADDRARDADDR11;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_ADDRARDADDR12;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_ADDRARDADDR13;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_ADDRARDADDR2;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_ADDRARDADDR3;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_ADDRARDADDR4;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_ADDRARDADDR5;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_ADDRARDADDR6;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_ADDRARDADDR7;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_ADDRARDADDR8;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_ADDRARDADDR9;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_ADDRATIEHIGH0;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_ADDRATIEHIGH1;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_ADDRBTIEHIGH0;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_ADDRBTIEHIGH1;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_ADDRBWRADDR0;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_ADDRBWRADDR1;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_ADDRBWRADDR10;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_ADDRBWRADDR11;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_ADDRBWRADDR12;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_ADDRBWRADDR13;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_ADDRBWRADDR2;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_ADDRBWRADDR3;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_ADDRBWRADDR4;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_ADDRBWRADDR5;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_ADDRBWRADDR6;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_ADDRBWRADDR7;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_ADDRBWRADDR8;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_ADDRBWRADDR9;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DIADI0;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DIADI1;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DIADI10;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DIADI11;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DIADI12;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DIADI13;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DIADI14;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DIADI15;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DIADI2;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DIADI3;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DIADI4;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DIADI5;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DIADI6;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DIADI7;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DIADI8;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DIADI9;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DIBDI0;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DIBDI1;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DIBDI10;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DIBDI11;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DIBDI12;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DIBDI13;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DIBDI14;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DIBDI15;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DIBDI2;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DIBDI3;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DIBDI4;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DIBDI5;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DIBDI6;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DIBDI7;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DIBDI8;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DIBDI9;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DIPADIP0;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DIPADIP1;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DIPBDIP0;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DIPBDIP1;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DO0;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DO1;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DO10;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DO11;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DO12;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DO13;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DO14;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DO15;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DO16;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DO17;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DO18;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DO19;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DO2;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DO20;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DO21;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DO22;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DO23;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DO24;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DO25;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DO26;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DO27;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DO28;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DO29;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DO3;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DO30;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DO31;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DO4;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DO5;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DO6;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DO7;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DO8;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DO9;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DOP0;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DOP1;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DOP2;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_DOP3;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_RDCLK;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_RDEN;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_RDRCLK;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_REGCE;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_REGCEB;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_REGCLKB;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_RST;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_RSTRAMB;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_RSTREG;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_RSTREGB;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_WEA0;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_WEA1;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_WEA2;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_WEA3;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_WEBWE0;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_WEBWE1;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_WEBWE2;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_WEBWE3;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_WEBWE4;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_WEBWE5;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_WEBWE6;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_WEBWE7;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_WRCLK;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y54_WREN;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_ADDRARDADDR0;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_ADDRARDADDR1;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_ADDRARDADDR10;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_ADDRARDADDR11;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_ADDRARDADDR12;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_ADDRARDADDR13;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_ADDRARDADDR2;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_ADDRARDADDR3;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_ADDRARDADDR4;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_ADDRARDADDR5;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_ADDRARDADDR6;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_ADDRARDADDR7;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_ADDRARDADDR8;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_ADDRARDADDR9;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_ADDRATIEHIGH0;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_ADDRATIEHIGH1;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_ADDRBTIEHIGH0;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_ADDRBTIEHIGH1;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_ADDRBWRADDR0;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_ADDRBWRADDR1;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_ADDRBWRADDR10;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_ADDRBWRADDR11;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_ADDRBWRADDR12;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_ADDRBWRADDR13;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_ADDRBWRADDR2;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_ADDRBWRADDR3;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_ADDRBWRADDR4;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_ADDRBWRADDR5;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_ADDRBWRADDR6;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_ADDRBWRADDR7;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_ADDRBWRADDR8;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_ADDRBWRADDR9;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_CLKARDCLK;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_CLKBWRCLK;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DIADI0;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DIADI1;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DIADI10;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DIADI11;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DIADI12;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DIADI13;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DIADI14;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DIADI15;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DIADI2;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DIADI3;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DIADI4;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DIADI5;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DIADI6;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DIADI7;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DIADI8;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DIADI9;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DIBDI0;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DIBDI1;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DIBDI10;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DIBDI11;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DIBDI12;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DIBDI13;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DIBDI14;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DIBDI15;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DIBDI2;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DIBDI3;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DIBDI4;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DIBDI5;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DIBDI6;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DIBDI7;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DIBDI8;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DIBDI9;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DIPADIP0;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DIPADIP1;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DIPBDIP0;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DIPBDIP1;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DOADO0;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DOADO1;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DOADO10;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DOADO11;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DOADO12;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DOADO13;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DOADO14;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DOADO15;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DOADO2;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DOADO3;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DOADO4;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DOADO5;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DOADO6;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DOADO7;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DOADO8;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DOADO9;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO0;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO1;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO10;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO11;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO12;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO13;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO14;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO15;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO2;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO3;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO4;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO5;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO6;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO7;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO8;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO9;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DOPADOP0;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DOPADOP1;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DOPBDOP0;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_DOPBDOP1;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_ENARDEN;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_ENBWREN;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_REGCEAREGCE;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_REGCEB;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_REGCLKARDRCLK;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_REGCLKB;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_RSTRAMARSTRAM;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_RSTRAMB;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_RSTREGARSTREG;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_RSTREGB;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_WEA0;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_WEA1;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_WEA2;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_WEA3;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_WEBWE0;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_WEBWE1;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_WEBWE2;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_WEBWE3;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_WEBWE4;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_WEBWE5;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_WEBWE6;
  wire [0:0] BRAM_R_X17Y135_RAMB18_X1Y55_WEBWE7;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_AO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_AO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_BO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_BO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_CO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_CO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_DO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_DO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A5Q;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_AMUX;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_AO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_AO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_AQ;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_BO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_BO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_BQ;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_CLK;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_CO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_CO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_DO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_DO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_SR;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_A;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_A1;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_A2;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_A3;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_A4;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_A5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_A6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_AO5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_AO6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_A_CY;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_A_XOR;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_B;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_B1;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_B2;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_B3;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_B4;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_B5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_B6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_BO5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_BO6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_B_CY;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_B_XOR;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_C;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_C1;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_C2;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_C3;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_C4;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_C5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_C6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_CO5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_CO6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_C_CY;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_C_XOR;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_D;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_D1;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_D2;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_D3;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_D4;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_D5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_D6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_DO5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_DO6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_D_CY;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_D_XOR;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_A;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_A1;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_A2;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_A3;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_A4;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_A5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_A6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_AO5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_AO6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_AQ;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_A_CY;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_A_XOR;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_B;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_B1;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_B2;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_B3;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_B4;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_B5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_B6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_BO5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_BO6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_B_CY;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_B_XOR;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_C;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_C1;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_C2;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_C3;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_C4;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_C5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_C6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_CLK;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_CO5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_CO6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_C_CY;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_C_XOR;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_D;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_D1;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_D2;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_D3;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_D4;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_D5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_D6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_DO5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_DO6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_D_CY;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_D_XOR;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_A;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_A1;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_A2;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_A3;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_A4;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_A5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_A6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_AO5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_AO6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_AQ;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_A_CY;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_A_XOR;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_B;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_B1;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_B2;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_B3;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_B4;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_B5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_B6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_BO5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_BO6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_B_CY;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_B_XOR;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_C;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_C1;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_C2;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_C3;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_C4;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_C5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_C6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_CLK;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_CO5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_CO6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_C_CY;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_C_XOR;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_D;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_D1;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_D2;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_D3;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_D4;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_D5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_D6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_DO5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_DO6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_D_CY;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_D_XOR;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_A;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_A1;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_A2;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_A3;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_A4;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_A5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_A6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_AO5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_AO6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_A_CY;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_A_XOR;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_B;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_B1;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_B2;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_B3;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_B4;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_B5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_B6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_BO5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_BO6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_B_CY;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_B_XOR;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_C;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_C1;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_C2;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_C3;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_C4;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_C5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_C6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_CO5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_CO6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_C_CY;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_C_XOR;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_D;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_D1;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_D2;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_D3;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_D4;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_D5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_D6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_DO5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_DO6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_D_CY;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_D_XOR;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_A;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_A1;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_A2;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_A3;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_A4;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_A5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_A6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_AO5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_AO6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_AQ;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_A_CY;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_A_XOR;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_B;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_B1;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_B2;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_B3;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_B4;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_B5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_B6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_BO5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_BO6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_BQ;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_B_CY;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_B_XOR;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_C;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_C1;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_C2;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_C3;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_C4;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_C5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_C6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_CLK;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_CO5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_CO6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_CQ;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_C_CY;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_C_XOR;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_D;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_D1;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_D2;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_D3;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_D4;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_D5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_D6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_DO5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_DO6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_DQ;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_D_CY;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_D_XOR;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_A;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_A1;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_A2;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_A3;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_A4;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_A5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_A6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_AO5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_AO6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_A_CY;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_A_XOR;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_B;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_B1;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_B2;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_B3;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_B4;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_B5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_B6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_BO5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_BO6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_B_CY;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_B_XOR;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_C;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_C1;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_C2;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_C3;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_C4;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_C5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_C6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_CO5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_CO6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_C_CY;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_C_XOR;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_D;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_D1;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_D2;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_D3;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_D4;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_D5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_D6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_DO5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_DO6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_D_CY;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_D_XOR;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_A;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_A1;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_A2;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_A3;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_A4;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_A5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_A6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_AO5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_AO6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_AQ;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_AX;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_A_CY;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_A_XOR;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_B;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_B1;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_B2;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_B3;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_B4;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_B5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_B6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_BO5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_BO6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_B_CY;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_B_XOR;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_C;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_C1;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_C2;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_C3;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_C4;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_C5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_C6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_CE;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_CLK;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_CO5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_CO6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_C_CY;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_C_XOR;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_D;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_D1;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_D2;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_D3;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_D4;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_D5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_D6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_DO5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_DO6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_D_CY;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_D_XOR;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_A;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_A1;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_A2;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_A3;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_A4;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_A5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_A6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_AO5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_AO6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_A_CY;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_A_XOR;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_B;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_B1;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_B2;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_B3;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_B4;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_B5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_B6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_BO5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_BO6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_B_CY;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_B_XOR;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_C;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_C1;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_C2;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_C3;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_C4;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_C5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_C6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_CO5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_CO6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_C_CY;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_C_XOR;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_D;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_D1;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_D2;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_D3;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_D4;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_D5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_D6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_DO5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_DO6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_D_CY;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_D_XOR;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_A;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_A1;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_A2;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_A3;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_A4;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_A5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_A6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_AO5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_AO6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_AQ;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_AX;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_A_CY;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_A_XOR;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_B;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_B1;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_B2;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_B3;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_B4;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_B5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_B6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_BO5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_BO6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_BQ;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_BX;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_B_CY;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_B_XOR;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_C;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_C1;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_C2;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_C3;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_C4;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_C5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_C6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_CE;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_CLK;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_CO5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_CO6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_CQ;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_CX;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_C_CY;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_C_XOR;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_D;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_D1;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_D2;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_D3;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_D4;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_D5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_D6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_DO5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_DO6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_DQ;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_DX;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_D_CY;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_D_XOR;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_A;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_A1;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_A2;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_A3;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_A4;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_A5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_A6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_AO5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_AO6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_AQ;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_AX;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_A_CY;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_A_XOR;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_B;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_B1;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_B2;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_B3;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_B4;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_B5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_B6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_BO5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_BO6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_BQ;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_BX;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_B_CY;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_B_XOR;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_C;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_C1;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_C2;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_C3;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_C4;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_C5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_C6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_CE;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_CLK;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_CO5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_CO6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_C_CY;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_C_XOR;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_D;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_D1;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_D2;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_D3;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_D4;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_D5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_D6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_DO5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_D_CY;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_D_XOR;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_A;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_A1;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_A2;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_A3;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_A4;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_A5;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_A6;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_AO5;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_AO6;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_AQ;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_AX;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_A_CY;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_A_XOR;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_B;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_B1;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_B2;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_B3;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_B4;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_B5;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_B6;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_BO5;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_BO6;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_BQ;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_BX;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_B_CY;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_B_XOR;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_C;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_C1;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_C2;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_C3;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_C4;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_C5;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_C6;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_CE;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_CLK;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_CO5;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_CO6;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_CQ;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_CX;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_C_CY;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_C_XOR;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_D;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_D1;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_D2;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_D3;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_D4;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_D5;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_D6;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_DO5;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_DO6;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_DQ;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_DX;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_D_CY;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_D_XOR;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_A;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_A1;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_A2;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_A3;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_A4;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_A5;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_A6;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_AO5;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_AO6;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_AQ;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_AX;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_A_CY;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_A_XOR;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_B;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_B1;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_B2;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_B3;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_B4;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_B5;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_B6;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_BO5;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_BO6;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_BQ;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_BX;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_B_CY;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_B_XOR;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_C;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_C1;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_C2;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_C3;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_C4;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_C5;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_C6;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_CE;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_CLK;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_CO5;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_CO6;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_C_CY;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_C_XOR;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_D;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_D1;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_D2;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_D3;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_D4;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_D5;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_D6;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_DO5;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_DO6;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_D_CY;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_D_XOR;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_A;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_A1;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_A2;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_A3;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_A4;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_A5;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_A6;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_AO5;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_AO6;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_AQ;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_AX;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_A_CY;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_A_XOR;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_B;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_B1;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_B2;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_B3;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_B4;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_B5;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_B6;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_BO5;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_BO6;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_BQ;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_BX;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_B_CY;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_B_XOR;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_C;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_C1;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_C2;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_C3;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_C4;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_C5;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_C6;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_CE;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_CLK;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_CO5;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_CO6;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_CQ;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_CX;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_C_CY;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_C_XOR;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_D;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_D1;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_D2;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_D3;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_D4;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_D5;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_D6;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_DO5;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_DO6;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_DQ;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_DX;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_D_CY;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_D_XOR;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_A;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_A1;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_A2;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_A3;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_A4;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_A5;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_A6;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_AO5;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_AO6;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_A_CY;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_A_XOR;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_B;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_B1;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_B2;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_B3;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_B4;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_B5;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_B6;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_BO5;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_BO6;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_B_CY;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_B_XOR;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_C;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_C1;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_C2;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_C3;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_C4;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_C5;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_C6;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_CO5;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_CO6;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_C_CY;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_C_XOR;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_D;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_D1;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_D2;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_D3;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_D4;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_D5;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_D6;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_DO5;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_DO6;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_D_CY;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_D_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_AO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_AO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_BO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_BO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_CO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_CO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_DO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_DO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_AO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_AO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_AQ;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_BO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_BO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_CLK;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_CO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_CO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_DO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_DO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_AO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_AO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_BO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_BO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_CO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_CO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_DO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_DO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_AMUX;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_AO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_AO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_AQ;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_BO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_BO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_BQ;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_CLK;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_CO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_CO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_DO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_DO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_AO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_AO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_AQ;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_AX;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_BO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_BO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_CLK;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_CO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_CO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_DO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_DO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_AMUX;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_AO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_AO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_AQ;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_BMUX;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_BO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_BO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_CLK;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_CO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_CO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_CQ;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_DO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_DO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_AMUX;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_AO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_AO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_BO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_BO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_BQ;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_CLK;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_CO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_CO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_DO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_DO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A5Q;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_AMUX;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_AO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_AO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_AQ;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_AX;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_BO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_BO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_BX;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_CLK;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_CO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_CO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_DMUX;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_DO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_DO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_AMUX;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_AO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_AO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_AQ;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_AX;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_BMUX;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_BO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_BQ;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_CLK;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_CO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_CO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_CQ;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_DO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_DO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_DQ;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_AMUX;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_AO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_AO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_AQ;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_AX;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B5Q;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_BMUX;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_BO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_BO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_BQ;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_BX;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_CLK;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_CO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_CO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_CQ;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_DO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_DO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_AMUX;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_AO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_AO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_AQ;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_BMUX;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_BO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_BO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_BQ;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_CLK;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_CO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_CO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_CQ;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_DMUX;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_DO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_DO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A5Q;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_AMUX;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_AO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_AO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_AX;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_BO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_BO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_BQ;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_CLK;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_CO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_CO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_DO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_DO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A5Q;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_AMUX;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_AO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_AO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_AQ;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_AX;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_BO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_BO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_BQ;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_CLK;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_CMUX;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_CO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_CO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_DO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_DO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_AMUX;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_AO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_AO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_AQ;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_BO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_BO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_BQ;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_CLK;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_CO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_CO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_DO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_DO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_AO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_AO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_AQ;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_AX;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_BO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_BO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_CLK;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_CO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_CO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_DO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_DO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_AO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_AO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_AQ;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_BO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_BO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_BQ;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_CLK;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_CO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_CO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_DO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_DO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_AMUX;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_AO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_AO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_BO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_BO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_CO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_CO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_DO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_DO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_AMUX;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_AO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_AO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_BO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_BO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_BQ;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_CLK;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_CO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_CO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_DO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_DO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_AO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_AO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_BO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_BO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_CO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_CO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_DO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_DO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_AO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_AO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_BO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_BO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_CMUX;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_CO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_CO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_DO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_DO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_AO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_AO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_BMUX;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_BO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_BO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_CO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_CO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_DO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_DO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_AMUX;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_AO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_AO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_BMUX;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_BO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_BO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_CO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_CO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_DO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_DO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_AO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_AO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_BMUX;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_BO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_BO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_CO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_CO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_DO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_DO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_AO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_AO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_BO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_BO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_CO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_CO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_DO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_DO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_AO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_AO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_BO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_BO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_CO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_CO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_DO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_DO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_AO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_AO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_BO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_BO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_CO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_CO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_DO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_DO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_AO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_AO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_BO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_BO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_CO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_CO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_DO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_DO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_AMUX;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_AO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_BO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_BO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_CO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_CO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_DO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_DO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_AO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_AO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_AQ;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_AX;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_BO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_BO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_BQ;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_BX;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_CE;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_CLK;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_CO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_CO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_DO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_DO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_AO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_AO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_BO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_BO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_CO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_CO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_DO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_DO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_AO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_AO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_AQ;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_AX;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_BO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_BO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_CE;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_CLK;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_CO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_CO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_DO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_DO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_AO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_AO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_BO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_BO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_CO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_CO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_DO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_DO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D_XOR;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_A;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_A1;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_A2;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_A3;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_A4;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_A5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_A6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_AO5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_AO6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_AQ;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_AX;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_A_CY;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_A_XOR;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_B;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_B1;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_B2;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_B3;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_B4;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_B5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_B6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_BO5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_BO6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_BQ;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_BX;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_B_CY;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_B_XOR;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_C;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_C1;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_C2;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_C3;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_C4;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_C5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_C6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_CE;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_CLK;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_CO5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_CO6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_CQ;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_CX;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_C_CY;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_C_XOR;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_D;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_D1;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_D2;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_D3;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_D4;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_D5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_D6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_DO5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_DO6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_DQ;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_DX;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_D_CY;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_D_XOR;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_A;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_A1;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_A2;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_A3;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_A4;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_A5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_A6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_AO5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_AO6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_A_CY;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_A_XOR;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_B;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_B1;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_B2;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_B3;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_B4;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_B5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_B6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_BO5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_BO6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_B_CY;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_B_XOR;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_C;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_C1;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_C2;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_C3;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_C4;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_C5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_C6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_CO5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_CO6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_C_CY;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_C_XOR;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_D;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_D1;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_D2;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_D3;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_D4;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_D5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_D6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_DO5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_DO6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_D_CY;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_D_XOR;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_A;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_A1;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_A2;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_A3;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_A4;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_A5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_A6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_AO5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_AO6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_AQ;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_AX;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_A_CY;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_A_XOR;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_B;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_B1;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_B2;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_B3;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_B4;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_B5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_B6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_BO5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_BO6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_BQ;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_BX;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_B_CY;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_B_XOR;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_C;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_C1;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_C2;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_C3;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_C4;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_C5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_C6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_CE;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_CLK;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_CO5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_CO6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_CQ;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_CX;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_C_CY;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_C_XOR;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_D;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_D1;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_D2;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_D3;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_D4;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_D5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_D6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_DO5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_DO6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_DQ;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_DX;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_D_CY;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_D_XOR;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_A;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_A1;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_A2;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_A3;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_A4;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_A5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_A5Q;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_A6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_AMUX;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_AO5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_AO6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_AQ;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_AX;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_A_CY;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_A_XOR;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_B;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_B1;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_B2;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_B3;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_B4;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_B5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_B6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_BO5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_BO6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_BQ;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_BX;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_B_CY;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_B_XOR;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_C;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_C1;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_C2;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_C3;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_C4;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_C5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_C6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_CE;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_CLK;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_CO5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_CO6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_CQ;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_CX;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_C_CY;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_C_XOR;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_D;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_D1;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_D2;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_D3;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_D4;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_D5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_D6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_DO5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_DO6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_DQ;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_DX;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_D_CY;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_D_XOR;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_A;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_A1;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_A2;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_A3;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_A4;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_A5;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_A6;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_AO5;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_AO6;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_AQ;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_AX;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_A_CY;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_A_XOR;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_B;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_B1;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_B2;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_B3;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_B4;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_B5;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_B6;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_BO5;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_BO6;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_B_CY;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_B_XOR;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_C;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_C1;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_C2;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_C3;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_C4;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_C5;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_C6;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_CLK;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_CO5;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_CO6;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_C_CY;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_C_XOR;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_D;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_D1;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_D2;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_D3;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_D4;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_D5;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_D6;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_DO5;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_DO6;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_D_CY;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_D_XOR;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_A;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_A1;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_A2;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_A3;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_A4;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_A5;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_A6;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_AO5;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_AO6;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_A_CY;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_A_XOR;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_B;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_B1;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_B2;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_B3;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_B4;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_B5;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_B6;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_BO5;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_BO6;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_B_CY;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_B_XOR;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_C;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_C1;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_C2;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_C3;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_C4;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_C5;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_C6;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_CO5;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_CO6;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_C_CY;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_C_XOR;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_D;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_D1;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_D2;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_D3;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_D4;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_D5;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_D6;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_DO5;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_DO6;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_D_CY;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_D_XOR;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_A;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_A1;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_A2;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_A3;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_A4;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_A5;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_A6;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_AO5;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_AO6;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_AQ;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_AX;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_A_CY;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_A_XOR;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_B;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_B1;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_B2;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_B3;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_B4;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_B5;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_B6;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_BO5;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_BO6;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_B_CY;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_B_XOR;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_C;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_C1;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_C2;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_C3;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_C4;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_C5;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_C6;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_CLK;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_CO5;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_CO6;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_C_CY;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_C_XOR;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_D;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_D1;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_D2;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_D3;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_D4;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_D5;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_D6;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_DO5;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_DO6;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_D_CY;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_D_XOR;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_A;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_A1;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_A2;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_A3;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_A4;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_A5;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_A6;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_AO5;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_AO6;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_A_CY;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_A_XOR;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_B;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_B1;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_B2;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_B3;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_B4;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_B5;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_B6;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_BO5;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_BO6;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_B_CY;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_B_XOR;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_C;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_C1;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_C2;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_C3;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_C4;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_C5;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_C6;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_CO5;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_CO6;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_C_CY;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_C_XOR;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_D;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_D1;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_D2;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_D3;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_D4;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_D5;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_D6;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_DO5;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_DO6;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_D_CY;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_D_XOR;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_A;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_A1;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_A2;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_A3;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_A4;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_A5;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_A6;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_AO5;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_AO6;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_AQ;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_AX;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_A_CY;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_A_XOR;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_B;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_B1;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_B2;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_B3;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_B4;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_B5;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_B6;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_BO5;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_BO6;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_B_CY;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_B_XOR;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_C;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_C1;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_C2;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_C3;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_C4;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_C5;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_C6;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_CLK;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_CO5;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_CO6;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_C_CY;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_C_XOR;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_D;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_D1;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_D2;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_D3;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_D4;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_D5;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_D6;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_DO5;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_DO6;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_D_CY;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X82Y116_D_XOR;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_A;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_A1;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_A2;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_A3;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_A4;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_A5;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_A6;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_AO5;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_AO6;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_A_CY;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_A_XOR;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_B;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_B1;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_B2;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_B3;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_B4;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_B5;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_B6;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_BO5;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_BO6;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_B_CY;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_B_XOR;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_C;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_C1;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_C2;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_C3;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_C4;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_C5;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_C6;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_CO5;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_CO6;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_C_CY;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_C_XOR;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_D;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_D1;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_D2;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_D3;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_D4;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_D5;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_D6;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_DO5;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_DO6;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_D_CY;
  wire [0:0] CLBLL_L_X54Y116_SLICE_X83Y116_D_XOR;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_A;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_A1;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_A2;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_A3;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_A4;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_A5;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_A6;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_AO5;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_AO6;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_AQ;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_AX;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_A_CY;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_A_XOR;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_B;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_B1;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_B2;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_B3;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_B4;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_B5;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_B6;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_BO5;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_BO6;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_B_CY;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_B_XOR;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_C;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_C1;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_C2;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_C3;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_C4;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_C5;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_C6;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_CLK;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_CO5;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_CO6;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_C_CY;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_C_XOR;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_D;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_D1;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_D2;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_D3;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_D4;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_D5;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_D6;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_DO5;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_DO6;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_D_CY;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X82Y119_D_XOR;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_A;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_A1;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_A2;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_A3;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_A4;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_A5;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_A6;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_AO5;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_AO6;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_A_CY;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_A_XOR;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_B;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_B1;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_B2;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_B3;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_B4;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_B5;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_B6;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_BO5;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_BO6;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_B_CY;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_B_XOR;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_C;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_C1;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_C2;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_C3;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_C4;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_C5;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_C6;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_CO5;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_CO6;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_C_CY;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_C_XOR;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_D;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_D1;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_D2;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_D3;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_D4;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_D5;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_D6;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_DO5;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_DO6;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_D_CY;
  wire [0:0] CLBLL_L_X54Y119_SLICE_X83Y119_D_XOR;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_A;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_A1;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_A2;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_A3;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_A4;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_A5;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_A6;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_AO5;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_AO6;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_AQ;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_AX;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_A_CY;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_A_XOR;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_B;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_B1;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_B2;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_B3;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_B4;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_B5;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_B6;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_BO5;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_BO6;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_B_CY;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_B_XOR;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_C;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_C1;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_C2;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_C3;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_C4;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_C5;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_C6;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_CLK;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_CO5;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_CO6;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_C_CY;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_C_XOR;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_D;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_D1;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_D2;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_D3;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_D4;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_D5;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_D6;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_DO5;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_DO6;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_D_CY;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X82Y123_D_XOR;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_A;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_A1;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_A2;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_A3;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_A4;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_A5;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_A6;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_AO5;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_AO6;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_A_CY;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_A_XOR;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_B;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_B1;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_B2;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_B3;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_B4;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_B5;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_B6;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_BO5;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_BO6;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_B_CY;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_B_XOR;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_C;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_C1;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_C2;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_C3;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_C4;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_C5;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_C6;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_CO5;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_CO6;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_C_CY;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_C_XOR;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_D;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_D1;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_D2;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_D3;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_D4;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_D5;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_D6;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_DO5;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_DO6;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_D_CY;
  wire [0:0] CLBLL_L_X54Y123_SLICE_X83Y123_D_XOR;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_A;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_A1;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_A2;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_A3;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_A4;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_A5;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_A6;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_AO5;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_AO6;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_AQ;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_AX;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_A_CY;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_A_XOR;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_B;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_B1;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_B2;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_B3;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_B4;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_B5;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_B6;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_BO5;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_BO6;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_B_CY;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_B_XOR;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_C;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_C1;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_C2;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_C3;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_C4;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_C5;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_C6;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_CLK;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_CO5;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_CO6;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_C_CY;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_C_XOR;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_D;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_D1;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_D2;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_D3;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_D4;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_D5;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_D6;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_DO5;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_DO6;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_D_CY;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X82Y133_D_XOR;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_A;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_A1;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_A2;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_A3;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_A4;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_A5;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_A6;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_AO5;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_AO6;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_A_CY;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_A_XOR;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_B;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_B1;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_B2;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_B3;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_B4;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_B5;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_B6;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_BO5;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_BO6;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_B_CY;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_B_XOR;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_C;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_C1;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_C2;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_C3;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_C4;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_C5;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_C6;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_CO5;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_CO6;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_C_CY;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_C_XOR;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_D;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_D1;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_D2;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_D3;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_D4;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_D5;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_D6;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_DO5;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_DO6;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_D_CY;
  wire [0:0] CLBLL_L_X54Y133_SLICE_X83Y133_D_XOR;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_A;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_A1;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_A2;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_A3;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_A4;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_A5;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_A6;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_AO5;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_AO6;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_AQ;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_AX;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_A_CY;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_A_XOR;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_B;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_B1;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_B2;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_B3;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_B4;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_B5;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_B6;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_BO5;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_BO6;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_B_CY;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_B_XOR;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_C;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_C1;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_C2;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_C3;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_C4;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_C5;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_C6;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_CLK;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_CO5;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_CO6;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_C_CY;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_C_XOR;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_D;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_D1;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_D2;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_D3;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_D4;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_D5;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_D6;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_DO5;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_DO6;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_D_CY;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X82Y138_D_XOR;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_A;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_A1;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_A2;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_A3;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_A4;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_A5;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_A6;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_AO5;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_AO6;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_A_CY;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_A_XOR;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_B;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_B1;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_B2;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_B3;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_B4;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_B5;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_B6;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_BO5;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_BO6;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_B_CY;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_B_XOR;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_C;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_C1;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_C2;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_C3;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_C4;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_C5;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_C6;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_CO5;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_CO6;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_C_CY;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_C_XOR;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_D;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_D1;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_D2;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_D3;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_D4;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_D5;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_D6;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_DO5;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_DO6;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_D_CY;
  wire [0:0] CLBLL_L_X54Y138_SLICE_X83Y138_D_XOR;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_A;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_A1;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_A2;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_A3;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_A4;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_A5;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_A6;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_AO5;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_AO6;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_AQ;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_AX;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_A_CY;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_A_XOR;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_B;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_B1;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_B2;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_B3;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_B4;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_B5;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_B6;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_BO5;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_BO6;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_B_CY;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_B_XOR;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_C;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_C1;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_C2;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_C3;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_C4;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_C5;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_C6;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_CLK;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_CO5;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_CO6;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_C_CY;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_C_XOR;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_D;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_D1;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_D2;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_D3;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_D4;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_D5;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_D6;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_DO5;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_DO6;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_D_CY;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X82Y141_D_XOR;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_A;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_A1;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_A2;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_A3;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_A4;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_A5;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_A6;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_AO5;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_AO6;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_A_CY;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_A_XOR;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_B;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_B1;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_B2;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_B3;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_B4;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_B5;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_B6;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_BO5;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_BO6;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_B_CY;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_B_XOR;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_C;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_C1;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_C2;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_C3;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_C4;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_C5;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_C6;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_CO5;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_CO6;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_C_CY;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_C_XOR;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_D;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_D1;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_D2;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_D3;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_D4;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_D5;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_D6;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_DO5;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_DO6;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_D_CY;
  wire [0:0] CLBLL_L_X54Y141_SLICE_X83Y141_D_XOR;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_A;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_A1;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_A2;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_A3;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_A4;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_A5;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_A6;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_AO5;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_AO6;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_AQ;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_AX;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_A_CY;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_A_XOR;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_B;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_B1;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_B2;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_B3;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_B4;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_B5;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_B6;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_BO5;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_BO6;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_B_CY;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_B_XOR;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_C;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_C1;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_C2;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_C3;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_C4;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_C5;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_C6;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_CLK;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_CO5;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_CO6;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_C_CY;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_C_XOR;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_D;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_D1;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_D2;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_D3;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_D4;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_D5;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_D6;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_DO5;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_DO6;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_D_CY;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X82Y96_D_XOR;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_A;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_A1;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_A2;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_A3;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_A4;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_A5;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_A6;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_AO5;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_AO6;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_A_CY;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_A_XOR;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_B;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_B1;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_B2;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_B3;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_B4;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_B5;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_B6;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_BO5;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_BO6;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_B_CY;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_B_XOR;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_C;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_C1;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_C2;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_C3;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_C4;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_C5;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_C6;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_CO5;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_CO6;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_C_CY;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_C_XOR;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_D;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_D1;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_D2;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_D3;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_D4;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_D5;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_D6;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_DO5;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_DO6;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_D_CY;
  wire [0:0] CLBLL_L_X54Y96_SLICE_X83Y96_D_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_AO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_AO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_BO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_BO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_BQ;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_CLK;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_CO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_CO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_DO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_DO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_AO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_AO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_BO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_BO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_CO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_CO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_DO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_DO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_AO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_AO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_AQ;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_BO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_BO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_CLK;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_CO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_CO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_DO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_DO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_AO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_AO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_AQ;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_BO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_BO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_CLK;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_CO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_CO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_DO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_DO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_AO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_AO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_AQ;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_BO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_BO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_BQ;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_CLK;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_CO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_CO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_CQ;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_DO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_DQ;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_AO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_AO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_BO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_BO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_CO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_CO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_DO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_DO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_AO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_AO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_BO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_BO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_CO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_CO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_DO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_DO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_AO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_AO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_AQ;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_BO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_BO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_BQ;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_CLK;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_CO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_CO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_CQ;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_DO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_AO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_AO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_BO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_BO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_CO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_CO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_DO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_DO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_AO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_AO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_BO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_BO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_CO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_CO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_DO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_DO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A5Q;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_AMUX;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_AO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_AO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_AQ;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_BO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_BO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_CLK;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_CO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_CO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_DO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_AO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_AO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_BO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_BO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_CO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_CO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_DO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_AO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_AO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_BO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_BO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_CO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_CO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_DO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_DO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_AMUX;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_AO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_AO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_BMUX;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_BO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_BO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_CO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_CO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_DO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_DO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_AMUX;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_AO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_AO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_BO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_BO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_CO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_CO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_DO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_DO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_AO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_AO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_BO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_BO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_CO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_CO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_DO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_DO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_AO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_AO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_AX;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_BO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_BO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_CLK;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_CO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_CO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_DO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_DO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_AO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_AO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_BO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_BO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_CO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_CO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_DO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_DO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_AO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_AO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_BO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_BO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_CLK;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_CO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_CO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_DO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_DO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_AO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_AO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_BO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_BO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_CO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_CO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_DO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_DO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_AO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_AO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_AQ;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_BO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_BO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_BQ;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_CLK;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_CO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_CO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_CQ;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_DO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_DO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_AO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_AO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_BO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_BO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_CO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_CO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_DO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_DO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_AO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_AO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_BO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_BO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_CO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_CO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_DO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_DO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_AO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_AO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_BO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_BO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_CO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_CO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_DO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_DO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D_XOR;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_A;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_A1;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_A2;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_A3;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_A4;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_A5;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_A6;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_AO5;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_AO6;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_AQ;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_A_CY;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_A_XOR;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_B;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_B1;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_B2;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_B3;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_B4;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_B5;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_B6;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_BO5;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_BO6;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_BQ;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_B_CY;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_B_XOR;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_C;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_C1;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_C2;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_C3;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_C4;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_C5;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_C6;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_CLK;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_CO5;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_CO6;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_C_CY;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_C_XOR;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_D;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_D1;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_D2;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_D3;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_D4;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_D5;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_D6;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_DO5;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_DO6;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_D_CY;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_D_XOR;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_A;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_A1;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_A2;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_A3;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_A4;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_A5;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_A6;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_AO5;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_AO6;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_A_CY;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_A_XOR;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_B;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_B1;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_B2;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_B3;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_B4;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_B5;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_B6;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_BO5;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_BO6;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_B_CY;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_B_XOR;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_C;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_C1;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_C2;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_C3;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_C4;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_C5;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_C6;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_CO5;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_CO6;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_C_CY;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_C_XOR;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_D;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_D1;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_D2;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_D3;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_D4;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_D5;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_D6;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_DO5;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_DO6;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_D_CY;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_D_XOR;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_A;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_A1;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_A2;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_A3;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_A4;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_A5;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_A6;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_AO5;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_AO6;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_AQ;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_A_CY;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_A_XOR;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_B;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_B1;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_B2;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_B3;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_B4;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_B5;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_B6;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_BO5;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_BO6;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_B_CY;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_B_XOR;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_C;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_C1;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_C2;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_C3;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_C4;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_C5;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_C6;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_CLK;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_CO5;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_CO6;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_C_CY;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_C_XOR;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_D;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_D1;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_D2;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_D3;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_D4;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_D5;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_D6;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_DO5;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_DO6;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_D_CY;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_D_XOR;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_A;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_A1;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_A2;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_A3;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_A4;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_A5;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_A6;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_AO5;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_AO6;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_A_CY;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_A_XOR;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_B;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_B1;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_B2;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_B3;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_B4;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_B5;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_B6;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_BO5;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_BO6;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_B_CY;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_B_XOR;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_C;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_C1;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_C2;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_C3;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_C4;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_C5;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_C6;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_CO5;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_CO6;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_C_CY;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_C_XOR;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_D;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_D1;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_D2;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_D3;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_D4;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_D5;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_D6;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_DO5;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_DO6;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_D_CY;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_D_XOR;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_A;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_A1;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_A2;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_A3;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_A4;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_A5;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_A6;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_AO5;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_AO6;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_AQ;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_A_CY;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_A_XOR;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_B;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_B1;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_B2;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_B3;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_B4;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_B5;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_B6;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_BO5;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_BO6;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_BQ;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_B_CY;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_B_XOR;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_C;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_C1;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_C2;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_C3;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_C4;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_C5;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_C6;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_CLK;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_CO5;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_CO6;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_C_CY;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_C_XOR;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_D;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_D1;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_D2;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_D3;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_D4;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_D5;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_D6;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_DO5;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_DO6;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_D_CY;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_D_XOR;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_A;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_A1;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_A2;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_A3;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_A4;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_A5;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_A6;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_AO5;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_AO6;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_A_CY;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_A_XOR;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_B;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_B1;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_B2;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_B3;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_B4;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_B5;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_B6;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_BO5;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_BO6;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_B_CY;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_B_XOR;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_C;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_C1;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_C2;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_C3;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_C4;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_C5;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_C6;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_CO5;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_CO6;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_C_CY;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_C_XOR;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_D;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_D1;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_D2;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_D3;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_D4;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_D5;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_D6;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_DO5;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_DO6;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_D_CY;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_D_XOR;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_A;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_A1;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_A2;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_A3;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_A4;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_A5;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_A6;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_AO5;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_AO6;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_AQ;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_AX;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_A_CY;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_A_XOR;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_B;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_B1;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_B2;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_B3;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_B4;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_B5;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_B6;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_BO5;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_BO6;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_BQ;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_BX;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_B_CY;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_B_XOR;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_C;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_C1;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_C2;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_C3;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_C4;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_C5;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_C6;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_CE;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_CLK;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_CO5;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_CO6;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_C_CY;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_C_XOR;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_D;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_D1;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_D2;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_D3;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_D4;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_D5;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_D6;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_DO5;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_DO6;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_D_CY;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X22Y149_D_XOR;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_A;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_A1;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_A2;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_A3;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_A4;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_A5;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_A6;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_AO5;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_AO6;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_A_CY;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_A_XOR;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_B;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_B1;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_B2;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_B3;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_B4;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_B5;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_B6;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_BO5;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_BO6;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_B_CY;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_B_XOR;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_C;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_C1;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_C2;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_C3;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_C4;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_C5;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_C6;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_CO5;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_CO6;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_C_CY;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_C_XOR;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_D;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_D1;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_D2;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_D3;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_D4;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_D5;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_D6;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_DO5;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_DO6;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_D_CY;
  wire [0:0] CLBLM_L_X16Y149_SLICE_X23Y149_D_XOR;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_A;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_A1;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_A2;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_A3;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_A4;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_A5;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_A6;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_AO5;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_AO6;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_AQ;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_AX;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_A_CY;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_A_XOR;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_B;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_B1;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_B2;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_B3;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_B4;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_B5;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_B6;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_BO5;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_BO6;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_BQ;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_BX;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_B_CY;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_B_XOR;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_C;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_C1;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_C2;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_C3;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_C4;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_C5;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_C6;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_CE;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_CLK;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_CO5;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_CO6;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_CQ;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_CX;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_C_CY;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_C_XOR;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_D;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_D1;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_D2;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_D3;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_D4;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_D5;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_D6;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_DO5;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_DO6;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_DQ;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_DX;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_D_CY;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_D_XOR;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_A;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_A1;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_A2;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_A3;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_A4;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_A5;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_A6;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_AO5;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_AO6;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_AQ;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_AX;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_A_CY;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_A_XOR;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_B;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_B1;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_B2;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_B3;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_B4;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_B5;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_B6;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_BO5;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_BO6;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_B_CY;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_B_XOR;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_C;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_C1;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_C2;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_C3;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_C4;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_C5;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_C6;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_CE;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_CLK;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_CO5;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_CO6;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_C_CY;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_C_XOR;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_D;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_D1;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_D2;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_D3;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_D4;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_D5;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_D6;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_DO5;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_DO6;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_D_CY;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_D_XOR;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_A;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_A1;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_A2;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_A3;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_A4;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_A5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_A6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_AO5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_AO6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_AQ;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_AX;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_A_CY;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_A_XOR;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_B;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_B1;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_B2;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_B3;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_B4;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_B5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_B6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_BO5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_BO6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_BQ;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_BX;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_B_CY;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_B_XOR;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_C;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_C1;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_C2;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_C3;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_C4;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_C5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_C6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_CE;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_CLK;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_CO5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_CO6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_C_CY;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_C_XOR;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_D;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_D1;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_D2;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_D3;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_D4;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_D5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_D6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_DO5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_DO6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_D_CY;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_D_XOR;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_A;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_A1;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_A2;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_A3;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_A4;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_A5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_A6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_AO5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_AO6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_A_CY;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_A_XOR;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_B;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_B1;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_B2;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_B3;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_B4;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_B5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_B6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_BO5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_BO6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_B_CY;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_B_XOR;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_C;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_C1;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_C2;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_C3;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_C4;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_C5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_C6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_CO5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_CO6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_C_CY;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_C_XOR;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_D;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_D1;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_D2;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_D3;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_D4;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_D5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_D6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_DO5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_DO6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_D_CY;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_D_XOR;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_A;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_A1;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_A2;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_A3;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_A4;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_A5;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_A6;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_AO5;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_AO6;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_AQ;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_AX;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_A_CY;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_A_XOR;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_B;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_B1;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_B2;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_B3;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_B4;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_B5;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_B6;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_BO5;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_BO6;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_B_CY;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_B_XOR;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_C;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_C1;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_C2;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_C3;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_C4;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_C5;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_C6;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_CE;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_CLK;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_CO5;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_CO6;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_C_CY;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_C_XOR;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_D;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_D1;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_D2;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_D3;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_D4;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_D5;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_D6;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_DO5;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_DO6;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_D_CY;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_D_XOR;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_A;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_A1;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_A2;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_A3;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_A4;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_A5;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_A6;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_AO5;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_AO6;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_A_CY;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_A_XOR;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_B;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_B1;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_B2;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_B3;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_B4;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_B5;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_B6;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_BO5;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_BO6;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_B_CY;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_B_XOR;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_C;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_C1;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_C2;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_C3;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_C4;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_C5;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_C6;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_CO5;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_CO6;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_C_CY;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_C_XOR;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_D;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_D1;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_D2;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_D3;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_D4;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_D5;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_D6;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_DO5;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_DO6;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_D_CY;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_D_XOR;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_A;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_A1;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_A2;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_A3;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_A4;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_A5;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_A6;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_AO5;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_AO6;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_AQ;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_AX;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_A_CY;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_A_XOR;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_B;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_B1;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_B2;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_B3;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_B4;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_B5;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_B6;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_BO5;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_BO6;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_BQ;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_BX;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_B_CY;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_B_XOR;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_C;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_C1;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_C2;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_C3;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_C4;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_C5;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_C6;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_CE;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_CLK;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_CO5;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_CO6;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_C_CY;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_C_XOR;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_D;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_D1;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_D2;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_D3;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_D4;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_D5;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_D6;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_DO5;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_DO6;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_D_CY;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_D_XOR;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_A;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_A1;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_A2;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_A3;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_A4;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_A5;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_A6;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_AO5;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_AO6;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_A_CY;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_A_XOR;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_B;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_B1;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_B2;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_B3;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_B4;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_B5;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_B6;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_BO5;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_BO6;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_B_CY;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_B_XOR;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_C;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_C1;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_C2;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_C3;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_C4;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_C5;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_C6;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_CO5;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_CO6;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_C_CY;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_C_XOR;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_D;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_D1;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_D2;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_D3;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_D4;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_D5;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_D6;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_DO5;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_DO6;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_D_CY;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_D_XOR;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_A;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_A1;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_A2;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_A3;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_A4;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_A5;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_A6;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_AO5;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_AO6;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_AQ;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_AX;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_A_CY;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_A_XOR;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_B;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_B1;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_B2;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_B3;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_B4;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_B5;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_B6;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_BO5;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_BO6;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_B_CY;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_B_XOR;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_C;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_C1;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_C2;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_C3;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_C4;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_C5;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_C6;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_CE;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_CLK;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_CO5;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_CO6;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_C_CY;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_C_XOR;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_D;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_D1;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_D2;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_D3;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_D4;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_D5;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_D6;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_DO5;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_DO6;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_D_CY;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X22Y155_D_XOR;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_A;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_A1;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_A2;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_A3;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_A4;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_A5;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_A6;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_AO5;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_AO6;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_A_CY;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_A_XOR;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_B;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_B1;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_B2;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_B3;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_B4;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_B5;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_B6;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_BO5;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_BO6;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_B_CY;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_B_XOR;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_C;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_C1;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_C2;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_C3;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_C4;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_C5;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_C6;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_CO5;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_CO6;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_C_CY;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_C_XOR;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_D;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_D1;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_D2;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_D3;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_D4;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_D5;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_D6;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_DO5;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_DO6;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_D_CY;
  wire [0:0] CLBLM_L_X16Y155_SLICE_X23Y155_D_XOR;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_A;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_A1;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_A2;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_A3;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_A4;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_A5;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_A6;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_AO5;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_AO6;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_AQ;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_AX;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_A_CY;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_A_XOR;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_B;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_B1;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_B2;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_B3;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_B4;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_B5;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_B6;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_BO5;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_BO6;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_B_CY;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_B_XOR;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_C;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_C1;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_C2;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_C3;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_C4;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_C5;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_C6;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_CE;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_CLK;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_CO5;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_CO6;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_C_CY;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_C_XOR;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_D;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_D1;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_D2;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_D3;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_D4;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_D5;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_D6;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_DO5;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_DO6;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_D_CY;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X22Y157_D_XOR;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_A;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_A1;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_A2;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_A3;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_A4;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_A5;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_A6;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_AO5;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_AO6;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_A_CY;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_A_XOR;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_B;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_B1;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_B2;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_B3;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_B4;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_B5;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_B6;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_BO5;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_BO6;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_B_CY;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_B_XOR;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_C;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_C1;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_C2;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_C3;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_C4;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_C5;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_C6;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_CO5;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_CO6;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_C_CY;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_C_XOR;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_D;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_D1;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_D2;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_D3;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_D4;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_D5;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_D6;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_DO5;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_DO6;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_D_CY;
  wire [0:0] CLBLM_L_X16Y157_SLICE_X23Y157_D_XOR;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_A;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_A1;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_A2;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_A3;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_A4;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_A5;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_A6;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_AO5;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_AO6;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_AQ;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_AX;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_A_CY;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_A_XOR;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_B;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_B1;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_B2;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_B3;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_B4;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_B5;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_B6;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_BO5;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_BO6;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_B_CY;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_B_XOR;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_C;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_C1;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_C2;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_C3;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_C4;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_C5;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_C6;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_CLK;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_CO5;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_CO6;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_C_CY;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_C_XOR;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_D;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_D1;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_D2;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_D3;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_D4;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_D5;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_D6;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_DO5;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_DO6;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_D_CY;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X84Y151_D_XOR;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_A;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_A1;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_A2;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_A3;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_A4;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_A5;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_A6;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_AO5;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_AO6;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_A_CY;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_A_XOR;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_B;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_B1;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_B2;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_B3;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_B4;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_B5;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_B6;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_BO5;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_BO6;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_B_CY;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_B_XOR;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_C;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_C1;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_C2;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_C3;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_C4;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_C5;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_C6;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_CO5;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_CO6;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_C_CY;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_C_XOR;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_D;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_D1;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_D2;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_D3;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_D4;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_D5;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_D6;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_DO5;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_DO6;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_D_CY;
  wire [0:0] CLBLM_L_X56Y151_SLICE_X85Y151_D_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_AO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_AO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_AQ;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_BO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_BO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_BQ;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_CLK;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_CO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_CO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_DO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_DO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_AO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_AO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_BO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_BO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_CO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_CO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_DO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_DO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_AO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_AO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_BO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_BO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_BQ;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_CLK;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_CO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_CO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_CQ;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_DO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_DO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_AO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_AO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_BO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_BO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_CO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_CO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_DO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_DO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A5Q;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_AMUX;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_AO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_AO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B5Q;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_BMUX;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_BO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_BO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_BQ;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_CLK;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_CO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_CO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_CQ;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_DO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_DO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_DQ;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_AMUX;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_AO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_AO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_BO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_BO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_BQ;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_CLK;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_CO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_CO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_CQ;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_DO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_DO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_DQ;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_AO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_AO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_BO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_BO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_BQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_CLK;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_CO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_CO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_DO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_DO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_AO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_AO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_BO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_BO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_BQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_CLK;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_CO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_CO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_CQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_DO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_AO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_AO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_BO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_BO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_CO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_CO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_DO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_DO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A5Q;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_AMUX;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_AO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_AO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_AQ;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_BO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_BO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_BQ;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_CLK;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_CO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_CO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_CQ;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_DO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_DO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_AO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_AO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_BO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_BO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_CO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_CO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_DO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_DO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_AMUX;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_AO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_AO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_BO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_BO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_CO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_CO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_DO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_DO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_AO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_AO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_AQ;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_BO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_BO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_CLK;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_CO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_CO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_DO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_DO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_AO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_AO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_BO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_BO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_CO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_CO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_DO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_DO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A5Q;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_AMUX;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_AO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_AO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_AQ;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_BMUX;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_BO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_BO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_CLK;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_CMUX;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_CO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_CO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_DO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_DO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_AO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_AO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_BO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_BO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_CO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_CO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_DO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_DO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A5Q;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_AMUX;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_AO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_AO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_AQ;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_BMUX;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_BO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_BO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_CLK;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_CO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_CO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_DO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_DO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_AO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_AO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_BO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_BO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_CO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_CO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_DO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_DO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A5Q;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_AMUX;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_AO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_AO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_AQ;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B5Q;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_BMUX;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_BO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_BO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_BQ;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_CLK;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_CO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_CO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_DO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_DO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_AO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_AO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_BO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_BO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_CO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_CO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_DO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_DO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_AO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_BO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_CLK;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_CO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_CO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_DO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_AO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_AO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_BO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_BO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_CO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_CO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_DO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_DO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_AO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_AO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_AQ;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_BO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_BO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_CLK;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_CO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_CO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_DO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_DO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_AO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_AO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_BO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_BO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_CO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_CO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_DO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_DO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_AO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_AO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_AQ;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_BO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_BO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_BQ;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_CLK;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_CO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_DO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_DO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_AO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_AO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_BO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_BO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_CO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_CO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_DO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_DO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_AO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_AO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_AQ;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_BO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_BO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_BQ;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_CLK;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_CO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_CO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_DO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_DO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_AO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_AO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_BO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_BO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_CO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_CO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_DO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_DO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_AO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_AO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_BO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_BO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_CO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_CO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_DO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_DO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_AO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_AO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_BO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_BO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_CO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_CO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_DO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_DO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_AO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_AO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_BO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_BO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_CO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_CO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_DO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_DO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_AO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_AO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_BO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_BO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_CO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_CO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_DO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_DO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D_XOR;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_A;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_A1;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_A2;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_A3;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_A4;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_A5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_A6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_AMUX;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_AO5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_AO6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_A_CY;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_A_XOR;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_B;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_B1;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_B2;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_B3;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_B4;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_B5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_B6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_BO5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_BO6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_B_CY;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_B_XOR;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_C;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_C1;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_C2;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_C3;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_C4;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_C5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_C6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_CO5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_CO6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_C_CY;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_C_XOR;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_D;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_D1;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_D2;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_D3;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_D4;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_D5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_D6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_DO5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_DO6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_D_CY;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_D_XOR;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_A;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_A1;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_A2;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_A3;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_A4;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_A5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_A6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_AO5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_AO6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_A_CY;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_A_XOR;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_B;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_B1;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_B2;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_B3;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_B4;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_B5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_B6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_BO5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_BO6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_B_CY;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_B_XOR;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_C;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_C1;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_C2;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_C3;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_C4;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_C5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_C6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_CO5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_CO6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_C_CY;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_C_XOR;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_D;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_D1;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_D2;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_D3;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_D4;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_D5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_D6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_DO5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_DO6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_D_CY;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_D_XOR;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_A;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_A1;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_A2;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_A3;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_A4;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_A5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_A6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_AO5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_AO6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_AQ;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_A_CY;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_A_XOR;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_B;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_B1;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_B2;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_B3;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_B4;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_B5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_B6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_BO5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_BO6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_B_CY;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_B_XOR;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_C;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_C1;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_C2;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_C3;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_C4;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_C5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_C6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_CLK;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_CO5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_CO6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_C_CY;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_C_XOR;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_D;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_D1;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_D2;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_D3;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_D4;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_D5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_D6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_DO5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_DO6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_D_CY;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_D_XOR;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_A;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_A1;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_A2;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_A3;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_A4;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_A5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_A6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_AO5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_AO6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_A_CY;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_A_XOR;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_B;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_B1;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_B2;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_B3;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_B4;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_B5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_B6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_BO5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_BO6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_B_CY;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_B_XOR;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_C;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_C1;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_C2;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_C3;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_C4;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_C5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_C6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_CO5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_CO6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_C_CY;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_C_XOR;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_D;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_D1;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_D2;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_D3;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_D4;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_D5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_D6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_DO5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_DO6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_D_CY;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_D_XOR;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_A;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_A1;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_A2;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_A3;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_A4;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_A5;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_A6;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_AO5;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_AO6;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_A_CY;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_A_XOR;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_B;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_B1;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_B2;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_B3;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_B4;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_B5;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_B6;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_BO5;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_BO6;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_B_CY;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_B_XOR;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_C;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_C1;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_C2;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_C3;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_C4;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_C5;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_C6;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_CO5;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_CO6;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_C_CY;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_C_XOR;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_D;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_D1;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_D2;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_D3;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_D4;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_D5;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_D6;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_DO5;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_DO6;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_D_CY;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_D_XOR;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_A;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_A1;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_A2;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_A3;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_A4;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_A5;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_A6;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_AO5;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_AO6;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_AQ;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_A_CY;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_A_XOR;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_B;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_B1;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_B2;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_B3;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_B4;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_B5;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_B6;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_BO5;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_BO6;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_B_CY;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_B_XOR;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_C;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_C1;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_C2;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_C3;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_C4;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_C5;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_C6;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_CLK;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_CO5;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_CO6;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_C_CY;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_C_XOR;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_D;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_D1;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_D2;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_D3;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_D4;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_D5;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_D6;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_DO5;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_DO6;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_D_CY;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_D_XOR;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_A;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_A1;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_A2;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_A3;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_A4;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_A5;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_A6;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_AO5;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_AO6;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_AQ;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_AX;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_A_CY;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_A_XOR;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_B;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_B1;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_B2;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_B3;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_B4;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_B5;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_B6;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_BO5;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_BO6;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_BQ;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_BX;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_B_CY;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_B_XOR;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_C;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_C1;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_C2;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_C3;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_C4;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_C5;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_C6;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_CE;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_CLK;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_CO5;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_CO6;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_C_CY;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_C_XOR;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_D;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_D1;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_D2;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_D3;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_D4;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_D5;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_D6;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_DO5;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_DO6;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_D_CY;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X36Y149_D_XOR;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_A;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_A1;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_A2;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_A3;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_A4;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_A5;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_A6;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_AO5;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_AO6;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_AQ;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_AX;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_A_CY;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_A_XOR;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_B;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_B1;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_B2;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_B3;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_B4;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_B5;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_B6;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_BO5;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_BO6;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_B_CY;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_B_XOR;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_C;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_C1;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_C2;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_C3;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_C4;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_C5;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_C6;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_CE;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_CLK;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_CO5;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_CO6;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_C_CY;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_C_XOR;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_D;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_D1;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_D2;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_D3;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_D4;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_D5;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_D6;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_DO5;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_DO6;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_D_CY;
  wire [0:0] CLBLM_R_X25Y149_SLICE_X37Y149_D_XOR;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_A;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_A1;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_A2;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_A3;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_A4;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_A5;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_A6;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_AO5;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_AO6;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_AQ;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_AX;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_A_CY;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_A_XOR;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_B;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_B1;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_B2;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_B3;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_B4;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_B5;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_B6;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_BO5;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_BO6;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_BQ;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_BX;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_B_CY;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_B_XOR;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_C;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_C1;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_C2;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_C3;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_C4;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_C5;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_C6;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_CE;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_CLK;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_CO5;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_CO6;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_CQ;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_CX;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_C_CY;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_C_XOR;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_D;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_D1;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_D2;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_D3;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_D4;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_D5;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_D6;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_DO5;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_DO6;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_D_CY;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X36Y151_D_XOR;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_A;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_A1;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_A2;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_A3;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_A4;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_A5;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_A6;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_AO5;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_AO6;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_A_CY;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_A_XOR;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_B;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_B1;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_B2;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_B3;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_B4;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_B5;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_B6;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_BO5;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_BO6;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_B_CY;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_B_XOR;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_C;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_C1;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_C2;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_C3;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_C4;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_C5;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_C6;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_CO5;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_CO6;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_C_CY;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_C_XOR;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_D;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_D1;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_D2;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_D3;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_D4;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_D5;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_D6;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_DO5;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_DO6;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_D_CY;
  wire [0:0] CLBLM_R_X25Y151_SLICE_X37Y151_D_XOR;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_A;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_A1;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_A2;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_A3;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_A4;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_A5;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_A6;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_AO5;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_AO6;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_AQ;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_AX;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_A_CY;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_A_XOR;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_B;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_B1;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_B2;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_B3;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_B4;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_B5;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_B6;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_BO5;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_BO6;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_BQ;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_BX;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_B_CY;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_B_XOR;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_C;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_C1;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_C2;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_C3;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_C4;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_C5;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_C6;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_CE;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_CLK;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_CO5;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_CO6;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_C_CY;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_C_XOR;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_D;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_D1;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_D2;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_D3;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_D4;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_D5;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_D6;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_DO5;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_DO6;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_D_CY;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X36Y153_D_XOR;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_A;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_A1;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_A2;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_A3;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_A4;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_A5;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_A6;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_AO5;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_AO6;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_A_CY;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_A_XOR;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_B;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_B1;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_B2;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_B3;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_B4;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_B5;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_B6;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_BO5;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_BO6;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_B_CY;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_B_XOR;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_C;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_C1;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_C2;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_C3;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_C4;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_C5;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_C6;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_CO5;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_CO6;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_C_CY;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_C_XOR;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_D;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_D1;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_D2;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_D3;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_D4;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_D5;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_D6;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_DO5;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_DO6;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_D_CY;
  wire [0:0] CLBLM_R_X25Y153_SLICE_X37Y153_D_XOR;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_A;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_A1;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_A2;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_A3;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_A4;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_A5;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_A6;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_AO5;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_AO6;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_AQ;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_AX;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_A_CY;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_A_XOR;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_B;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_B1;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_B2;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_B3;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_B4;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_B5;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_B6;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_BO5;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_BO6;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_BQ;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_BX;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_B_CY;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_B_XOR;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_C;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_C1;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_C2;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_C3;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_C4;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_C5;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_C6;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_CE;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_CLK;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_CO5;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_CO6;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_CQ;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_CX;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_C_CY;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_C_XOR;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_D;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_D1;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_D2;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_D3;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_D4;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_D5;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_D6;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_DO5;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_DO6;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_D_CY;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X36Y154_D_XOR;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_A;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_A1;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_A2;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_A3;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_A4;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_A5;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_A6;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_AO5;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_AO6;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_A_CY;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_A_XOR;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_B;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_B1;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_B2;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_B3;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_B4;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_B5;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_B6;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_BO5;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_BO6;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_B_CY;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_B_XOR;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_C;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_C1;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_C2;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_C3;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_C4;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_C5;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_C6;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_CO5;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_CO6;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_C_CY;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_C_XOR;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_D;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_D1;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_D2;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_D3;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_D4;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_D5;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_D6;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_DO5;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_DO6;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_D_CY;
  wire [0:0] CLBLM_R_X25Y154_SLICE_X37Y154_D_XOR;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_A;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_A1;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_A2;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_A3;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_A4;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_A5;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_A6;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_AO5;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_AO6;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_AQ;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_AX;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_A_CY;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_A_XOR;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_B;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_B1;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_B2;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_B3;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_B4;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_B5;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_B6;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_BO5;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_BO6;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_BQ;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_BX;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_B_CY;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_B_XOR;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_C;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_C1;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_C2;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_C3;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_C4;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_C5;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_C6;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_CE;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_CLK;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_CO5;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_CO6;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_C_CY;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_C_XOR;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_D;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_D1;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_D2;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_D3;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_D4;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_D5;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_D6;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_DO5;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_DO6;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_D_CY;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X36Y157_D_XOR;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_A;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_A1;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_A2;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_A3;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_A4;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_A5;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_A6;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_AO5;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_AO6;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_AQ;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_AX;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_A_CY;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_A_XOR;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_B;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_B1;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_B2;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_B3;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_B4;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_B5;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_B6;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_BO5;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_BO6;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_B_CY;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_B_XOR;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_C;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_C1;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_C2;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_C3;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_C4;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_C5;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_C6;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_CE;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_CLK;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_CO5;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_CO6;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_C_CY;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_C_XOR;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_D;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_D1;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_D2;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_D3;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_D4;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_D5;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_D6;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_DO5;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_DO6;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_D_CY;
  wire [0:0] CLBLM_R_X25Y157_SLICE_X37Y157_D_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A5Q;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_AMUX;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_AO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_AO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_AQ;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_BO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_BO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_BQ;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_CLK;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_CO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_CO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_DO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_DO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_SR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_AO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_AO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_BO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_BO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_CO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_CO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_DO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_AO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_AO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_AQ;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_BO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_BO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_CLK;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_CO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_CO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_DO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_DO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_AMUX;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_AO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_AO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_AQ;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_BO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_BO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_BQ;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_CLK;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_CO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_CO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_DO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_DO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A5Q;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_AMUX;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_AO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_AO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_AQ;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B5Q;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_BMUX;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_BO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_BO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_BQ;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C5Q;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_CLK;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_CMUX;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_CO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_CO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_CQ;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_DMUX;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_DO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_DO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_SR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_AMUX;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_AO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_AO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_AQ;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_AX;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B5Q;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_BMUX;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_BO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_BO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_BQ;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_BX;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_CLK;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_CO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_CO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_CQ;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_DO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_DO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_DQ;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_AMUX;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_AO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_AO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_AQ;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_BMUX;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_BO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_BO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_BQ;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_CLK;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_CO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_CO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_CQ;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_DO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_DO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_DQ;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_AMUX;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_AO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_AO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_AQ;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_BO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_BO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_BQ;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_CLK;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_CO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_CO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_CQ;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_DO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_DO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_AO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_AO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_BO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_BO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_CO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_CO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_DO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_DO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_AMUX;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_AO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_AO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_AQ;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_BO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_BO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_BQ;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_CLK;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_CO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_CO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_DO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_DO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D_XOR;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_A;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_A1;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_A2;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_A3;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_A4;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_A5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_A6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_AMUX;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_AO5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_AO6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_AQ;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_A_CY;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_A_XOR;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_B;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_B1;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_B2;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_B3;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_B4;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_B5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_B6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_BO5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_BO6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_BQ;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_B_CY;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_B_XOR;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_C;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_C1;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_C2;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_C3;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_C4;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_C5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_C6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_CLK;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_CO5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_CO6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_C_CY;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_C_XOR;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_D;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_D1;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_D2;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_D3;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_D4;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_D5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_D6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_DO5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_DO6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_D_CY;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_D_XOR;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_A;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_A1;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_A2;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_A3;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_A4;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_A5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_A6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_AMUX;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_AO5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_AO6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_A_CY;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_A_XOR;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_B;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_B1;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_B2;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_B3;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_B4;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_B5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_B6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_BO5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_BO6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_B_CY;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_B_XOR;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_C;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_C1;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_C2;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_C3;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_C4;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_C5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_C6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_CO5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_CO6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_C_CY;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_C_XOR;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_D;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_D1;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_D2;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_D3;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_D4;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_D5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_D6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_DO5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_DO6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_D_CY;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_D_XOR;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_A;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_A1;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_A2;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_A3;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_A4;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_A5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_A6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_AO5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_AO6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_A_CY;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_A_XOR;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_B;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_B1;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_B2;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_B3;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_B4;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_B5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_B6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_BO5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_BO6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_B_CY;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_B_XOR;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_C;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_C1;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_C2;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_C3;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_C4;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_C5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_C6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_CO5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_CO6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_C_CY;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_C_XOR;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_D;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_D1;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_D2;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_D3;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_D4;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_D5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_D6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_DO5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_DO6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_D_CY;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_D_XOR;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_A;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_A1;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_A2;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_A3;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_A4;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_A5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_A6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_AMUX;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_AO5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_AO6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_A_CY;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_A_XOR;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_B;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_B1;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_B2;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_B3;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_B4;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_B5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_B6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_BMUX;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_BO5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_BO6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_B_CY;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_B_XOR;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_C;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_C1;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_C2;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_C3;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_C4;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_C5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_C6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_CO5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_CO6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_C_CY;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_C_XOR;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_D;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_D1;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_D2;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_D3;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_D4;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_D5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_D6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_DO5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_DO6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_D_CY;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_D_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_AO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_AO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_BO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_BO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_CO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_CO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_DO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_DO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_AMUX;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_AO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_AO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_BO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_BO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_CO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_CO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_DO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_DO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_AO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_AO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_BO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_BO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_CO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_CO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_DO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_DO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_AO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_AO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_BO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_BO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_CO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_CO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_DO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_DO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_AO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_AO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_BO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_BO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_CO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_CO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_DO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_DO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_AO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_AO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_BO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_BO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_CO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_CO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_DO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_DO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_AO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_AO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_AQ;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_AX;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_BO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_BO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_BQ;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_BX;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_CE;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_CLK;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_CO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_CO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_CQ;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_CX;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_DO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_DO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_AO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_AO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_BO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_BO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_CO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_CO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_DO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_DO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_AO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_AQ;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_AX;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_BO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_BO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_BQ;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_BX;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_CE;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_CLK;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_CO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_CO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_CQ;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_CX;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_DO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_DO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_DQ;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_DX;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_AO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_AO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_BO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_BO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_CO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_CO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_DO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_DO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_AO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_AO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_AX;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_BO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_BO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_BQ;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_BX;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_CE;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_CLK;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_CO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_CO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_CQ;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_CX;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_DO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_DO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_DQ;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_DX;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_AO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_AO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_AQ;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_AX;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_BO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_BO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_BQ;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_BX;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_CE;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_CLK;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_CO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_CO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_DO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_DO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_AO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_AO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_AQ;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_AX;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_BO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_BO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_BQ;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_BX;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_CE;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_CLK;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_CO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_CO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_CQ;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_CX;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_DO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_DO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_DQ;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_DX;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_AO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_AQ;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_AX;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_BO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_BO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_BQ;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_BX;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_CE;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_CLK;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_CO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_CO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_CQ;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_CX;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_DO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_DO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_DQ;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_DX;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_AO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_AO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_AQ;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_AX;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_BO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_BO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_BQ;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_BX;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_CE;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_CLK;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_CO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_CO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_CQ;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_CX;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_DO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_DQ;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_DX;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_AO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_AO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_AQ;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_AX;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_BO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_BO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_CE;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_CLK;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_CO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_CO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_DO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_AO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_AO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_AQ;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_AX;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_BO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_BO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_BQ;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_BX;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_CE;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_CLK;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_CO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_CO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_CQ;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_CX;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_DO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_DO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_DQ;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_DX;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_AO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_AO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_AQ;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_AX;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_BO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_BO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_BX;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_CE;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_CLK;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_CO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_CO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_DO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_DO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_AO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_AO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_AQ;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_AX;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_BO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_BO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_BQ;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_BX;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_CE;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_CLK;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_CO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_CO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_CQ;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_CX;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_DO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_DO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_DQ;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_DX;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_AO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_AO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_AQ;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_AX;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_BO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_BO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_BQ;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_BX;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_CE;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_CLK;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_CO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_CO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_CQ;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_CX;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_DO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_DO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_DQ;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_DX;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D_XOR;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_A;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_A1;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_A2;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_A3;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_A4;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_A5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_A6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_AO5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_AO6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_AQ;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_AX;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_A_CY;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_A_XOR;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_B;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_B1;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_B2;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_B3;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_B4;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_B5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_B6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_BO5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_BO6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_BQ;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_BX;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_B_CY;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_B_XOR;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_C;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_C1;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_C2;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_C3;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_C4;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_C5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_C6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_CE;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_CLK;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_CO5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_CO6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_CQ;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_CX;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_C_CY;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_C_XOR;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_D;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_D1;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_D2;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_D3;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_D4;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_D5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_D6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_DO5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_DO6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_DQ;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_DX;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_D_CY;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_D_XOR;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_A;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_A1;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_A2;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_A3;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_A4;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_A5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_A6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_AO5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_AO6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_AQ;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_AX;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_A_CY;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_A_XOR;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_B;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_B1;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_B2;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_B3;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_B4;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_B5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_B6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_BO5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_BO6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_BQ;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_BX;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_B_CY;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_B_XOR;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_C;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_C1;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_C2;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_C3;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_C4;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_C5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_C6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_CE;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_CLK;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_CO5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_CO6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_CQ;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_CX;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_C_CY;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_C_XOR;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_D;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_D1;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_D2;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_D3;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_D4;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_D5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_D6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_DO5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_DO6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_D_CY;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_D_XOR;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_A;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_A1;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_A2;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_A3;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_A4;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_A5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_A6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_AO5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_AO6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_AQ;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_AX;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_A_CY;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_A_XOR;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_B;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_B1;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_B2;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_B3;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_B4;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_B5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_B6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_BO5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_BO6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_BQ;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_BX;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_B_CY;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_B_XOR;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_C;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_C1;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_C2;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_C3;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_C4;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_C5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_C6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_CE;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_CLK;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_CO5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_CO6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_CQ;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_CX;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_C_CY;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_C_XOR;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_D;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_D1;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_D2;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_D3;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_D4;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_D5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_D6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_DO5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_DO6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_DQ;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_DX;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_D_CY;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_D_XOR;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_A;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_A1;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_A2;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_A3;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_A4;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_A5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_A6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_AO5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_AO6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_AQ;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_AX;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_A_CY;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_A_XOR;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_B;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_B1;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_B2;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_B3;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_B4;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_B5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_B6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_BO5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_BO6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_BQ;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_BX;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_B_CY;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_B_XOR;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_C;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_C1;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_C2;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_C3;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_C4;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_C5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_C6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_CE;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_CLK;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_CO5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_CO6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_CQ;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_CX;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_C_CY;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_C_XOR;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_D;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_D1;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_D2;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_D3;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_D4;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_D5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_D6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_DO5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_DO6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_DQ;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_DX;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_D_CY;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_D_XOR;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_A;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_A1;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_A2;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_A3;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_A4;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_A5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_A6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_AO5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_AO6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_AQ;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_AX;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_A_CY;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_A_XOR;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_B;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_B1;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_B2;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_B3;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_B4;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_B5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_B6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_BO5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_BO6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_BQ;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_BX;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_B_CY;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_B_XOR;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_C;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_C1;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_C2;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_C3;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_C4;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_C5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_C6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_CE;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_CLK;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_CO5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_CO6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_CQ;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_CX;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_C_CY;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_C_XOR;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_D;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_D1;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_D2;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_D3;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_D4;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_D5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_D6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_DO5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_DO6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_DQ;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_DX;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_D_CY;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_D_XOR;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_A;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_A1;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_A2;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_A3;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_A4;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_A5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_A6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_AO5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_AO6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_AQ;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_AX;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_A_CY;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_A_XOR;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_B;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_B1;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_B2;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_B3;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_B4;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_B5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_B6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_BO5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_BO6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_BQ;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_BX;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_B_CY;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_B_XOR;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_C;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_C1;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_C2;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_C3;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_C4;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_C5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_C6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_CE;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_CLK;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_CO5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_CO6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_CQ;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_CX;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_C_CY;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_C_XOR;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_D;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_D1;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_D2;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_D3;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_D4;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_D5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_D6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_DO5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_DO6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_DQ;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_DX;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_D_CY;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_D_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_AO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_AO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_BO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_BO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_CLK;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_CO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_CO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_DO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_DO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_AMUX;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_AO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_AO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_AQ;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_BMUX;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_BO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_BO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_BQ;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_CLK;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_CO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_CO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_CQ;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_DO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_DO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_AMUX;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_AO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_AO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_AQ;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_BO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_BO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_BQ;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_CLK;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_CMUX;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_CO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_CO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_DO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_DO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_AMUX;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_AO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_AO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_AQ;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B5Q;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_BMUX;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_BO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_BO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_BQ;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_BX;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_CLK;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_CO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_DO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_DO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_AMUX;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_AO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_AO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_AX;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B5Q;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_BMUX;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_BO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_BO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_BX;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_CLK;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_CMUX;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_CO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_CO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_CQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_CX;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_DO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_DO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_AMUX;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_AO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_AO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B5Q;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_BMUX;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_BO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_BO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_BQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_BX;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_CLK;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_CO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_CO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_CQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_DO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_DO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_DQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_DX;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_AMUX;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_AO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_AO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_AQ;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_BO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_BO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_CLK;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_CO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_CO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_DO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_DO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_AO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_AO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_AQ;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_AX;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_BO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_BO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_CLK;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_CO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_CO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_DO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_DO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A5Q;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_AMUX;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_AO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_AO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_AQ;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_AX;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_BO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_BO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_BQ;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_CLK;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_CO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_CO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_DO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_DO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_AMUX;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_AO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_AO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_AQ;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_AX;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B5Q;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_BMUX;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_BO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_BO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_BQ;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_BX;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_CLK;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_CO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_CO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_DO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_DO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_AMUX;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_AO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_AO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_AQ;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B5Q;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_BMUX;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_BO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_BO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_BX;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_CLK;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_CO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_CO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_CQ;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_DMUX;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_DO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_DO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_DQ;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_DX;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A5Q;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_AMUX;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_AO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_AO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_AQ;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_AX;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_BO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_BO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_BQ;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_BX;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_CLK;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_CO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_CO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_CQ;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_CX;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_DO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_DO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A5Q;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_AMUX;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_AO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_AO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_AQ;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_AX;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_BMUX;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_BO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_BO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_CLK;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_CO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_CO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_CQ;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_DO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_DO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A5Q;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_AMUX;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_AO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_AO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_AQ;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_AX;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_BMUX;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_BO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_BO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_CLK;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_CO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_CO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_CQ;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_DO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_DO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_AMUX;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_AO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_AO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_AQ;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B5Q;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_BMUX;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_BO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_BO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_BQ;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_BX;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_CLK;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_CO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_CO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_DO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_DO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A5Q;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_AMUX;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_AO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_AO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_AQ;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_AX;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B5Q;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_BMUX;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_BO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_BO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_BQ;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_BX;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_CLK;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_CO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_CO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_DO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_AMUX;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_AO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_AO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_AQ;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_BO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_BO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_BQ;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_BX;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_CLK;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_CO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_CO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_DO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_DO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_AO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_AO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_AQ;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_BO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_BO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_BQ;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_CLK;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_CO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_CO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_CQ;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_DO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_DO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_AMUX;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_AO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_AO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_BMUX;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_BO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_BO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_CO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_CO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_DMUX;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_DO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_DO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A5Q;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_AMUX;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_AO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_AO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_AQ;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_BO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_BO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_BQ;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_CLK;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_CO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_CO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_CQ;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_DO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_DO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_AO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_AO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_BO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_BO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_CO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_CO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_DO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_DO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_AO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_AO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_AQ;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_BO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_BO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_CLK;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_CO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_CO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_DO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_DO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_AO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_AO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_BO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_BO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_CMUX;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_CO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_CO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_DO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_DO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_AO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_AO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_BO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_BO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_CO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_CO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_DO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_DO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_AMUX;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_AO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_AO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_BO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_BO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_CO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_CO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_DO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_DO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_AO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_AO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_AQ;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_BO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_BO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_CLK;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_CO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_CO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_DO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_AO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_AO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_BO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_BQ;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_CLK;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_CO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_CO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_DO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_DO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_AO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_AO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_AQ;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_BO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_BO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_CLK;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_CO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_CO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_DO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_DO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_AO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_AO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_BMUX;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_BO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_BO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_CO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_CO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_DO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_DO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_AO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_AO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_BO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_BO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_CO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_CO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_DO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_DO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_AO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_AO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_BO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_BO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_CO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_CO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_DO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_DO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_AO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_AO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_BO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_BO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_CO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_CO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_DO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_DO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D_XOR;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_A;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_A1;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_A2;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_A3;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_A4;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_A5;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_A6;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_AO5;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_AO6;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_AQ;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_AX;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_A_CY;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_A_XOR;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_B;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_B1;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_B2;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_B3;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_B4;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_B5;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_B6;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_BO5;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_BO6;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_BQ;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_BX;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_B_CY;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_B_XOR;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_C;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_C1;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_C2;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_C3;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_C4;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_C5;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_C6;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_CE;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_CLK;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_CO5;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_CO6;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_CQ;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_CX;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_C_CY;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_C_XOR;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_D;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_D1;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_D2;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_D3;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_D4;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_D5;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_D6;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_DO5;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_DO6;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_DQ;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_DX;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_D_CY;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_D_XOR;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_A;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_A1;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_A2;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_A3;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_A4;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_A5;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_A6;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_AO5;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_AO6;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_A_CY;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_A_XOR;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_B;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_B1;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_B2;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_B3;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_B4;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_B5;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_B6;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_BO5;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_BO6;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_B_CY;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_B_XOR;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_C;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_C1;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_C2;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_C3;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_C4;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_C5;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_C6;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_CO5;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_CO6;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_C_CY;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_C_XOR;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_D;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_D1;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_D2;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_D3;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_D4;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_D5;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_D6;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_DO5;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_DO6;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_D_CY;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_D_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_AO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_AO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_AQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B5Q;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_BMUX;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_BO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_BO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_BQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C5Q;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_CLK;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_CMUX;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_CO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_CO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_CQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_DO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_DO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_AO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_AO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_AQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_AX;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_BO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_BO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_BX;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_CLK;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_CO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_CO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_DO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_DO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_AO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_AO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_AQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_BO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_BO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_CLK;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_CO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_CO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_CQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D5Q;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_DMUX;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_DO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_DO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_DQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_AO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_AO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_AX;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_BO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_BO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_CLK;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_CO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_CO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_DO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_DO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A5Q;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_AMUX;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_AO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_AO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_BO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_BO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_CLK;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_CO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_CO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_DO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_DO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_AO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_AO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_BO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_BO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_CO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_CO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_DO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_DO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A5Q;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_AMUX;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_AO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_AO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_BO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_BO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_BQ;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_CLK;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_CO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_CO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_DO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_DO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_AO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_AO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_AQ;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_BO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_BO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_CLK;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_CO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_CO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_DO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_DO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A5Q;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_AMUX;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_AO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_AO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B5Q;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_BMUX;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_BO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_BO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_BQ;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_CLK;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_CO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_CO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_CQ;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_DO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_DO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_DQ;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A5Q;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_AMUX;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_AO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_AO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_AQ;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B5Q;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_BMUX;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_BO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_BO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_BQ;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_CLK;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_CO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_CO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_CQ;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_DO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_DO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_AMUX;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_AO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_AO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_AX;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B5Q;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_BMUX;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_BO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_BO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_BQ;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_BX;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_CLK;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_CO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_DO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_DO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_AO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_AO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_AQ;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_BO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_BO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_BQ;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_CLK;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_CO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_CO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_CQ;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_DO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_DO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_DQ;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_AMUX;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_AO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_AO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_BO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_BO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_CO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_CO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_DO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_DO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A5Q;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_AMUX;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_AO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_AO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_BO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_BO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_BQ;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_CLK;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_CO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_CO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_CQ;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_DO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_DO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_DQ;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A5Q;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_AMUX;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_AO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_AO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_BO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_BO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_BQ;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_BX;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_CLK;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_CO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_CO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_CQ;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_CX;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_DO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_DO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_AO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_AO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_AQ;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_BMUX;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_BO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_BO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_CLK;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_CO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_CO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_DO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_DO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_AO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_AO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_BO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_BO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_CO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_CO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_DO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_DO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_AO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_AO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_AQ;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_BO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_BQ;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_CLK;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_CO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_CO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_DO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_DO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_AMUX;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_AO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_AO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_BO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_BO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_CO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_CO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_DMUX;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_DO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_DO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A5Q;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_AMUX;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_AO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_AO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_AQ;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B5Q;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_BMUX;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_BO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_BO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_BQ;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_CLK;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_CO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_CO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_DO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_DO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_AO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_AO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_BO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_BO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_CO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_CO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_DO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_DO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_AO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_AO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_BO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_BO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_CMUX;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_CO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_DO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_DO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A5Q;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_AMUX;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_AO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_AO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_AQ;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_BO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_BO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_BQ;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_CLK;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_CO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_CO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_DO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_DO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_AMUX;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_AO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_AO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_BMUX;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_BO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_BO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_CO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_CO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_DO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_DO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A5Q;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_AMUX;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_AO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_AO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_AQ;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_BO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_BO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_BQ;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_CLK;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_CO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_CO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_DO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_DO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_AO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_AO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_AQ;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_BO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_BO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_BQ;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_CLK;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_CO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_CO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_CQ;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_DO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_DO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_DQ;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_AMUX;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_AO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_AO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_BO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_BO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_CO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_CO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_DO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_DO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_AO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_AO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_AQ;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_BO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_BQ;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_CLK;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_CO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_CO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_CQ;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_DO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_DO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_DQ;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_AO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_AO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_BO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_BO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_CO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_CO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_DMUX;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_DO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_DO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_AO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_AO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_BO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_BO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_CO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_CO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_DO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_AO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_AO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_BO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_BO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_CO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_CO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_DO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_DO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_AO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_AO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_BO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_BO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_CO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_CO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_DO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_DO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D_XOR;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  wire [0:0] CLK_HROW_BOT_R_X139Y78_BUFHCE_X0Y20_CE;
  wire [0:0] CLK_HROW_BOT_R_X139Y78_BUFHCE_X0Y20_I;
  wire [0:0] CLK_HROW_BOT_R_X139Y78_BUFHCE_X0Y20_O;
  wire [0:0] CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_CE;
  wire [0:0] CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_I;
  wire [0:0] CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  wire [0:0] CLK_HROW_TOP_R_X139Y182_BUFHCE_X1Y44_CE;
  wire [0:0] CLK_HROW_TOP_R_X139Y182_BUFHCE_X1Y44_I;
  wire [0:0] CLK_HROW_TOP_R_X139Y182_BUFHCE_X1Y44_O;
  wire [0:0] LIOB33_SING_X0Y0_IOB_X0Y0_I;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_O;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_I;
  wire [0:0] LIOB33_SING_X0Y150_IOB_X0Y150_I;
  wire [0:0] LIOB33_SING_X0Y199_IOB_X0Y199_I;
  wire [0:0] LIOB33_SING_X0Y200_IOB_X0Y200_I;
  wire [0:0] LIOB33_SING_X0Y249_IOB_X0Y249_I;
  wire [0:0] LIOB33_SING_X0Y50_IOB_X0Y50_I;
  wire [0:0] LIOB33_SING_X0Y99_IOB_X0Y99_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_I;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_I;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_I;
  wire [0:0] LIOB33_X0Y11_IOB_X0Y11_I;
  wire [0:0] LIOB33_X0Y11_IOB_X0Y12_I;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_I;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_I;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_I;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_I;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_I;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_I;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_I;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_I;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_I;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_I;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_I;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_I;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_I;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_I;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_I;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_I;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_I;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_I;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_I;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_I;
  wire [0:0] LIOB33_X0Y13_IOB_X0Y13_I;
  wire [0:0] LIOB33_X0Y13_IOB_X0Y14_I;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_I;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_I;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_I;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_I;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_I;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_I;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_I;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y151_I;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y152_I;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y153_I;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y154_I;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y155_I;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y156_I;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y157_I;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y158_I;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y159_I;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y160_I;
  wire [0:0] LIOB33_X0Y15_IOB_X0Y15_I;
  wire [0:0] LIOB33_X0Y15_IOB_X0Y16_I;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y161_I;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y162_I;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y163_I;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y164_I;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y165_I;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y166_I;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y167_I;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y168_I;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y169_I;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y170_I;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y171_I;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y172_I;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y173_I;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y174_I;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y175_I;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y176_I;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y177_I;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y178_I;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y179_I;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y180_I;
  wire [0:0] LIOB33_X0Y17_IOB_X0Y17_I;
  wire [0:0] LIOB33_X0Y17_IOB_X0Y18_I;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y181_I;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y182_I;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y183_I;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y184_I;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y185_I;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y186_I;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y187_I;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y188_I;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y189_I;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y190_I;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y191_I;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y192_I;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y193_I;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y194_I;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y195_I;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y196_I;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y197_I;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y198_I;
  wire [0:0] LIOB33_X0Y19_IOB_X0Y19_I;
  wire [0:0] LIOB33_X0Y19_IOB_X0Y20_I;
  wire [0:0] LIOB33_X0Y1_IOB_X0Y1_I;
  wire [0:0] LIOB33_X0Y1_IOB_X0Y2_I;
  wire [0:0] LIOB33_X0Y201_IOB_X0Y201_I;
  wire [0:0] LIOB33_X0Y201_IOB_X0Y202_I;
  wire [0:0] LIOB33_X0Y203_IOB_X0Y203_I;
  wire [0:0] LIOB33_X0Y203_IOB_X0Y204_I;
  wire [0:0] LIOB33_X0Y205_IOB_X0Y205_I;
  wire [0:0] LIOB33_X0Y205_IOB_X0Y206_I;
  wire [0:0] LIOB33_X0Y207_IOB_X0Y207_I;
  wire [0:0] LIOB33_X0Y207_IOB_X0Y208_I;
  wire [0:0] LIOB33_X0Y209_IOB_X0Y209_I;
  wire [0:0] LIOB33_X0Y209_IOB_X0Y210_I;
  wire [0:0] LIOB33_X0Y211_IOB_X0Y211_I;
  wire [0:0] LIOB33_X0Y211_IOB_X0Y212_I;
  wire [0:0] LIOB33_X0Y213_IOB_X0Y213_I;
  wire [0:0] LIOB33_X0Y213_IOB_X0Y214_I;
  wire [0:0] LIOB33_X0Y215_IOB_X0Y215_I;
  wire [0:0] LIOB33_X0Y215_IOB_X0Y216_I;
  wire [0:0] LIOB33_X0Y217_IOB_X0Y217_I;
  wire [0:0] LIOB33_X0Y217_IOB_X0Y218_I;
  wire [0:0] LIOB33_X0Y219_IOB_X0Y219_I;
  wire [0:0] LIOB33_X0Y219_IOB_X0Y220_I;
  wire [0:0] LIOB33_X0Y21_IOB_X0Y21_I;
  wire [0:0] LIOB33_X0Y21_IOB_X0Y22_I;
  wire [0:0] LIOB33_X0Y221_IOB_X0Y221_I;
  wire [0:0] LIOB33_X0Y221_IOB_X0Y222_I;
  wire [0:0] LIOB33_X0Y223_IOB_X0Y223_I;
  wire [0:0] LIOB33_X0Y223_IOB_X0Y224_I;
  wire [0:0] LIOB33_X0Y225_IOB_X0Y225_I;
  wire [0:0] LIOB33_X0Y225_IOB_X0Y226_I;
  wire [0:0] LIOB33_X0Y227_IOB_X0Y227_I;
  wire [0:0] LIOB33_X0Y227_IOB_X0Y228_I;
  wire [0:0] LIOB33_X0Y229_IOB_X0Y229_I;
  wire [0:0] LIOB33_X0Y229_IOB_X0Y230_I;
  wire [0:0] LIOB33_X0Y231_IOB_X0Y231_I;
  wire [0:0] LIOB33_X0Y231_IOB_X0Y232_I;
  wire [0:0] LIOB33_X0Y233_IOB_X0Y233_I;
  wire [0:0] LIOB33_X0Y233_IOB_X0Y234_I;
  wire [0:0] LIOB33_X0Y235_IOB_X0Y235_I;
  wire [0:0] LIOB33_X0Y235_IOB_X0Y236_I;
  wire [0:0] LIOB33_X0Y237_IOB_X0Y237_I;
  wire [0:0] LIOB33_X0Y237_IOB_X0Y238_I;
  wire [0:0] LIOB33_X0Y239_IOB_X0Y239_I;
  wire [0:0] LIOB33_X0Y239_IOB_X0Y240_I;
  wire [0:0] LIOB33_X0Y23_IOB_X0Y23_I;
  wire [0:0] LIOB33_X0Y23_IOB_X0Y24_I;
  wire [0:0] LIOB33_X0Y241_IOB_X0Y241_I;
  wire [0:0] LIOB33_X0Y241_IOB_X0Y242_I;
  wire [0:0] LIOB33_X0Y243_IOB_X0Y243_I;
  wire [0:0] LIOB33_X0Y243_IOB_X0Y244_I;
  wire [0:0] LIOB33_X0Y245_IOB_X0Y245_I;
  wire [0:0] LIOB33_X0Y245_IOB_X0Y246_I;
  wire [0:0] LIOB33_X0Y247_IOB_X0Y247_I;
  wire [0:0] LIOB33_X0Y247_IOB_X0Y248_I;
  wire [0:0] LIOB33_X0Y25_IOB_X0Y25_I;
  wire [0:0] LIOB33_X0Y25_IOB_X0Y26_I;
  wire [0:0] LIOB33_X0Y27_IOB_X0Y27_I;
  wire [0:0] LIOB33_X0Y27_IOB_X0Y28_I;
  wire [0:0] LIOB33_X0Y29_IOB_X0Y29_I;
  wire [0:0] LIOB33_X0Y29_IOB_X0Y30_I;
  wire [0:0] LIOB33_X0Y31_IOB_X0Y31_I;
  wire [0:0] LIOB33_X0Y3_IOB_X0Y3_I;
  wire [0:0] LIOB33_X0Y3_IOB_X0Y4_I;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y51_I;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y52_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y53_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y54_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y55_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y56_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y57_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y58_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y59_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y60_I;
  wire [0:0] LIOB33_X0Y5_IOB_X0Y5_I;
  wire [0:0] LIOB33_X0Y5_IOB_X0Y6_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y61_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y62_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y63_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y64_I;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y65_I;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y66_I;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y67_I;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y68_I;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y69_I;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y70_I;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y71_I;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y72_I;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y73_I;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y74_I;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y75_I;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y76_I;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y77_I;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y78_I;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y79_I;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y80_I;
  wire [0:0] LIOB33_X0Y7_IOB_X0Y7_I;
  wire [0:0] LIOB33_X0Y7_IOB_X0Y8_I;
  wire [0:0] LIOB33_X0Y81_IOB_X0Y81_I;
  wire [0:0] LIOB33_X0Y81_IOB_X0Y82_I;
  wire [0:0] LIOB33_X0Y83_IOB_X0Y83_I;
  wire [0:0] LIOB33_X0Y83_IOB_X0Y84_I;
  wire [0:0] LIOB33_X0Y85_IOB_X0Y85_I;
  wire [0:0] LIOB33_X0Y85_IOB_X0Y86_I;
  wire [0:0] LIOB33_X0Y87_IOB_X0Y87_I;
  wire [0:0] LIOB33_X0Y87_IOB_X0Y88_I;
  wire [0:0] LIOB33_X0Y89_IOB_X0Y89_I;
  wire [0:0] LIOB33_X0Y89_IOB_X0Y90_I;
  wire [0:0] LIOB33_X0Y91_IOB_X0Y91_I;
  wire [0:0] LIOB33_X0Y91_IOB_X0Y92_I;
  wire [0:0] LIOB33_X0Y93_IOB_X0Y93_I;
  wire [0:0] LIOB33_X0Y93_IOB_X0Y94_I;
  wire [0:0] LIOB33_X0Y95_IOB_X0Y95_I;
  wire [0:0] LIOB33_X0Y95_IOB_X0Y96_I;
  wire [0:0] LIOB33_X0Y97_IOB_X0Y97_I;
  wire [0:0] LIOB33_X0Y97_IOB_X0Y98_I;
  wire [0:0] LIOB33_X0Y9_IOB_X0Y10_I;
  wire [0:0] LIOB33_X0Y9_IOB_X0Y9_I;
  wire [0:0] LIOI3_SING_X0Y0_ILOGIC_X0Y0_D;
  wire [0:0] LIOI3_SING_X0Y0_ILOGIC_X0Y0_O;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ;
  wire [0:0] LIOI3_SING_X0Y149_ILOGIC_X0Y149_D;
  wire [0:0] LIOI3_SING_X0Y149_ILOGIC_X0Y149_O;
  wire [0:0] LIOI3_SING_X0Y150_ILOGIC_X0Y150_D;
  wire [0:0] LIOI3_SING_X0Y150_ILOGIC_X0Y150_O;
  wire [0:0] LIOI3_SING_X0Y199_ILOGIC_X0Y199_D;
  wire [0:0] LIOI3_SING_X0Y199_ILOGIC_X0Y199_O;
  wire [0:0] LIOI3_SING_X0Y200_ILOGIC_X0Y200_D;
  wire [0:0] LIOI3_SING_X0Y200_ILOGIC_X0Y200_O;
  wire [0:0] LIOI3_SING_X0Y249_ILOGIC_X0Y249_D;
  wire [0:0] LIOI3_SING_X0Y249_ILOGIC_X0Y249_O;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_D;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_O;
  wire [0:0] LIOI3_SING_X0Y99_ILOGIC_X0Y99_D;
  wire [0:0] LIOI3_SING_X0Y99_ILOGIC_X0Y99_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y119_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y119_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y131_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y131_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y132_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y132_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_ILOGIC_X0Y143_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_ILOGIC_X0Y143_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_ILOGIC_X0Y144_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_ILOGIC_X0Y144_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y157_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y157_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y158_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y158_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y169_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y169_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y170_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y170_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y181_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y181_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y182_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y182_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y193_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y193_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y194_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y194_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y19_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y19_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y20_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y20_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y207_ILOGIC_X0Y207_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y207_ILOGIC_X0Y207_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y207_ILOGIC_X0Y208_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y207_ILOGIC_X0Y208_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y219_ILOGIC_X0Y219_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y219_ILOGIC_X0Y219_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y219_ILOGIC_X0Y220_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y219_ILOGIC_X0Y220_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y231_ILOGIC_X0Y231_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y231_ILOGIC_X0Y231_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y231_ILOGIC_X0Y232_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y231_ILOGIC_X0Y232_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y243_ILOGIC_X0Y243_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y243_ILOGIC_X0Y243_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y243_ILOGIC_X0Y244_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y243_ILOGIC_X0Y244_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y31_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y31_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y7_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y7_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y8_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y8_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y81_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y81_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y82_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y82_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_ILOGIC_X0Y93_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_ILOGIC_X0Y93_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_ILOGIC_X0Y94_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_ILOGIC_X0Y94_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y138_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y138_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y13_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y13_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y14_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y14_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y163_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y163_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y164_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y164_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y187_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y187_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y188_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y188_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y213_ILOGIC_X0Y213_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y213_ILOGIC_X0Y213_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y213_ILOGIC_X0Y214_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y213_ILOGIC_X0Y214_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y237_ILOGIC_X0Y237_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y237_ILOGIC_X0Y237_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y237_ILOGIC_X0Y238_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y237_ILOGIC_X0Y238_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_ILOGIC_X0Y87_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_ILOGIC_X0Y87_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_ILOGIC_X0Y88_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_ILOGIC_X0Y88_O;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_O;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_O;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_D;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_O;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y118_D;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y118_O;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y11_D;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y11_O;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y12_D;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y12_O;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y121_D;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y121_O;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y122_D;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y122_O;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y123_D;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y123_O;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y124_D;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y124_O;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y125_D;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y125_O;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y126_D;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y126_O;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y127_D;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y127_O;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y128_D;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y128_O;
  wire [0:0] LIOI3_X0Y129_ILOGIC_X0Y129_D;
  wire [0:0] LIOI3_X0Y129_ILOGIC_X0Y129_O;
  wire [0:0] LIOI3_X0Y129_ILOGIC_X0Y130_D;
  wire [0:0] LIOI3_X0Y129_ILOGIC_X0Y130_O;
  wire [0:0] LIOI3_X0Y133_ILOGIC_X0Y133_D;
  wire [0:0] LIOI3_X0Y133_ILOGIC_X0Y133_O;
  wire [0:0] LIOI3_X0Y133_ILOGIC_X0Y134_D;
  wire [0:0] LIOI3_X0Y133_ILOGIC_X0Y134_O;
  wire [0:0] LIOI3_X0Y135_ILOGIC_X0Y135_D;
  wire [0:0] LIOI3_X0Y135_ILOGIC_X0Y135_O;
  wire [0:0] LIOI3_X0Y135_ILOGIC_X0Y136_D;
  wire [0:0] LIOI3_X0Y135_ILOGIC_X0Y136_O;
  wire [0:0] LIOI3_X0Y139_ILOGIC_X0Y139_D;
  wire [0:0] LIOI3_X0Y139_ILOGIC_X0Y139_O;
  wire [0:0] LIOI3_X0Y139_ILOGIC_X0Y140_D;
  wire [0:0] LIOI3_X0Y139_ILOGIC_X0Y140_O;
  wire [0:0] LIOI3_X0Y141_ILOGIC_X0Y141_D;
  wire [0:0] LIOI3_X0Y141_ILOGIC_X0Y141_O;
  wire [0:0] LIOI3_X0Y141_ILOGIC_X0Y142_D;
  wire [0:0] LIOI3_X0Y141_ILOGIC_X0Y142_O;
  wire [0:0] LIOI3_X0Y145_ILOGIC_X0Y145_D;
  wire [0:0] LIOI3_X0Y145_ILOGIC_X0Y145_O;
  wire [0:0] LIOI3_X0Y145_ILOGIC_X0Y146_D;
  wire [0:0] LIOI3_X0Y145_ILOGIC_X0Y146_O;
  wire [0:0] LIOI3_X0Y147_ILOGIC_X0Y147_D;
  wire [0:0] LIOI3_X0Y147_ILOGIC_X0Y147_O;
  wire [0:0] LIOI3_X0Y147_ILOGIC_X0Y148_D;
  wire [0:0] LIOI3_X0Y147_ILOGIC_X0Y148_O;
  wire [0:0] LIOI3_X0Y151_ILOGIC_X0Y151_D;
  wire [0:0] LIOI3_X0Y151_ILOGIC_X0Y151_O;
  wire [0:0] LIOI3_X0Y151_ILOGIC_X0Y152_D;
  wire [0:0] LIOI3_X0Y151_ILOGIC_X0Y152_O;
  wire [0:0] LIOI3_X0Y153_ILOGIC_X0Y153_D;
  wire [0:0] LIOI3_X0Y153_ILOGIC_X0Y153_O;
  wire [0:0] LIOI3_X0Y153_ILOGIC_X0Y154_D;
  wire [0:0] LIOI3_X0Y153_ILOGIC_X0Y154_O;
  wire [0:0] LIOI3_X0Y155_ILOGIC_X0Y155_D;
  wire [0:0] LIOI3_X0Y155_ILOGIC_X0Y155_O;
  wire [0:0] LIOI3_X0Y155_ILOGIC_X0Y156_D;
  wire [0:0] LIOI3_X0Y155_ILOGIC_X0Y156_O;
  wire [0:0] LIOI3_X0Y159_ILOGIC_X0Y159_D;
  wire [0:0] LIOI3_X0Y159_ILOGIC_X0Y159_O;
  wire [0:0] LIOI3_X0Y159_ILOGIC_X0Y160_D;
  wire [0:0] LIOI3_X0Y159_ILOGIC_X0Y160_O;
  wire [0:0] LIOI3_X0Y15_ILOGIC_X0Y15_D;
  wire [0:0] LIOI3_X0Y15_ILOGIC_X0Y15_O;
  wire [0:0] LIOI3_X0Y15_ILOGIC_X0Y16_D;
  wire [0:0] LIOI3_X0Y15_ILOGIC_X0Y16_O;
  wire [0:0] LIOI3_X0Y161_ILOGIC_X0Y161_D;
  wire [0:0] LIOI3_X0Y161_ILOGIC_X0Y161_O;
  wire [0:0] LIOI3_X0Y161_ILOGIC_X0Y162_D;
  wire [0:0] LIOI3_X0Y161_ILOGIC_X0Y162_O;
  wire [0:0] LIOI3_X0Y165_ILOGIC_X0Y165_D;
  wire [0:0] LIOI3_X0Y165_ILOGIC_X0Y165_O;
  wire [0:0] LIOI3_X0Y165_ILOGIC_X0Y166_D;
  wire [0:0] LIOI3_X0Y165_ILOGIC_X0Y166_O;
  wire [0:0] LIOI3_X0Y167_ILOGIC_X0Y167_D;
  wire [0:0] LIOI3_X0Y167_ILOGIC_X0Y167_O;
  wire [0:0] LIOI3_X0Y167_ILOGIC_X0Y168_D;
  wire [0:0] LIOI3_X0Y167_ILOGIC_X0Y168_O;
  wire [0:0] LIOI3_X0Y171_ILOGIC_X0Y171_D;
  wire [0:0] LIOI3_X0Y171_ILOGIC_X0Y171_O;
  wire [0:0] LIOI3_X0Y171_ILOGIC_X0Y172_D;
  wire [0:0] LIOI3_X0Y171_ILOGIC_X0Y172_O;
  wire [0:0] LIOI3_X0Y173_ILOGIC_X0Y173_D;
  wire [0:0] LIOI3_X0Y173_ILOGIC_X0Y173_O;
  wire [0:0] LIOI3_X0Y173_ILOGIC_X0Y174_D;
  wire [0:0] LIOI3_X0Y173_ILOGIC_X0Y174_O;
  wire [0:0] LIOI3_X0Y175_ILOGIC_X0Y175_D;
  wire [0:0] LIOI3_X0Y175_ILOGIC_X0Y175_O;
  wire [0:0] LIOI3_X0Y175_ILOGIC_X0Y176_D;
  wire [0:0] LIOI3_X0Y175_ILOGIC_X0Y176_O;
  wire [0:0] LIOI3_X0Y177_ILOGIC_X0Y177_D;
  wire [0:0] LIOI3_X0Y177_ILOGIC_X0Y177_O;
  wire [0:0] LIOI3_X0Y177_ILOGIC_X0Y178_D;
  wire [0:0] LIOI3_X0Y177_ILOGIC_X0Y178_O;
  wire [0:0] LIOI3_X0Y179_ILOGIC_X0Y179_D;
  wire [0:0] LIOI3_X0Y179_ILOGIC_X0Y179_O;
  wire [0:0] LIOI3_X0Y179_ILOGIC_X0Y180_D;
  wire [0:0] LIOI3_X0Y179_ILOGIC_X0Y180_O;
  wire [0:0] LIOI3_X0Y17_ILOGIC_X0Y17_D;
  wire [0:0] LIOI3_X0Y17_ILOGIC_X0Y17_O;
  wire [0:0] LIOI3_X0Y17_ILOGIC_X0Y18_D;
  wire [0:0] LIOI3_X0Y17_ILOGIC_X0Y18_O;
  wire [0:0] LIOI3_X0Y183_ILOGIC_X0Y183_D;
  wire [0:0] LIOI3_X0Y183_ILOGIC_X0Y183_O;
  wire [0:0] LIOI3_X0Y183_ILOGIC_X0Y184_D;
  wire [0:0] LIOI3_X0Y183_ILOGIC_X0Y184_O;
  wire [0:0] LIOI3_X0Y185_ILOGIC_X0Y185_D;
  wire [0:0] LIOI3_X0Y185_ILOGIC_X0Y185_O;
  wire [0:0] LIOI3_X0Y185_ILOGIC_X0Y186_D;
  wire [0:0] LIOI3_X0Y185_ILOGIC_X0Y186_O;
  wire [0:0] LIOI3_X0Y189_ILOGIC_X0Y189_D;
  wire [0:0] LIOI3_X0Y189_ILOGIC_X0Y189_O;
  wire [0:0] LIOI3_X0Y189_ILOGIC_X0Y190_D;
  wire [0:0] LIOI3_X0Y189_ILOGIC_X0Y190_O;
  wire [0:0] LIOI3_X0Y191_ILOGIC_X0Y191_D;
  wire [0:0] LIOI3_X0Y191_ILOGIC_X0Y191_O;
  wire [0:0] LIOI3_X0Y191_ILOGIC_X0Y192_D;
  wire [0:0] LIOI3_X0Y191_ILOGIC_X0Y192_O;
  wire [0:0] LIOI3_X0Y195_ILOGIC_X0Y195_D;
  wire [0:0] LIOI3_X0Y195_ILOGIC_X0Y195_O;
  wire [0:0] LIOI3_X0Y195_ILOGIC_X0Y196_D;
  wire [0:0] LIOI3_X0Y195_ILOGIC_X0Y196_O;
  wire [0:0] LIOI3_X0Y197_ILOGIC_X0Y197_D;
  wire [0:0] LIOI3_X0Y197_ILOGIC_X0Y197_O;
  wire [0:0] LIOI3_X0Y197_ILOGIC_X0Y198_D;
  wire [0:0] LIOI3_X0Y197_ILOGIC_X0Y198_O;
  wire [0:0] LIOI3_X0Y1_ILOGIC_X0Y1_D;
  wire [0:0] LIOI3_X0Y1_ILOGIC_X0Y1_O;
  wire [0:0] LIOI3_X0Y1_ILOGIC_X0Y2_D;
  wire [0:0] LIOI3_X0Y1_ILOGIC_X0Y2_O;
  wire [0:0] LIOI3_X0Y201_ILOGIC_X0Y201_D;
  wire [0:0] LIOI3_X0Y201_ILOGIC_X0Y201_O;
  wire [0:0] LIOI3_X0Y201_ILOGIC_X0Y202_D;
  wire [0:0] LIOI3_X0Y201_ILOGIC_X0Y202_O;
  wire [0:0] LIOI3_X0Y203_ILOGIC_X0Y203_D;
  wire [0:0] LIOI3_X0Y203_ILOGIC_X0Y203_O;
  wire [0:0] LIOI3_X0Y203_ILOGIC_X0Y204_D;
  wire [0:0] LIOI3_X0Y203_ILOGIC_X0Y204_O;
  wire [0:0] LIOI3_X0Y205_ILOGIC_X0Y205_D;
  wire [0:0] LIOI3_X0Y205_ILOGIC_X0Y205_O;
  wire [0:0] LIOI3_X0Y205_ILOGIC_X0Y206_D;
  wire [0:0] LIOI3_X0Y205_ILOGIC_X0Y206_O;
  wire [0:0] LIOI3_X0Y209_ILOGIC_X0Y209_D;
  wire [0:0] LIOI3_X0Y209_ILOGIC_X0Y209_O;
  wire [0:0] LIOI3_X0Y209_ILOGIC_X0Y210_D;
  wire [0:0] LIOI3_X0Y209_ILOGIC_X0Y210_O;
  wire [0:0] LIOI3_X0Y211_ILOGIC_X0Y211_D;
  wire [0:0] LIOI3_X0Y211_ILOGIC_X0Y211_O;
  wire [0:0] LIOI3_X0Y211_ILOGIC_X0Y212_D;
  wire [0:0] LIOI3_X0Y211_ILOGIC_X0Y212_O;
  wire [0:0] LIOI3_X0Y215_ILOGIC_X0Y215_D;
  wire [0:0] LIOI3_X0Y215_ILOGIC_X0Y215_O;
  wire [0:0] LIOI3_X0Y215_ILOGIC_X0Y216_D;
  wire [0:0] LIOI3_X0Y215_ILOGIC_X0Y216_O;
  wire [0:0] LIOI3_X0Y217_ILOGIC_X0Y217_D;
  wire [0:0] LIOI3_X0Y217_ILOGIC_X0Y217_O;
  wire [0:0] LIOI3_X0Y217_ILOGIC_X0Y218_D;
  wire [0:0] LIOI3_X0Y217_ILOGIC_X0Y218_O;
  wire [0:0] LIOI3_X0Y21_ILOGIC_X0Y21_D;
  wire [0:0] LIOI3_X0Y21_ILOGIC_X0Y21_O;
  wire [0:0] LIOI3_X0Y21_ILOGIC_X0Y22_D;
  wire [0:0] LIOI3_X0Y21_ILOGIC_X0Y22_O;
  wire [0:0] LIOI3_X0Y221_ILOGIC_X0Y221_D;
  wire [0:0] LIOI3_X0Y221_ILOGIC_X0Y221_O;
  wire [0:0] LIOI3_X0Y221_ILOGIC_X0Y222_D;
  wire [0:0] LIOI3_X0Y221_ILOGIC_X0Y222_O;
  wire [0:0] LIOI3_X0Y223_ILOGIC_X0Y223_D;
  wire [0:0] LIOI3_X0Y223_ILOGIC_X0Y223_O;
  wire [0:0] LIOI3_X0Y223_ILOGIC_X0Y224_D;
  wire [0:0] LIOI3_X0Y223_ILOGIC_X0Y224_O;
  wire [0:0] LIOI3_X0Y225_ILOGIC_X0Y225_D;
  wire [0:0] LIOI3_X0Y225_ILOGIC_X0Y225_O;
  wire [0:0] LIOI3_X0Y225_ILOGIC_X0Y226_D;
  wire [0:0] LIOI3_X0Y225_ILOGIC_X0Y226_O;
  wire [0:0] LIOI3_X0Y227_ILOGIC_X0Y227_D;
  wire [0:0] LIOI3_X0Y227_ILOGIC_X0Y227_O;
  wire [0:0] LIOI3_X0Y227_ILOGIC_X0Y228_D;
  wire [0:0] LIOI3_X0Y227_ILOGIC_X0Y228_O;
  wire [0:0] LIOI3_X0Y229_ILOGIC_X0Y229_D;
  wire [0:0] LIOI3_X0Y229_ILOGIC_X0Y229_O;
  wire [0:0] LIOI3_X0Y229_ILOGIC_X0Y230_D;
  wire [0:0] LIOI3_X0Y229_ILOGIC_X0Y230_O;
  wire [0:0] LIOI3_X0Y233_ILOGIC_X0Y233_D;
  wire [0:0] LIOI3_X0Y233_ILOGIC_X0Y233_O;
  wire [0:0] LIOI3_X0Y233_ILOGIC_X0Y234_D;
  wire [0:0] LIOI3_X0Y233_ILOGIC_X0Y234_O;
  wire [0:0] LIOI3_X0Y235_ILOGIC_X0Y235_D;
  wire [0:0] LIOI3_X0Y235_ILOGIC_X0Y235_O;
  wire [0:0] LIOI3_X0Y235_ILOGIC_X0Y236_D;
  wire [0:0] LIOI3_X0Y235_ILOGIC_X0Y236_O;
  wire [0:0] LIOI3_X0Y239_ILOGIC_X0Y239_D;
  wire [0:0] LIOI3_X0Y239_ILOGIC_X0Y239_O;
  wire [0:0] LIOI3_X0Y239_ILOGIC_X0Y240_D;
  wire [0:0] LIOI3_X0Y239_ILOGIC_X0Y240_O;
  wire [0:0] LIOI3_X0Y23_ILOGIC_X0Y23_D;
  wire [0:0] LIOI3_X0Y23_ILOGIC_X0Y23_O;
  wire [0:0] LIOI3_X0Y23_ILOGIC_X0Y24_D;
  wire [0:0] LIOI3_X0Y23_ILOGIC_X0Y24_O;
  wire [0:0] LIOI3_X0Y241_ILOGIC_X0Y241_D;
  wire [0:0] LIOI3_X0Y241_ILOGIC_X0Y241_O;
  wire [0:0] LIOI3_X0Y241_ILOGIC_X0Y242_D;
  wire [0:0] LIOI3_X0Y241_ILOGIC_X0Y242_O;
  wire [0:0] LIOI3_X0Y245_ILOGIC_X0Y245_D;
  wire [0:0] LIOI3_X0Y245_ILOGIC_X0Y245_O;
  wire [0:0] LIOI3_X0Y245_ILOGIC_X0Y246_D;
  wire [0:0] LIOI3_X0Y245_ILOGIC_X0Y246_O;
  wire [0:0] LIOI3_X0Y247_ILOGIC_X0Y247_D;
  wire [0:0] LIOI3_X0Y247_ILOGIC_X0Y247_O;
  wire [0:0] LIOI3_X0Y247_ILOGIC_X0Y248_D;
  wire [0:0] LIOI3_X0Y247_ILOGIC_X0Y248_O;
  wire [0:0] LIOI3_X0Y25_ILOGIC_X0Y25_D;
  wire [0:0] LIOI3_X0Y25_ILOGIC_X0Y25_O;
  wire [0:0] LIOI3_X0Y25_ILOGIC_X0Y26_D;
  wire [0:0] LIOI3_X0Y25_ILOGIC_X0Y26_O;
  wire [0:0] LIOI3_X0Y27_ILOGIC_X0Y27_D;
  wire [0:0] LIOI3_X0Y27_ILOGIC_X0Y27_O;
  wire [0:0] LIOI3_X0Y27_ILOGIC_X0Y28_D;
  wire [0:0] LIOI3_X0Y27_ILOGIC_X0Y28_O;
  wire [0:0] LIOI3_X0Y29_ILOGIC_X0Y29_D;
  wire [0:0] LIOI3_X0Y29_ILOGIC_X0Y29_O;
  wire [0:0] LIOI3_X0Y29_ILOGIC_X0Y30_D;
  wire [0:0] LIOI3_X0Y29_ILOGIC_X0Y30_O;
  wire [0:0] LIOI3_X0Y3_ILOGIC_X0Y3_D;
  wire [0:0] LIOI3_X0Y3_ILOGIC_X0Y3_O;
  wire [0:0] LIOI3_X0Y3_ILOGIC_X0Y4_D;
  wire [0:0] LIOI3_X0Y3_ILOGIC_X0Y4_O;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_O;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_O;
  wire [0:0] LIOI3_X0Y5_ILOGIC_X0Y5_D;
  wire [0:0] LIOI3_X0Y5_ILOGIC_X0Y5_O;
  wire [0:0] LIOI3_X0Y5_ILOGIC_X0Y6_D;
  wire [0:0] LIOI3_X0Y5_ILOGIC_X0Y6_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_O;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y65_D;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y65_O;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y66_D;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y66_O;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y67_D;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y67_O;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y68_D;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y68_O;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y71_D;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y71_O;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y72_D;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y72_O;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y73_D;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y73_O;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y74_D;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y74_O;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y75_D;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y75_O;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y76_D;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y76_O;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y77_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y77_O;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_O;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y79_D;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y79_O;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y80_D;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y80_O;
  wire [0:0] LIOI3_X0Y83_ILOGIC_X0Y83_D;
  wire [0:0] LIOI3_X0Y83_ILOGIC_X0Y83_O;
  wire [0:0] LIOI3_X0Y83_ILOGIC_X0Y84_D;
  wire [0:0] LIOI3_X0Y83_ILOGIC_X0Y84_O;
  wire [0:0] LIOI3_X0Y85_ILOGIC_X0Y85_D;
  wire [0:0] LIOI3_X0Y85_ILOGIC_X0Y85_O;
  wire [0:0] LIOI3_X0Y85_ILOGIC_X0Y86_D;
  wire [0:0] LIOI3_X0Y85_ILOGIC_X0Y86_O;
  wire [0:0] LIOI3_X0Y89_ILOGIC_X0Y89_D;
  wire [0:0] LIOI3_X0Y89_ILOGIC_X0Y89_O;
  wire [0:0] LIOI3_X0Y89_ILOGIC_X0Y90_D;
  wire [0:0] LIOI3_X0Y89_ILOGIC_X0Y90_O;
  wire [0:0] LIOI3_X0Y91_ILOGIC_X0Y91_D;
  wire [0:0] LIOI3_X0Y91_ILOGIC_X0Y91_O;
  wire [0:0] LIOI3_X0Y91_ILOGIC_X0Y92_D;
  wire [0:0] LIOI3_X0Y91_ILOGIC_X0Y92_O;
  wire [0:0] LIOI3_X0Y95_ILOGIC_X0Y95_D;
  wire [0:0] LIOI3_X0Y95_ILOGIC_X0Y95_O;
  wire [0:0] LIOI3_X0Y95_ILOGIC_X0Y96_D;
  wire [0:0] LIOI3_X0Y95_ILOGIC_X0Y96_O;
  wire [0:0] LIOI3_X0Y97_ILOGIC_X0Y97_D;
  wire [0:0] LIOI3_X0Y97_ILOGIC_X0Y97_O;
  wire [0:0] LIOI3_X0Y97_ILOGIC_X0Y98_D;
  wire [0:0] LIOI3_X0Y97_ILOGIC_X0Y98_O;
  wire [0:0] LIOI3_X0Y9_ILOGIC_X0Y10_D;
  wire [0:0] LIOI3_X0Y9_ILOGIC_X0Y10_O;
  wire [0:0] LIOI3_X0Y9_ILOGIC_X0Y9_D;
  wire [0:0] LIOI3_X0Y9_ILOGIC_X0Y9_O;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_O;
  wire [0:0] RIOB33_SING_X105Y149_IOB_X1Y149_O;
  wire [0:0] RIOB33_SING_X105Y150_IOB_X1Y150_O;
  wire [0:0] RIOB33_SING_X105Y199_IOB_X1Y199_I;
  wire [0:0] RIOB33_SING_X105Y200_IOB_X1Y200_I;
  wire [0:0] RIOB33_SING_X105Y50_IOB_X1Y50_O;
  wire [0:0] RIOB33_SING_X105Y99_IOB_X1Y99_O;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_O;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_O;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_O;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_O;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_O;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_O;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_O;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_O;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_O;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_O;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_O;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_O;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_O;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y114_O;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y115_O;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y116_O;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y117_O;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y118_O;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y119_O;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y120_O;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y121_O;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y122_O;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y123_O;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y124_O;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y125_O;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y126_O;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y127_O;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y128_O;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y129_O;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y130_O;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y131_O;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y132_O;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y133_O;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y134_O;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y135_O;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y136_O;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y137_O;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y138_O;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y139_O;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y140_O;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y141_O;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y142_O;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y143_O;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y144_O;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y145_O;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y146_O;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y147_O;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y148_O;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y151_O;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y152_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y153_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y154_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y155_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y156_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y157_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y158_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y159_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y160_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y161_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y162_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y163_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y164_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y165_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y166_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y167_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y168_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y169_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y170_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y171_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y172_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y173_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y174_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y175_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y176_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y177_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y178_I;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y179_I;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y180_I;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y181_I;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y182_I;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y183_I;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y184_I;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y185_I;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y186_I;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y187_I;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y188_I;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y189_I;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y190_I;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y191_I;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y192_I;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y193_I;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y194_I;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y195_I;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y196_I;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y197_I;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y198_I;
  wire [0:0] RIOB33_X105Y201_IOB_X1Y201_I;
  wire [0:0] RIOB33_X105Y201_IOB_X1Y202_I;
  wire [0:0] RIOB33_X105Y203_IOB_X1Y203_I;
  wire [0:0] RIOB33_X105Y203_IOB_X1Y204_I;
  wire [0:0] RIOB33_X105Y205_IOB_X1Y205_I;
  wire [0:0] RIOB33_X105Y51_IOB_X1Y51_O;
  wire [0:0] RIOB33_X105Y51_IOB_X1Y52_O;
  wire [0:0] RIOB33_X105Y53_IOB_X1Y53_O;
  wire [0:0] RIOB33_X105Y53_IOB_X1Y54_O;
  wire [0:0] RIOB33_X105Y55_IOB_X1Y55_O;
  wire [0:0] RIOB33_X105Y55_IOB_X1Y56_O;
  wire [0:0] RIOB33_X105Y57_IOB_X1Y57_O;
  wire [0:0] RIOB33_X105Y57_IOB_X1Y58_O;
  wire [0:0] RIOB33_X105Y59_IOB_X1Y59_O;
  wire [0:0] RIOB33_X105Y59_IOB_X1Y60_O;
  wire [0:0] RIOB33_X105Y61_IOB_X1Y61_O;
  wire [0:0] RIOB33_X105Y61_IOB_X1Y62_O;
  wire [0:0] RIOB33_X105Y63_IOB_X1Y63_O;
  wire [0:0] RIOB33_X105Y63_IOB_X1Y64_O;
  wire [0:0] RIOB33_X105Y65_IOB_X1Y65_O;
  wire [0:0] RIOB33_X105Y65_IOB_X1Y66_O;
  wire [0:0] RIOB33_X105Y67_IOB_X1Y67_O;
  wire [0:0] RIOB33_X105Y67_IOB_X1Y68_O;
  wire [0:0] RIOB33_X105Y69_IOB_X1Y69_O;
  wire [0:0] RIOB33_X105Y69_IOB_X1Y70_O;
  wire [0:0] RIOB33_X105Y71_IOB_X1Y71_O;
  wire [0:0] RIOB33_X105Y71_IOB_X1Y72_O;
  wire [0:0] RIOB33_X105Y73_IOB_X1Y73_O;
  wire [0:0] RIOB33_X105Y73_IOB_X1Y74_O;
  wire [0:0] RIOB33_X105Y75_IOB_X1Y75_O;
  wire [0:0] RIOB33_X105Y75_IOB_X1Y76_O;
  wire [0:0] RIOB33_X105Y77_IOB_X1Y77_O;
  wire [0:0] RIOB33_X105Y77_IOB_X1Y78_O;
  wire [0:0] RIOB33_X105Y79_IOB_X1Y79_O;
  wire [0:0] RIOB33_X105Y79_IOB_X1Y80_O;
  wire [0:0] RIOB33_X105Y81_IOB_X1Y81_O;
  wire [0:0] RIOB33_X105Y81_IOB_X1Y82_O;
  wire [0:0] RIOB33_X105Y83_IOB_X1Y83_O;
  wire [0:0] RIOB33_X105Y83_IOB_X1Y84_O;
  wire [0:0] RIOB33_X105Y85_IOB_X1Y85_O;
  wire [0:0] RIOB33_X105Y85_IOB_X1Y86_O;
  wire [0:0] RIOB33_X105Y87_IOB_X1Y87_O;
  wire [0:0] RIOB33_X105Y87_IOB_X1Y88_O;
  wire [0:0] RIOB33_X105Y89_IOB_X1Y89_O;
  wire [0:0] RIOB33_X105Y89_IOB_X1Y90_O;
  wire [0:0] RIOB33_X105Y91_IOB_X1Y91_O;
  wire [0:0] RIOB33_X105Y91_IOB_X1Y92_O;
  wire [0:0] RIOB33_X105Y93_IOB_X1Y93_O;
  wire [0:0] RIOB33_X105Y93_IOB_X1Y94_O;
  wire [0:0] RIOB33_X105Y95_IOB_X1Y95_O;
  wire [0:0] RIOB33_X105Y95_IOB_X1Y96_O;
  wire [0:0] RIOB33_X105Y97_IOB_X1Y97_O;
  wire [0:0] RIOB33_X105Y97_IOB_X1Y98_O;
  wire [0:0] RIOI3_SING_X105Y100_OLOGIC_X1Y100_D1;
  wire [0:0] RIOI3_SING_X105Y100_OLOGIC_X1Y100_OQ;
  wire [0:0] RIOI3_SING_X105Y100_OLOGIC_X1Y100_T1;
  wire [0:0] RIOI3_SING_X105Y100_OLOGIC_X1Y100_TQ;
  wire [0:0] RIOI3_SING_X105Y149_OLOGIC_X1Y149_D1;
  wire [0:0] RIOI3_SING_X105Y149_OLOGIC_X1Y149_OQ;
  wire [0:0] RIOI3_SING_X105Y149_OLOGIC_X1Y149_T1;
  wire [0:0] RIOI3_SING_X105Y149_OLOGIC_X1Y149_TQ;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ;
  wire [0:0] RIOI3_SING_X105Y199_ILOGIC_X1Y199_D;
  wire [0:0] RIOI3_SING_X105Y199_ILOGIC_X1Y199_O;
  wire [0:0] RIOI3_SING_X105Y200_ILOGIC_X1Y200_D;
  wire [0:0] RIOI3_SING_X105Y200_ILOGIC_X1Y200_O;
  wire [0:0] RIOI3_SING_X105Y50_OLOGIC_X1Y50_D1;
  wire [0:0] RIOI3_SING_X105Y50_OLOGIC_X1Y50_OQ;
  wire [0:0] RIOI3_SING_X105Y50_OLOGIC_X1Y50_T1;
  wire [0:0] RIOI3_SING_X105Y50_OLOGIC_X1Y50_TQ;
  wire [0:0] RIOI3_SING_X105Y99_OLOGIC_X1Y99_D1;
  wire [0:0] RIOI3_SING_X105Y99_OLOGIC_X1Y99_OQ;
  wire [0:0] RIOI3_SING_X105Y99_OLOGIC_X1Y99_T1;
  wire [0:0] RIOI3_SING_X105Y99_OLOGIC_X1Y99_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_ILOGIC_X1Y181_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_ILOGIC_X1Y181_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_ILOGIC_X1Y182_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_ILOGIC_X1Y182_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_ILOGIC_X1Y193_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_ILOGIC_X1Y193_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_ILOGIC_X1Y194_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_ILOGIC_X1Y194_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_ILOGIC_X1Y187_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_ILOGIC_X1Y187_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_ILOGIC_X1Y188_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_ILOGIC_X1Y188_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_TQ;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y101_D1;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y101_OQ;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y101_T1;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y101_TQ;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y102_D1;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y102_OQ;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y102_T1;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y102_TQ;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y103_D1;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y103_OQ;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y103_T1;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y103_TQ;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y104_D1;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y104_OQ;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y104_T1;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y104_TQ;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y105_D1;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y105_OQ;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y105_T1;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y105_TQ;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y106_D1;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y106_OQ;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y106_T1;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y106_TQ;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y109_D1;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y109_OQ;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y109_T1;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y109_TQ;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y110_D1;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y110_OQ;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y110_T1;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y110_TQ;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y111_D1;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y111_OQ;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y111_T1;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y111_TQ;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y112_D1;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y112_OQ;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y112_T1;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y112_TQ;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y115_D1;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y115_OQ;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y115_T1;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y115_TQ;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y116_D1;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y116_OQ;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y116_T1;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y116_TQ;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y117_D1;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y117_OQ;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y117_T1;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y117_TQ;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y118_D1;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y118_OQ;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y118_T1;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y118_TQ;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y121_D1;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y121_OQ;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y121_T1;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y121_TQ;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y122_D1;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y122_OQ;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y122_T1;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y122_TQ;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y123_D1;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y123_OQ;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y123_T1;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y123_TQ;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y124_D1;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y124_OQ;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y124_T1;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y124_TQ;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y125_D1;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y125_OQ;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y125_T1;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y125_TQ;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y126_D1;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y126_OQ;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y126_T1;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y126_TQ;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_D1;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_OQ;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_T1;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_TQ;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y128_D1;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y128_OQ;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y128_T1;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y128_TQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_D1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_OQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_T1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_TQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_D1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_OQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_T1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_TQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_D1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_OQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_T1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_TQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_D1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_OQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_T1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_TQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_D1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_OQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_T1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_TQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_D1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_OQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_T1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_TQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_D1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_OQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_T1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_TQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_D1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_OQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_T1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_TQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_D1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_OQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_T1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_TQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_D1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_OQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_T1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_TQ;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_D1;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_OQ;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_T1;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_TQ;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y146_D1;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y146_OQ;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y146_T1;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y146_TQ;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y147_D1;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y147_OQ;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y147_T1;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y147_TQ;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y148_D1;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y148_OQ;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y148_T1;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y148_TQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_TQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_TQ;
  wire [0:0] RIOI3_X105Y177_ILOGIC_X1Y178_D;
  wire [0:0] RIOI3_X105Y177_ILOGIC_X1Y178_O;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_TQ;
  wire [0:0] RIOI3_X105Y179_ILOGIC_X1Y179_D;
  wire [0:0] RIOI3_X105Y179_ILOGIC_X1Y179_O;
  wire [0:0] RIOI3_X105Y179_ILOGIC_X1Y180_D;
  wire [0:0] RIOI3_X105Y179_ILOGIC_X1Y180_O;
  wire [0:0] RIOI3_X105Y183_ILOGIC_X1Y183_D;
  wire [0:0] RIOI3_X105Y183_ILOGIC_X1Y183_O;
  wire [0:0] RIOI3_X105Y183_ILOGIC_X1Y184_D;
  wire [0:0] RIOI3_X105Y183_ILOGIC_X1Y184_O;
  wire [0:0] RIOI3_X105Y185_ILOGIC_X1Y185_D;
  wire [0:0] RIOI3_X105Y185_ILOGIC_X1Y185_O;
  wire [0:0] RIOI3_X105Y185_ILOGIC_X1Y186_D;
  wire [0:0] RIOI3_X105Y185_ILOGIC_X1Y186_O;
  wire [0:0] RIOI3_X105Y189_ILOGIC_X1Y189_D;
  wire [0:0] RIOI3_X105Y189_ILOGIC_X1Y189_O;
  wire [0:0] RIOI3_X105Y189_ILOGIC_X1Y190_D;
  wire [0:0] RIOI3_X105Y189_ILOGIC_X1Y190_O;
  wire [0:0] RIOI3_X105Y191_ILOGIC_X1Y191_D;
  wire [0:0] RIOI3_X105Y191_ILOGIC_X1Y191_O;
  wire [0:0] RIOI3_X105Y191_ILOGIC_X1Y192_D;
  wire [0:0] RIOI3_X105Y191_ILOGIC_X1Y192_O;
  wire [0:0] RIOI3_X105Y195_ILOGIC_X1Y195_D;
  wire [0:0] RIOI3_X105Y195_ILOGIC_X1Y195_O;
  wire [0:0] RIOI3_X105Y195_ILOGIC_X1Y196_D;
  wire [0:0] RIOI3_X105Y195_ILOGIC_X1Y196_O;
  wire [0:0] RIOI3_X105Y197_ILOGIC_X1Y197_D;
  wire [0:0] RIOI3_X105Y197_ILOGIC_X1Y197_O;
  wire [0:0] RIOI3_X105Y197_ILOGIC_X1Y198_D;
  wire [0:0] RIOI3_X105Y197_ILOGIC_X1Y198_O;
  wire [0:0] RIOI3_X105Y201_ILOGIC_X1Y201_D;
  wire [0:0] RIOI3_X105Y201_ILOGIC_X1Y201_O;
  wire [0:0] RIOI3_X105Y201_ILOGIC_X1Y202_D;
  wire [0:0] RIOI3_X105Y201_ILOGIC_X1Y202_O;
  wire [0:0] RIOI3_X105Y203_ILOGIC_X1Y203_D;
  wire [0:0] RIOI3_X105Y203_ILOGIC_X1Y203_O;
  wire [0:0] RIOI3_X105Y203_ILOGIC_X1Y204_D;
  wire [0:0] RIOI3_X105Y203_ILOGIC_X1Y204_O;
  wire [0:0] RIOI3_X105Y205_ILOGIC_X1Y205_D;
  wire [0:0] RIOI3_X105Y205_ILOGIC_X1Y205_O;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y51_D1;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y51_OQ;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y51_T1;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y51_TQ;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y52_D1;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y52_OQ;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y52_T1;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y52_TQ;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y53_D1;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y53_OQ;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y53_T1;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y53_TQ;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y54_D1;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y54_OQ;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y54_T1;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y54_TQ;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y55_D1;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y55_OQ;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y55_T1;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y55_TQ;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y56_D1;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y56_OQ;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y56_T1;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y56_TQ;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y59_D1;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y59_OQ;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y59_T1;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y59_TQ;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y60_D1;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y60_OQ;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y60_T1;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y60_TQ;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y61_D1;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y61_OQ;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y61_T1;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y61_TQ;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y62_D1;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y62_OQ;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y62_T1;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y62_TQ;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y65_D1;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y65_OQ;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y65_T1;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y65_TQ;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y66_D1;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y66_OQ;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y66_T1;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y66_TQ;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y67_D1;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y67_OQ;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y67_T1;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y67_TQ;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y68_D1;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y68_OQ;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y68_T1;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y68_TQ;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y71_D1;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y71_OQ;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y71_T1;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y71_TQ;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y72_D1;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y72_OQ;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y72_T1;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y72_TQ;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y73_D1;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y73_OQ;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y73_T1;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y73_TQ;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y74_D1;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y74_OQ;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y74_T1;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y74_TQ;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y75_D1;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y75_OQ;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y75_T1;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y75_TQ;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y76_D1;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y76_OQ;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y76_T1;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y76_TQ;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y77_D1;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y77_OQ;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y77_T1;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y77_TQ;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y78_D1;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y78_OQ;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y78_T1;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y78_TQ;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y79_D1;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y79_OQ;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y79_T1;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y79_TQ;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y80_D1;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y80_OQ;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y80_T1;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y80_TQ;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y83_D1;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y83_OQ;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y83_T1;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y83_TQ;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y84_D1;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y84_OQ;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y84_T1;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y84_TQ;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y85_D1;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y85_OQ;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y85_T1;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y85_TQ;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y86_D1;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y86_OQ;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y86_T1;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y86_TQ;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y89_D1;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y89_OQ;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y89_T1;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y89_TQ;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y90_D1;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y90_OQ;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y90_T1;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y90_TQ;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y91_D1;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y91_OQ;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y91_T1;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y91_TQ;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y92_D1;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y92_OQ;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y92_T1;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y92_TQ;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y95_D1;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y95_OQ;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y95_T1;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y95_TQ;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y96_D1;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y96_OQ;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y96_T1;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y96_TQ;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y97_D1;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y97_OQ;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y97_T1;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y97_TQ;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y98_D1;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y98_OQ;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y98_T1;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y98_TQ;


  (* KEEP, DONT_TOUCH, BEL = "RAMB18E1" *)
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .IS_CLKARDCLK_INVERTED(0),
    .IS_CLKBWRCLK_INVERTED(0),
    .IS_ENARDEN_INVERTED(0),
    .IS_ENBWREN_INVERTED(0),
    .IS_RSTRAMARSTRAM_INVERTED(1),
    .IS_RSTRAMB_INVERTED(1),
    .IS_RSTREGARSTREG_INVERTED(1),
    .IS_RSTREGB_INVERTED(1),
    .RAM_MODE("TDP"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(1)
  ) BRAM_L_X6Y125_RAMB18_X0Y50_RAMB18E1 (
.ADDRARDADDR({1'b0, 1'b0, CLBLL_L_X4Y132_SLICE_X5Y132_BO6, CLBLL_L_X4Y132_SLICE_X5Y132_CO6, CLBLL_L_X4Y133_SLICE_X4Y133_CO6, CLBLL_L_X4Y133_SLICE_X5Y133_DO6, CLBLM_R_X5Y129_SLICE_X6Y129_DO6, CLBLL_L_X4Y130_SLICE_X5Y130_DO6, CLBLL_L_X4Y132_SLICE_X5Y132_DO6, CLBLM_R_X3Y130_SLICE_X3Y130_CO6, 1'b0, 1'b0, 1'b0, 1'b0}),
.ADDRBWRADDR({1'b0, 1'b0, CLBLL_L_X4Y127_SLICE_X5Y127_BO6, CLBLM_R_X5Y127_SLICE_X7Y127_CO6, CLBLM_R_X5Y127_SLICE_X7Y127_DO6, CLBLM_R_X5Y126_SLICE_X7Y126_CO6, CLBLM_R_X5Y126_SLICE_X6Y126_CO6, CLBLM_R_X5Y125_SLICE_X7Y125_DO6, CLBLM_R_X7Y125_SLICE_X8Y125_DO6, CLBLM_R_X5Y127_SLICE_X6Y127_DO6, 1'b0, 1'b0, 1'b0, 1'b0}),
.CLKARDCLK(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CLKBWRCLK(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.DIADI({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
.DIBDI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
.DIPADIP({1'b0, 1'b0}),
.DIPBDIP({1'b1, 1'b1}),
.DOADO({BRAM_L_X6Y125_RAMB18_X0Y50_DO15, BRAM_L_X6Y125_RAMB18_X0Y50_DO14, BRAM_L_X6Y125_RAMB18_X0Y50_DO13, BRAM_L_X6Y125_RAMB18_X0Y50_DO12, BRAM_L_X6Y125_RAMB18_X0Y50_DO11, BRAM_L_X6Y125_RAMB18_X0Y50_DO10, BRAM_L_X6Y125_RAMB18_X0Y50_DO9, BRAM_L_X6Y125_RAMB18_X0Y50_DO8, BRAM_L_X6Y125_RAMB18_X0Y50_DO7, BRAM_L_X6Y125_RAMB18_X0Y50_DO6, BRAM_L_X6Y125_RAMB18_X0Y50_DO5, BRAM_L_X6Y125_RAMB18_X0Y50_DO4, BRAM_L_X6Y125_RAMB18_X0Y50_DO3, BRAM_L_X6Y125_RAMB18_X0Y50_DO2, BRAM_L_X6Y125_RAMB18_X0Y50_DO1, BRAM_L_X6Y125_RAMB18_X0Y50_DO0}),
.DOBDO({BRAM_L_X6Y125_RAMB18_X0Y50_DO31, BRAM_L_X6Y125_RAMB18_X0Y50_DO30, BRAM_L_X6Y125_RAMB18_X0Y50_DO29, BRAM_L_X6Y125_RAMB18_X0Y50_DO28, BRAM_L_X6Y125_RAMB18_X0Y50_DO27, BRAM_L_X6Y125_RAMB18_X0Y50_DO26, BRAM_L_X6Y125_RAMB18_X0Y50_DO25, BRAM_L_X6Y125_RAMB18_X0Y50_DO24, BRAM_L_X6Y125_RAMB18_X0Y50_DO23, BRAM_L_X6Y125_RAMB18_X0Y50_DO22, BRAM_L_X6Y125_RAMB18_X0Y50_DO21, BRAM_L_X6Y125_RAMB18_X0Y50_DO20, BRAM_L_X6Y125_RAMB18_X0Y50_DO19, BRAM_L_X6Y125_RAMB18_X0Y50_DO18, BRAM_L_X6Y125_RAMB18_X0Y50_DO17, BRAM_L_X6Y125_RAMB18_X0Y50_DO16}),
.DOPADOP({BRAM_L_X6Y125_RAMB18_X0Y50_DOP1, BRAM_L_X6Y125_RAMB18_X0Y50_DOP0}),
.DOPBDOP({BRAM_L_X6Y125_RAMB18_X0Y50_DOP3, BRAM_L_X6Y125_RAMB18_X0Y50_DOP2}),
.ENARDEN(1'b1),
.ENBWREN(1'b1),
.REGCEAREGCE(1'b0),
.REGCEB(1'b0),
.RSTRAMARSTRAM(1'b1),
.RSTRAMB(1'b1),
.RSTREGARSTREG(1'b1),
.RSTREGB(1'b1),
.WEA({1'b0, 1'b0}),
.WEBWE({1'b0})
  );


  (* KEEP, DONT_TOUCH, BEL = "RAMB18E1" *)
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .IS_CLKARDCLK_INVERTED(0),
    .IS_CLKBWRCLK_INVERTED(0),
    .IS_ENARDEN_INVERTED(0),
    .IS_ENBWREN_INVERTED(0),
    .IS_RSTRAMARSTRAM_INVERTED(1),
    .IS_RSTRAMB_INVERTED(1),
    .IS_RSTREGARSTREG_INVERTED(1),
    .IS_RSTREGB_INVERTED(1),
    .RAM_MODE("TDP"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(1)
  ) BRAM_L_X6Y125_RAMB18_X0Y51_RAMB18E1 (
.ADDRARDADDR({1'b0, 1'b0, CLBLM_L_X8Y137_SLICE_X11Y137_DO6, CLBLM_L_X8Y136_SLICE_X11Y136_DO6, CLBLM_L_X10Y137_SLICE_X12Y137_DO6, CLBLM_L_X10Y134_SLICE_X13Y134_BO6, CLBLM_R_X7Y134_SLICE_X8Y134_CO6, CLBLM_R_X7Y134_SLICE_X8Y134_DO6, CLBLM_R_X7Y136_SLICE_X8Y136_CO6, CLBLM_R_X7Y136_SLICE_X8Y136_DO6, 1'b0, 1'b0, 1'b0, 1'b0}),
.ADDRBWRADDR({1'b0, 1'b0, CLBLL_L_X4Y131_SLICE_X5Y131_DO6, CLBLM_R_X5Y132_SLICE_X7Y132_DO6, CLBLM_R_X7Y133_SLICE_X8Y133_DO6, CLBLM_R_X7Y132_SLICE_X8Y132_CO6, CLBLM_R_X7Y131_SLICE_X8Y131_CO6, CLBLM_R_X7Y130_SLICE_X8Y130_DO6, CLBLM_R_X7Y131_SLICE_X8Y131_DO6, CLBLM_R_X7Y132_SLICE_X8Y132_DO6, 1'b0, 1'b0, 1'b0, 1'b0}),
.CLKARDCLK(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CLKBWRCLK(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.DIADI({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
.DIBDI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
.DIPADIP({1'b0, 1'b0}),
.DIPBDIP({1'b1, 1'b1}),
.DOADO({BRAM_L_X6Y125_RAMB18_X0Y51_DOADO15, BRAM_L_X6Y125_RAMB18_X0Y51_DOADO14, BRAM_L_X6Y125_RAMB18_X0Y51_DOADO13, BRAM_L_X6Y125_RAMB18_X0Y51_DOADO12, BRAM_L_X6Y125_RAMB18_X0Y51_DOADO11, BRAM_L_X6Y125_RAMB18_X0Y51_DOADO10, BRAM_L_X6Y125_RAMB18_X0Y51_DOADO9, BRAM_L_X6Y125_RAMB18_X0Y51_DOADO8, BRAM_L_X6Y125_RAMB18_X0Y51_DOADO7, BRAM_L_X6Y125_RAMB18_X0Y51_DOADO6, BRAM_L_X6Y125_RAMB18_X0Y51_DOADO5, BRAM_L_X6Y125_RAMB18_X0Y51_DOADO4, BRAM_L_X6Y125_RAMB18_X0Y51_DOADO3, BRAM_L_X6Y125_RAMB18_X0Y51_DOADO2, BRAM_L_X6Y125_RAMB18_X0Y51_DOADO1, BRAM_L_X6Y125_RAMB18_X0Y51_DOADO0}),
.DOBDO({BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO15, BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO14, BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO13, BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO12, BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO11, BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO10, BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO9, BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO8, BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO7, BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO6, BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO5, BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO4, BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO3, BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO2, BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO1, BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO0}),
.DOPADOP({BRAM_L_X6Y125_RAMB18_X0Y51_DOPADOP1, BRAM_L_X6Y125_RAMB18_X0Y51_DOPADOP0}),
.DOPBDOP({BRAM_L_X6Y125_RAMB18_X0Y51_DOPBDOP1, BRAM_L_X6Y125_RAMB18_X0Y51_DOPBDOP0}),
.ENARDEN(1'b1),
.ENBWREN(1'b1),
.REGCEAREGCE(1'b0),
.REGCEB(1'b0),
.RSTRAMARSTRAM(1'b1),
.RSTRAMB(1'b1),
.RSTREGARSTREG(1'b1),
.RSTREGB(1'b1),
.WEA({1'b0, 1'b0}),
.WEBWE({1'b0})
  );


  (* KEEP, DONT_TOUCH, BEL = "RAMB18E1" *)
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .IS_CLKARDCLK_INVERTED(0),
    .IS_CLKBWRCLK_INVERTED(0),
    .IS_ENARDEN_INVERTED(0),
    .IS_ENBWREN_INVERTED(0),
    .IS_RSTRAMARSTRAM_INVERTED(1),
    .IS_RSTRAMB_INVERTED(1),
    .IS_RSTREGARSTREG_INVERTED(1),
    .IS_RSTREGB_INVERTED(1),
    .RAM_MODE("TDP"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(1)
  ) BRAM_L_X6Y130_RAMB18_X0Y52_RAMB18E1 (
.ADDRARDADDR({1'b0, 1'b0, CLBLM_R_X3Y134_SLICE_X3Y134_AO6, CLBLL_L_X4Y130_SLICE_X5Y130_CO6, CLBLL_L_X4Y130_SLICE_X4Y130_DO6, CLBLM_R_X5Y130_SLICE_X6Y130_DO6, CLBLM_R_X5Y129_SLICE_X6Y129_CO6, CLBLL_L_X4Y129_SLICE_X5Y129_DO6, CLBLM_R_X5Y129_SLICE_X7Y129_CO6, CLBLM_R_X5Y129_SLICE_X7Y129_DO6, 1'b0, 1'b0, 1'b0, 1'b0}),
.ADDRBWRADDR({1'b0, 1'b0, CLBLL_L_X4Y133_SLICE_X5Y133_CO6, CLBLL_L_X4Y132_SLICE_X4Y132_DO6, CLBLM_R_X5Y132_SLICE_X6Y132_CO6, CLBLM_R_X5Y131_SLICE_X6Y131_DO6, CLBLM_R_X5Y132_SLICE_X6Y132_DO6, CLBLL_L_X4Y130_SLICE_X4Y130_CO6, CLBLL_L_X4Y130_SLICE_X5Y130_BO6, CLBLM_R_X5Y130_SLICE_X6Y130_CO6, 1'b0, 1'b0, 1'b0, 1'b0}),
.CLKARDCLK(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CLKBWRCLK(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.DIADI({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
.DIBDI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
.DIPADIP({1'b0, 1'b0}),
.DIPBDIP({1'b1, 1'b1}),
.DOADO({BRAM_L_X6Y130_RAMB18_X0Y52_DO15, BRAM_L_X6Y130_RAMB18_X0Y52_DO14, BRAM_L_X6Y130_RAMB18_X0Y52_DO13, BRAM_L_X6Y130_RAMB18_X0Y52_DO12, BRAM_L_X6Y130_RAMB18_X0Y52_DO11, BRAM_L_X6Y130_RAMB18_X0Y52_DO10, BRAM_L_X6Y130_RAMB18_X0Y52_DO9, BRAM_L_X6Y130_RAMB18_X0Y52_DO8, BRAM_L_X6Y130_RAMB18_X0Y52_DO7, BRAM_L_X6Y130_RAMB18_X0Y52_DO6, BRAM_L_X6Y130_RAMB18_X0Y52_DO5, BRAM_L_X6Y130_RAMB18_X0Y52_DO4, BRAM_L_X6Y130_RAMB18_X0Y52_DO3, BRAM_L_X6Y130_RAMB18_X0Y52_DO2, BRAM_L_X6Y130_RAMB18_X0Y52_DO1, BRAM_L_X6Y130_RAMB18_X0Y52_DO0}),
.DOBDO({BRAM_L_X6Y130_RAMB18_X0Y52_DO31, BRAM_L_X6Y130_RAMB18_X0Y52_DO30, BRAM_L_X6Y130_RAMB18_X0Y52_DO29, BRAM_L_X6Y130_RAMB18_X0Y52_DO28, BRAM_L_X6Y130_RAMB18_X0Y52_DO27, BRAM_L_X6Y130_RAMB18_X0Y52_DO26, BRAM_L_X6Y130_RAMB18_X0Y52_DO25, BRAM_L_X6Y130_RAMB18_X0Y52_DO24, BRAM_L_X6Y130_RAMB18_X0Y52_DO23, BRAM_L_X6Y130_RAMB18_X0Y52_DO22, BRAM_L_X6Y130_RAMB18_X0Y52_DO21, BRAM_L_X6Y130_RAMB18_X0Y52_DO20, BRAM_L_X6Y130_RAMB18_X0Y52_DO19, BRAM_L_X6Y130_RAMB18_X0Y52_DO18, BRAM_L_X6Y130_RAMB18_X0Y52_DO17, BRAM_L_X6Y130_RAMB18_X0Y52_DO16}),
.DOPADOP({BRAM_L_X6Y130_RAMB18_X0Y52_DOP1, BRAM_L_X6Y130_RAMB18_X0Y52_DOP0}),
.DOPBDOP({BRAM_L_X6Y130_RAMB18_X0Y52_DOP3, BRAM_L_X6Y130_RAMB18_X0Y52_DOP2}),
.ENARDEN(1'b1),
.ENBWREN(1'b1),
.REGCEAREGCE(1'b0),
.REGCEB(1'b0),
.RSTRAMARSTRAM(1'b1),
.RSTRAMB(1'b1),
.RSTREGARSTREG(1'b1),
.RSTREGB(1'b1),
.WEA({1'b0, 1'b0}),
.WEBWE({1'b0})
  );


  (* KEEP, DONT_TOUCH, BEL = "RAMB18E1" *)
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .IS_CLKARDCLK_INVERTED(0),
    .IS_CLKBWRCLK_INVERTED(0),
    .IS_ENARDEN_INVERTED(0),
    .IS_ENBWREN_INVERTED(0),
    .IS_RSTRAMARSTRAM_INVERTED(1),
    .IS_RSTRAMB_INVERTED(1),
    .IS_RSTREGARSTREG_INVERTED(1),
    .IS_RSTREGB_INVERTED(1),
    .RAM_MODE("TDP"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(1)
  ) BRAM_L_X6Y130_RAMB18_X0Y53_RAMB18E1 (
.ADDRARDADDR({1'b0, 1'b0, CLBLM_R_X3Y137_SLICE_X3Y137_DO6, CLBLL_L_X4Y135_SLICE_X4Y135_DO6, CLBLM_R_X5Y134_SLICE_X6Y134_DO6, CLBLL_L_X4Y135_SLICE_X4Y135_CO6, CLBLM_R_X5Y136_SLICE_X6Y136_BO6, CLBLM_R_X3Y137_SLICE_X2Y137_CO6, CLBLL_L_X4Y138_SLICE_X4Y138_BO6, CLBLL_L_X4Y137_SLICE_X4Y137_CO6, 1'b0, 1'b0, 1'b0, 1'b0}),
.ADDRBWRADDR({1'b0, 1'b0, CLBLL_L_X4Y134_SLICE_X5Y134_DO6, CLBLM_R_X3Y135_SLICE_X3Y135_AO6, CLBLM_R_X5Y134_SLICE_X7Y134_DO6, CLBLM_R_X7Y135_SLICE_X8Y135_AO6, CLBLM_R_X7Y133_SLICE_X8Y133_AO6, CLBLM_R_X5Y133_SLICE_X6Y133_DO6, CLBLM_R_X5Y133_SLICE_X6Y133_BO6, CLBLL_L_X4Y134_SLICE_X5Y134_CO6, 1'b0, 1'b0, 1'b0, 1'b0}),
.CLKARDCLK(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CLKBWRCLK(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.DIADI({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
.DIBDI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
.DIPADIP({1'b0, 1'b0}),
.DIPBDIP({1'b1, 1'b1}),
.DOADO({BRAM_L_X6Y130_RAMB18_X0Y53_DOADO15, BRAM_L_X6Y130_RAMB18_X0Y53_DOADO14, BRAM_L_X6Y130_RAMB18_X0Y53_DOADO13, BRAM_L_X6Y130_RAMB18_X0Y53_DOADO12, BRAM_L_X6Y130_RAMB18_X0Y53_DOADO11, BRAM_L_X6Y130_RAMB18_X0Y53_DOADO10, BRAM_L_X6Y130_RAMB18_X0Y53_DOADO9, BRAM_L_X6Y130_RAMB18_X0Y53_DOADO8, BRAM_L_X6Y130_RAMB18_X0Y53_DOADO7, BRAM_L_X6Y130_RAMB18_X0Y53_DOADO6, BRAM_L_X6Y130_RAMB18_X0Y53_DOADO5, BRAM_L_X6Y130_RAMB18_X0Y53_DOADO4, BRAM_L_X6Y130_RAMB18_X0Y53_DOADO3, BRAM_L_X6Y130_RAMB18_X0Y53_DOADO2, BRAM_L_X6Y130_RAMB18_X0Y53_DOADO1, BRAM_L_X6Y130_RAMB18_X0Y53_DOADO0}),
.DOBDO({BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO15, BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO14, BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO13, BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO12, BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO11, BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO10, BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO9, BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO8, BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO7, BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO6, BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO5, BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO4, BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO3, BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO2, BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO1, BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO0}),
.DOPADOP({BRAM_L_X6Y130_RAMB18_X0Y53_DOPADOP1, BRAM_L_X6Y130_RAMB18_X0Y53_DOPADOP0}),
.DOPBDOP({BRAM_L_X6Y130_RAMB18_X0Y53_DOPBDOP1, BRAM_L_X6Y130_RAMB18_X0Y53_DOPBDOP0}),
.ENARDEN(1'b1),
.ENBWREN(1'b1),
.REGCEAREGCE(1'b0),
.REGCEB(1'b0),
.RSTRAMARSTRAM(1'b1),
.RSTRAMB(1'b1),
.RSTREGARSTREG(1'b1),
.RSTREGB(1'b1),
.WEA({1'b0, 1'b0}),
.WEBWE({1'b0})
  );


  (* KEEP, DONT_TOUCH, BEL = "RAMB18E1" *)
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .IS_CLKARDCLK_INVERTED(0),
    .IS_CLKBWRCLK_INVERTED(0),
    .IS_ENARDEN_INVERTED(0),
    .IS_ENBWREN_INVERTED(0),
    .IS_RSTRAMARSTRAM_INVERTED(1),
    .IS_RSTRAMB_INVERTED(1),
    .IS_RSTREGARSTREG_INVERTED(1),
    .IS_RSTREGB_INVERTED(1),
    .RAM_MODE("TDP"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(1)
  ) BRAM_L_X6Y135_RAMB18_X0Y54_RAMB18E1 (
.ADDRARDADDR({1'b0, 1'b0, CLBLM_R_X3Y137_SLICE_X2Y137_DO6, CLBLM_R_X5Y136_SLICE_X7Y136_DO6, CLBLM_R_X5Y137_SLICE_X6Y137_CO6, CLBLL_L_X4Y137_SLICE_X5Y137_CO6, CLBLL_L_X4Y136_SLICE_X4Y136_CO6, CLBLL_L_X4Y136_SLICE_X5Y136_DO6, CLBLM_R_X5Y136_SLICE_X6Y136_DO6, CLBLL_L_X4Y137_SLICE_X5Y137_DO6, 1'b0, 1'b0, 1'b0, 1'b0}),
.ADDRBWRADDR({1'b0, 1'b0, CLBLM_R_X5Y137_SLICE_X6Y137_DO6, CLBLM_R_X3Y135_SLICE_X3Y135_DO6, CLBLM_R_X7Y137_SLICE_X8Y137_DO6, CLBLM_R_X7Y138_SLICE_X8Y138_AO6, CLBLM_R_X5Y135_SLICE_X7Y135_CO6, CLBLL_L_X4Y136_SLICE_X5Y136_CO6, CLBLM_R_X5Y136_SLICE_X7Y136_AO6, CLBLL_L_X4Y135_SLICE_X5Y135_DO6, 1'b0, 1'b0, 1'b0, 1'b0}),
.CLKARDCLK(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CLKBWRCLK(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.DIADI({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
.DIBDI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
.DIPADIP({1'b0, 1'b0}),
.DIPBDIP({1'b1, 1'b1}),
.DOADO({BRAM_L_X6Y135_RAMB18_X0Y54_DO15, BRAM_L_X6Y135_RAMB18_X0Y54_DO14, BRAM_L_X6Y135_RAMB18_X0Y54_DO13, BRAM_L_X6Y135_RAMB18_X0Y54_DO12, BRAM_L_X6Y135_RAMB18_X0Y54_DO11, BRAM_L_X6Y135_RAMB18_X0Y54_DO10, BRAM_L_X6Y135_RAMB18_X0Y54_DO9, BRAM_L_X6Y135_RAMB18_X0Y54_DO8, BRAM_L_X6Y135_RAMB18_X0Y54_DO7, BRAM_L_X6Y135_RAMB18_X0Y54_DO6, BRAM_L_X6Y135_RAMB18_X0Y54_DO5, BRAM_L_X6Y135_RAMB18_X0Y54_DO4, BRAM_L_X6Y135_RAMB18_X0Y54_DO3, BRAM_L_X6Y135_RAMB18_X0Y54_DO2, BRAM_L_X6Y135_RAMB18_X0Y54_DO1, BRAM_L_X6Y135_RAMB18_X0Y54_DO0}),
.DOBDO({BRAM_L_X6Y135_RAMB18_X0Y54_DO31, BRAM_L_X6Y135_RAMB18_X0Y54_DO30, BRAM_L_X6Y135_RAMB18_X0Y54_DO29, BRAM_L_X6Y135_RAMB18_X0Y54_DO28, BRAM_L_X6Y135_RAMB18_X0Y54_DO27, BRAM_L_X6Y135_RAMB18_X0Y54_DO26, BRAM_L_X6Y135_RAMB18_X0Y54_DO25, BRAM_L_X6Y135_RAMB18_X0Y54_DO24, BRAM_L_X6Y135_RAMB18_X0Y54_DO23, BRAM_L_X6Y135_RAMB18_X0Y54_DO22, BRAM_L_X6Y135_RAMB18_X0Y54_DO21, BRAM_L_X6Y135_RAMB18_X0Y54_DO20, BRAM_L_X6Y135_RAMB18_X0Y54_DO19, BRAM_L_X6Y135_RAMB18_X0Y54_DO18, BRAM_L_X6Y135_RAMB18_X0Y54_DO17, BRAM_L_X6Y135_RAMB18_X0Y54_DO16}),
.DOPADOP({BRAM_L_X6Y135_RAMB18_X0Y54_DOP1, BRAM_L_X6Y135_RAMB18_X0Y54_DOP0}),
.DOPBDOP({BRAM_L_X6Y135_RAMB18_X0Y54_DOP3, BRAM_L_X6Y135_RAMB18_X0Y54_DOP2}),
.ENARDEN(1'b1),
.ENBWREN(1'b1),
.REGCEAREGCE(1'b0),
.REGCEB(1'b0),
.RSTRAMARSTRAM(1'b1),
.RSTRAMB(1'b1),
.RSTREGARSTREG(1'b1),
.RSTREGB(1'b1),
.WEA({1'b0, 1'b0}),
.WEBWE({1'b0})
  );


  (* KEEP, DONT_TOUCH, BEL = "RAMB18E1" *)
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .IS_CLKARDCLK_INVERTED(0),
    .IS_CLKBWRCLK_INVERTED(0),
    .IS_ENARDEN_INVERTED(0),
    .IS_ENBWREN_INVERTED(0),
    .IS_RSTRAMARSTRAM_INVERTED(1),
    .IS_RSTRAMB_INVERTED(1),
    .IS_RSTREGARSTREG_INVERTED(1),
    .IS_RSTREGB_INVERTED(1),
    .RAM_MODE("TDP"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(1)
  ) BRAM_L_X6Y135_RAMB18_X0Y55_RAMB18E1 (
.ADDRARDADDR({1'b0, 1'b0, CLBLM_L_X8Y137_SLICE_X11Y137_CO6, CLBLM_L_X10Y137_SLICE_X12Y137_CO6, CLBLM_L_X10Y137_SLICE_X13Y137_BO6, CLBLM_L_X8Y136_SLICE_X11Y136_BO6, CLBLM_L_X8Y136_SLICE_X10Y136_CO6, CLBLM_R_X7Y136_SLICE_X9Y136_DO6, CLBLM_L_X8Y137_SLICE_X10Y137_DO6, CLBLM_L_X10Y136_SLICE_X12Y136_DO6, 1'b0, 1'b0, 1'b0, 1'b0}),
.ADDRBWRADDR({1'b0, 1'b0, CLBLM_R_X3Y135_SLICE_X3Y135_CO6, CLBLM_R_X3Y135_SLICE_X3Y135_BO6, CLBLM_R_X7Y135_SLICE_X8Y135_CO6, CLBLM_R_X7Y135_SLICE_X8Y135_BO6, CLBLM_R_X7Y133_SLICE_X8Y133_CO6, CLBLM_R_X7Y135_SLICE_X8Y135_DO6, CLBLM_R_X7Y132_SLICE_X8Y132_BO6, CLBLM_R_X7Y131_SLICE_X8Y131_AO6, 1'b0, 1'b0, 1'b0, 1'b0}),
.CLKARDCLK(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CLKBWRCLK(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.DIADI({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
.DIBDI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
.DIPADIP({1'b0, 1'b0}),
.DIPBDIP({1'b1, 1'b1}),
.DOADO({BRAM_L_X6Y135_RAMB18_X0Y55_DOADO15, BRAM_L_X6Y135_RAMB18_X0Y55_DOADO14, BRAM_L_X6Y135_RAMB18_X0Y55_DOADO13, BRAM_L_X6Y135_RAMB18_X0Y55_DOADO12, BRAM_L_X6Y135_RAMB18_X0Y55_DOADO11, BRAM_L_X6Y135_RAMB18_X0Y55_DOADO10, BRAM_L_X6Y135_RAMB18_X0Y55_DOADO9, BRAM_L_X6Y135_RAMB18_X0Y55_DOADO8, BRAM_L_X6Y135_RAMB18_X0Y55_DOADO7, BRAM_L_X6Y135_RAMB18_X0Y55_DOADO6, BRAM_L_X6Y135_RAMB18_X0Y55_DOADO5, BRAM_L_X6Y135_RAMB18_X0Y55_DOADO4, BRAM_L_X6Y135_RAMB18_X0Y55_DOADO3, BRAM_L_X6Y135_RAMB18_X0Y55_DOADO2, BRAM_L_X6Y135_RAMB18_X0Y55_DOADO1, BRAM_L_X6Y135_RAMB18_X0Y55_DOADO0}),
.DOBDO({BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO15, BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO14, BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO13, BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO12, BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO11, BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO10, BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO9, BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO8, BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO7, BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO6, BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO5, BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO4, BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO3, BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO2, BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO1, BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO0}),
.DOPADOP({BRAM_L_X6Y135_RAMB18_X0Y55_DOPADOP1, BRAM_L_X6Y135_RAMB18_X0Y55_DOPADOP0}),
.DOPBDOP({BRAM_L_X6Y135_RAMB18_X0Y55_DOPBDOP1, BRAM_L_X6Y135_RAMB18_X0Y55_DOPBDOP0}),
.ENARDEN(1'b1),
.ENBWREN(1'b1),
.REGCEAREGCE(1'b0),
.REGCEB(1'b0),
.RSTRAMARSTRAM(1'b1),
.RSTRAMB(1'b1),
.RSTREGARSTREG(1'b1),
.RSTREGB(1'b1),
.WEA({1'b0, 1'b0}),
.WEBWE({1'b0})
  );


  (* KEEP, DONT_TOUCH, BEL = "RAMB18E1" *)
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .IS_CLKARDCLK_INVERTED(0),
    .IS_CLKBWRCLK_INVERTED(0),
    .IS_ENARDEN_INVERTED(0),
    .IS_ENBWREN_INVERTED(0),
    .IS_RSTRAMARSTRAM_INVERTED(1),
    .IS_RSTRAMB_INVERTED(1),
    .IS_RSTREGARSTREG_INVERTED(1),
    .IS_RSTREGB_INVERTED(1),
    .RAM_MODE("TDP"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(1)
  ) BRAM_L_X6Y140_RAMB18_X0Y56_RAMB18E1 (
.ADDRARDADDR({1'b0, 1'b0, CLBLM_R_X5Y140_SLICE_X7Y140_AO6, CLBLM_R_X3Y138_SLICE_X2Y138_AO6, CLBLL_L_X4Y140_SLICE_X5Y140_BO6, CLBLM_R_X3Y138_SLICE_X3Y138_AO6, CLBLL_L_X4Y139_SLICE_X4Y139_AO6, CLBLL_L_X4Y139_SLICE_X5Y139_CO6, CLBLL_L_X4Y139_SLICE_X4Y139_BO6, CLBLM_R_X3Y139_SLICE_X2Y139_AO6, 1'b0, 1'b0, 1'b0, 1'b0}),
.ADDRBWRADDR({1'b0, 1'b0, CLBLM_R_X5Y140_SLICE_X6Y140_CO6, CLBLM_R_X7Y139_SLICE_X9Y139_DO6, CLBLM_R_X7Y140_SLICE_X8Y140_CO6, CLBLM_R_X7Y140_SLICE_X8Y140_AO6, CLBLM_R_X5Y139_SLICE_X7Y139_AO6, CLBLM_R_X5Y140_SLICE_X6Y140_BO6, CLBLM_R_X5Y140_SLICE_X6Y140_AO6, CLBLL_L_X4Y140_SLICE_X5Y140_AO6, 1'b0, 1'b0, 1'b0, 1'b0}),
.CLKARDCLK(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CLKBWRCLK(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.DIADI({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
.DIBDI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
.DIPADIP({1'b0, 1'b0}),
.DIPBDIP({1'b1, 1'b1}),
.DOADO({BRAM_L_X6Y140_RAMB18_X0Y56_DO15, BRAM_L_X6Y140_RAMB18_X0Y56_DO14, BRAM_L_X6Y140_RAMB18_X0Y56_DO13, BRAM_L_X6Y140_RAMB18_X0Y56_DO12, BRAM_L_X6Y140_RAMB18_X0Y56_DO11, BRAM_L_X6Y140_RAMB18_X0Y56_DO10, BRAM_L_X6Y140_RAMB18_X0Y56_DO9, BRAM_L_X6Y140_RAMB18_X0Y56_DO8, BRAM_L_X6Y140_RAMB18_X0Y56_DO7, BRAM_L_X6Y140_RAMB18_X0Y56_DO6, BRAM_L_X6Y140_RAMB18_X0Y56_DO5, BRAM_L_X6Y140_RAMB18_X0Y56_DO4, BRAM_L_X6Y140_RAMB18_X0Y56_DO3, BRAM_L_X6Y140_RAMB18_X0Y56_DO2, BRAM_L_X6Y140_RAMB18_X0Y56_DO1, BRAM_L_X6Y140_RAMB18_X0Y56_DO0}),
.DOBDO({BRAM_L_X6Y140_RAMB18_X0Y56_DO31, BRAM_L_X6Y140_RAMB18_X0Y56_DO30, BRAM_L_X6Y140_RAMB18_X0Y56_DO29, BRAM_L_X6Y140_RAMB18_X0Y56_DO28, BRAM_L_X6Y140_RAMB18_X0Y56_DO27, BRAM_L_X6Y140_RAMB18_X0Y56_DO26, BRAM_L_X6Y140_RAMB18_X0Y56_DO25, BRAM_L_X6Y140_RAMB18_X0Y56_DO24, BRAM_L_X6Y140_RAMB18_X0Y56_DO23, BRAM_L_X6Y140_RAMB18_X0Y56_DO22, BRAM_L_X6Y140_RAMB18_X0Y56_DO21, BRAM_L_X6Y140_RAMB18_X0Y56_DO20, BRAM_L_X6Y140_RAMB18_X0Y56_DO19, BRAM_L_X6Y140_RAMB18_X0Y56_DO18, BRAM_L_X6Y140_RAMB18_X0Y56_DO17, BRAM_L_X6Y140_RAMB18_X0Y56_DO16}),
.DOPADOP({BRAM_L_X6Y140_RAMB18_X0Y56_DOP1, BRAM_L_X6Y140_RAMB18_X0Y56_DOP0}),
.DOPBDOP({BRAM_L_X6Y140_RAMB18_X0Y56_DOP3, BRAM_L_X6Y140_RAMB18_X0Y56_DOP2}),
.ENARDEN(1'b1),
.ENBWREN(1'b1),
.REGCEAREGCE(1'b0),
.REGCEB(1'b0),
.RSTRAMARSTRAM(1'b1),
.RSTRAMB(1'b1),
.RSTREGARSTREG(1'b1),
.RSTREGB(1'b1),
.WEA({1'b0, 1'b0}),
.WEBWE({1'b0})
  );


  (* KEEP, DONT_TOUCH, BEL = "RAMB18E1" *)
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .IS_CLKARDCLK_INVERTED(0),
    .IS_CLKBWRCLK_INVERTED(0),
    .IS_ENARDEN_INVERTED(0),
    .IS_ENBWREN_INVERTED(0),
    .IS_RSTRAMARSTRAM_INVERTED(1),
    .IS_RSTRAMB_INVERTED(1),
    .IS_RSTREGARSTREG_INVERTED(1),
    .IS_RSTREGB_INVERTED(1),
    .RAM_MODE("TDP"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(1)
  ) BRAM_L_X6Y140_RAMB18_X0Y57_RAMB18E1 (
.ADDRARDADDR({1'b0, 1'b0, CLBLM_R_X3Y138_SLICE_X3Y138_DO6, CLBLM_R_X5Y138_SLICE_X6Y138_DO6, CLBLL_L_X4Y139_SLICE_X5Y139_DO6, CLBLM_R_X5Y137_SLICE_X7Y137_DO6, CLBLM_R_X3Y138_SLICE_X3Y138_BO6, CLBLL_L_X4Y140_SLICE_X4Y140_AO6, CLBLM_R_X3Y138_SLICE_X3Y138_CO6, CLBLL_L_X4Y140_SLICE_X4Y140_BO6, 1'b0, 1'b0, 1'b0, 1'b0}),
.ADDRBWRADDR({1'b0, 1'b0, CLBLM_R_X5Y140_SLICE_X6Y140_DO6, CLBLM_R_X5Y139_SLICE_X7Y139_DO6, CLBLM_R_X7Y138_SLICE_X8Y138_DO6, CLBLM_R_X7Y140_SLICE_X8Y140_BO6, CLBLM_R_X5Y138_SLICE_X7Y138_CO6, CLBLM_R_X7Y140_SLICE_X8Y140_DO6, CLBLM_R_X7Y139_SLICE_X8Y139_AO6, CLBLL_L_X4Y139_SLICE_X4Y139_DO6, 1'b0, 1'b0, 1'b0, 1'b0}),
.CLKARDCLK(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CLKBWRCLK(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.DIADI({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
.DIBDI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
.DIPADIP({1'b0, 1'b0}),
.DIPBDIP({1'b1, 1'b1}),
.DOADO({BRAM_L_X6Y140_RAMB18_X0Y57_DOADO15, BRAM_L_X6Y140_RAMB18_X0Y57_DOADO14, BRAM_L_X6Y140_RAMB18_X0Y57_DOADO13, BRAM_L_X6Y140_RAMB18_X0Y57_DOADO12, BRAM_L_X6Y140_RAMB18_X0Y57_DOADO11, BRAM_L_X6Y140_RAMB18_X0Y57_DOADO10, BRAM_L_X6Y140_RAMB18_X0Y57_DOADO9, BRAM_L_X6Y140_RAMB18_X0Y57_DOADO8, BRAM_L_X6Y140_RAMB18_X0Y57_DOADO7, BRAM_L_X6Y140_RAMB18_X0Y57_DOADO6, BRAM_L_X6Y140_RAMB18_X0Y57_DOADO5, BRAM_L_X6Y140_RAMB18_X0Y57_DOADO4, BRAM_L_X6Y140_RAMB18_X0Y57_DOADO3, BRAM_L_X6Y140_RAMB18_X0Y57_DOADO2, BRAM_L_X6Y140_RAMB18_X0Y57_DOADO1, BRAM_L_X6Y140_RAMB18_X0Y57_DOADO0}),
.DOBDO({BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO15, BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO14, BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO13, BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO12, BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO11, BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO10, BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO9, BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO8, BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO7, BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO6, BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO5, BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO4, BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO3, BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO2, BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO1, BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO0}),
.DOPADOP({BRAM_L_X6Y140_RAMB18_X0Y57_DOPADOP1, BRAM_L_X6Y140_RAMB18_X0Y57_DOPADOP0}),
.DOPBDOP({BRAM_L_X6Y140_RAMB18_X0Y57_DOPBDOP1, BRAM_L_X6Y140_RAMB18_X0Y57_DOPBDOP0}),
.ENARDEN(1'b1),
.ENBWREN(1'b1),
.REGCEAREGCE(1'b0),
.REGCEB(1'b0),
.RSTRAMARSTRAM(1'b1),
.RSTRAMB(1'b1),
.RSTREGARSTREG(1'b1),
.RSTREGB(1'b1),
.WEA({1'b0, 1'b0}),
.WEBWE({1'b0})
  );


  (* KEEP, DONT_TOUCH, BEL = "RAMB18E1" *)
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .IS_CLKARDCLK_INVERTED(0),
    .IS_CLKBWRCLK_INVERTED(0),
    .IS_ENARDEN_INVERTED(0),
    .IS_ENBWREN_INVERTED(0),
    .IS_RSTRAMARSTRAM_INVERTED(1),
    .IS_RSTRAMB_INVERTED(1),
    .IS_RSTREGARSTREG_INVERTED(1),
    .IS_RSTREGB_INVERTED(1),
    .RAM_MODE("TDP"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(1)
  ) BRAM_R_X17Y135_RAMB18_X1Y54_RAMB18E1 (
.ADDRARDADDR({1'b0, 1'b0, CLBLM_L_X16Y136_SLICE_X22Y136_BO6, CLBLM_L_X16Y136_SLICE_X22Y136_CO6, CLBLM_R_X13Y135_SLICE_X18Y135_AO6, CLBLM_L_X16Y135_SLICE_X22Y135_CO6, CLBLM_L_X16Y135_SLICE_X22Y135_DO6, CLBLM_L_X16Y136_SLICE_X22Y136_DO6, CLBLM_R_X15Y135_SLICE_X21Y135_BO6, CLBLM_L_X12Y135_SLICE_X16Y135_AO6, 1'b0, 1'b0, 1'b0, 1'b0}),
.ADDRBWRADDR({1'b0, 1'b0, CLBLM_R_X7Y135_SLICE_X9Y135_DO6, CLBLM_L_X8Y135_SLICE_X11Y135_CO6, CLBLM_L_X8Y134_SLICE_X11Y134_DO6, CLBLM_L_X8Y135_SLICE_X11Y135_AO6, CLBLM_L_X8Y132_SLICE_X10Y132_AO6, CLBLM_L_X10Y134_SLICE_X12Y134_CO6, CLBLM_L_X8Y132_SLICE_X10Y132_BO6, CLBLM_L_X8Y133_SLICE_X11Y133_DO6, 1'b0, 1'b0, 1'b0, 1'b0}),
.CLKARDCLK(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CLKBWRCLK(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.DIADI({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
.DIBDI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
.DIPADIP({1'b0, 1'b0}),
.DIPBDIP({1'b1, 1'b1}),
.DOADO({BRAM_R_X17Y135_RAMB18_X1Y54_DO15, BRAM_R_X17Y135_RAMB18_X1Y54_DO14, BRAM_R_X17Y135_RAMB18_X1Y54_DO13, BRAM_R_X17Y135_RAMB18_X1Y54_DO12, BRAM_R_X17Y135_RAMB18_X1Y54_DO11, BRAM_R_X17Y135_RAMB18_X1Y54_DO10, BRAM_R_X17Y135_RAMB18_X1Y54_DO9, BRAM_R_X17Y135_RAMB18_X1Y54_DO8, BRAM_R_X17Y135_RAMB18_X1Y54_DO7, BRAM_R_X17Y135_RAMB18_X1Y54_DO6, BRAM_R_X17Y135_RAMB18_X1Y54_DO5, BRAM_R_X17Y135_RAMB18_X1Y54_DO4, BRAM_R_X17Y135_RAMB18_X1Y54_DO3, BRAM_R_X17Y135_RAMB18_X1Y54_DO2, BRAM_R_X17Y135_RAMB18_X1Y54_DO1, BRAM_R_X17Y135_RAMB18_X1Y54_DO0}),
.DOBDO({BRAM_R_X17Y135_RAMB18_X1Y54_DO31, BRAM_R_X17Y135_RAMB18_X1Y54_DO30, BRAM_R_X17Y135_RAMB18_X1Y54_DO29, BRAM_R_X17Y135_RAMB18_X1Y54_DO28, BRAM_R_X17Y135_RAMB18_X1Y54_DO27, BRAM_R_X17Y135_RAMB18_X1Y54_DO26, BRAM_R_X17Y135_RAMB18_X1Y54_DO25, BRAM_R_X17Y135_RAMB18_X1Y54_DO24, BRAM_R_X17Y135_RAMB18_X1Y54_DO23, BRAM_R_X17Y135_RAMB18_X1Y54_DO22, BRAM_R_X17Y135_RAMB18_X1Y54_DO21, BRAM_R_X17Y135_RAMB18_X1Y54_DO20, BRAM_R_X17Y135_RAMB18_X1Y54_DO19, BRAM_R_X17Y135_RAMB18_X1Y54_DO18, BRAM_R_X17Y135_RAMB18_X1Y54_DO17, BRAM_R_X17Y135_RAMB18_X1Y54_DO16}),
.DOPADOP({BRAM_R_X17Y135_RAMB18_X1Y54_DOP1, BRAM_R_X17Y135_RAMB18_X1Y54_DOP0}),
.DOPBDOP({BRAM_R_X17Y135_RAMB18_X1Y54_DOP3, BRAM_R_X17Y135_RAMB18_X1Y54_DOP2}),
.ENARDEN(1'b1),
.ENBWREN(1'b1),
.REGCEAREGCE(1'b0),
.REGCEB(1'b0),
.RSTRAMARSTRAM(1'b1),
.RSTRAMB(1'b1),
.RSTREGARSTREG(1'b1),
.RSTREGB(1'b1),
.WEA({1'b0, 1'b0}),
.WEBWE({1'b0})
  );


  (* KEEP, DONT_TOUCH, BEL = "RAMB18E1" *)
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .IS_CLKARDCLK_INVERTED(0),
    .IS_CLKBWRCLK_INVERTED(0),
    .IS_ENARDEN_INVERTED(0),
    .IS_ENBWREN_INVERTED(0),
    .IS_RSTRAMARSTRAM_INVERTED(1),
    .IS_RSTRAMB_INVERTED(1),
    .IS_RSTREGARSTREG_INVERTED(1),
    .IS_RSTREGB_INVERTED(1),
    .RAM_MODE("TDP"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(1)
  ) BRAM_R_X17Y135_RAMB18_X1Y55_RAMB18E1 (
.ADDRARDADDR({1'b0, 1'b0, CLBLM_R_X13Y136_SLICE_X18Y136_BO6, CLBLM_R_X11Y136_SLICE_X14Y136_DO6, CLBLM_R_X11Y135_SLICE_X14Y135_CO6, CLBLM_L_X10Y136_SLICE_X12Y136_CO6, CLBLM_L_X10Y134_SLICE_X12Y134_BO6, CLBLM_L_X12Y135_SLICE_X16Y135_BO6, CLBLM_R_X11Y135_SLICE_X14Y135_BO6, CLBLM_L_X10Y136_SLICE_X13Y136_DO6, 1'b0, 1'b0, 1'b0, 1'b0}),
.ADDRBWRADDR({1'b0, 1'b0, CLBLM_R_X7Y136_SLICE_X9Y136_CO6, CLBLM_L_X8Y135_SLICE_X10Y135_CO6, CLBLM_L_X8Y135_SLICE_X11Y135_DO6, CLBLM_L_X8Y133_SLICE_X10Y133_AO6, CLBLM_L_X8Y133_SLICE_X10Y133_BO6, CLBLM_L_X8Y135_SLICE_X10Y135_DO6, CLBLM_L_X8Y134_SLICE_X11Y134_BO6, CLBLM_L_X8Y133_SLICE_X11Y133_CO6, 1'b0, 1'b0, 1'b0, 1'b0}),
.CLKARDCLK(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CLKBWRCLK(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.DIADI({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
.DIBDI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
.DIPADIP({1'b0, 1'b0}),
.DIPBDIP({1'b1, 1'b1}),
.DOADO({BRAM_R_X17Y135_RAMB18_X1Y55_DOADO15, BRAM_R_X17Y135_RAMB18_X1Y55_DOADO14, BRAM_R_X17Y135_RAMB18_X1Y55_DOADO13, BRAM_R_X17Y135_RAMB18_X1Y55_DOADO12, BRAM_R_X17Y135_RAMB18_X1Y55_DOADO11, BRAM_R_X17Y135_RAMB18_X1Y55_DOADO10, BRAM_R_X17Y135_RAMB18_X1Y55_DOADO9, BRAM_R_X17Y135_RAMB18_X1Y55_DOADO8, BRAM_R_X17Y135_RAMB18_X1Y55_DOADO7, BRAM_R_X17Y135_RAMB18_X1Y55_DOADO6, BRAM_R_X17Y135_RAMB18_X1Y55_DOADO5, BRAM_R_X17Y135_RAMB18_X1Y55_DOADO4, BRAM_R_X17Y135_RAMB18_X1Y55_DOADO3, BRAM_R_X17Y135_RAMB18_X1Y55_DOADO2, BRAM_R_X17Y135_RAMB18_X1Y55_DOADO1, BRAM_R_X17Y135_RAMB18_X1Y55_DOADO0}),
.DOBDO({BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO15, BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO14, BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO13, BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO12, BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO11, BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO10, BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO9, BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO8, BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO7, BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO6, BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO5, BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO4, BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO3, BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO2, BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO1, BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO0}),
.DOPADOP({BRAM_R_X17Y135_RAMB18_X1Y55_DOPADOP1, BRAM_R_X17Y135_RAMB18_X1Y55_DOPADOP0}),
.DOPBDOP({BRAM_R_X17Y135_RAMB18_X1Y55_DOPBDOP1, BRAM_R_X17Y135_RAMB18_X1Y55_DOPBDOP0}),
.ENARDEN(1'b1),
.ENBWREN(1'b1),
.REGCEAREGCE(1'b0),
.REGCEB(1'b0),
.RSTRAMARSTRAM(1'b1),
.RSTRAMB(1'b1),
.RSTREGARSTREG(1'b1),
.RSTREGB(1'b1),
.WEA({1'b0, 1'b0}),
.WEBWE({1'b0})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X0Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X0Y131_DO5),
.O6(CLBLL_L_X2Y131_SLICE_X0Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X0Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X0Y131_CO5),
.O6(CLBLL_L_X2Y131_SLICE_X0Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X0Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X0Y131_BO5),
.O6(CLBLL_L_X2Y131_SLICE_X0Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X0Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X0Y131_AO5),
.O6(CLBLL_L_X2Y131_SLICE_X0Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y131_SLICE_X1Y131_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y131_SLICE_X1Y131_AO5),
.Q(CLBLL_L_X2Y131_SLICE_X1Y131_A5Q),
.R(LIOB33_X0Y147_IOB_X0Y148_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y131_SLICE_X1Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y131_SLICE_X1Y131_AO6),
.Q(CLBLL_L_X2Y131_SLICE_X1Y131_AQ),
.R(LIOB33_X0Y147_IOB_X0Y148_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y131_SLICE_X1Y131_B_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y131_SLICE_X1Y131_BO6),
.Q(CLBLL_L_X2Y131_SLICE_X1Y131_BQ),
.S(LIOB33_X0Y147_IOB_X0Y148_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X1Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X1Y131_DO5),
.O6(CLBLL_L_X2Y131_SLICE_X1Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X1Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X1Y131_CO5),
.O6(CLBLL_L_X2Y131_SLICE_X1Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8080808080808080)
  ) CLBLL_L_X2Y131_SLICE_X1Y131_BLUT (
.I0(CLBLM_R_X3Y129_SLICE_X2Y129_A5Q),
.I1(CLBLM_R_X3Y129_SLICE_X2Y129_AQ),
.I2(CLBLM_R_X3Y129_SLICE_X2Y129_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X1Y131_BO5),
.O6(CLBLL_L_X2Y131_SLICE_X1Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000600066ccc6ccc)
  ) CLBLL_L_X2Y131_SLICE_X1Y131_ALUT (
.I0(CLBLM_R_X3Y129_SLICE_X2Y129_A5Q),
.I1(CLBLL_L_X2Y131_SLICE_X1Y131_A5Q),
.I2(CLBLM_R_X3Y129_SLICE_X2Y129_BQ),
.I3(CLBLM_R_X3Y129_SLICE_X2Y129_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X1Y131_AO5),
.O6(CLBLL_L_X2Y131_SLICE_X1Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y132_SLICE_X0Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y132_SLICE_X0Y132_DO5),
.O6(CLBLL_L_X2Y132_SLICE_X0Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y132_SLICE_X0Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y132_SLICE_X0Y132_CO5),
.O6(CLBLL_L_X2Y132_SLICE_X0Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y132_SLICE_X0Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y132_SLICE_X0Y132_BO5),
.O6(CLBLL_L_X2Y132_SLICE_X0Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y132_SLICE_X0Y132_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y132_SLICE_X0Y132_AO5),
.O6(CLBLL_L_X2Y132_SLICE_X0Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y132_SLICE_X1Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y132_SLICE_X1Y132_AO6),
.Q(CLBLL_L_X2Y132_SLICE_X1Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y132_SLICE_X1Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y132_SLICE_X1Y132_DO5),
.O6(CLBLL_L_X2Y132_SLICE_X1Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y132_SLICE_X1Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y132_SLICE_X1Y132_CO5),
.O6(CLBLL_L_X2Y132_SLICE_X1Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y132_SLICE_X1Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y132_SLICE_X1Y132_BO5),
.O6(CLBLL_L_X2Y132_SLICE_X1Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff96ff9600960096)
  ) CLBLL_L_X2Y132_SLICE_X1Y132_ALUT (
.I0(CLBLM_R_X3Y132_SLICE_X2Y132_CQ),
.I1(CLBLM_R_X3Y132_SLICE_X2Y132_AO5),
.I2(CLBLL_L_X2Y132_SLICE_X1Y132_AQ),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X2Y132_SLICE_X1Y132_AO5),
.O6(CLBLL_L_X2Y132_SLICE_X1Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y141_SLICE_X0Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y141_SLICE_X0Y141_AO6),
.Q(CLBLL_L_X2Y141_SLICE_X0Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y141_SLICE_X0Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y141_SLICE_X0Y141_DO5),
.O6(CLBLL_L_X2Y141_SLICE_X0Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y141_SLICE_X0Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y141_SLICE_X0Y141_CO5),
.O6(CLBLL_L_X2Y141_SLICE_X0Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y141_SLICE_X0Y141_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y141_SLICE_X0Y141_BO5),
.O6(CLBLL_L_X2Y141_SLICE_X0Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000020002)
  ) CLBLL_L_X2Y141_SLICE_X0Y141_ALUT (
.I0(CLBLL_L_X2Y142_SLICE_X0Y142_DQ),
.I1(CLBLL_L_X2Y142_SLICE_X0Y142_BQ),
.I2(CLBLL_L_X2Y142_SLICE_X0Y142_AQ),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(1'b1),
.I5(CLBLL_L_X2Y142_SLICE_X0Y142_CQ),
.O5(CLBLL_L_X2Y141_SLICE_X0Y141_AO5),
.O6(CLBLL_L_X2Y141_SLICE_X0Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y141_SLICE_X1Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y141_SLICE_X1Y141_DO5),
.O6(CLBLL_L_X2Y141_SLICE_X1Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y141_SLICE_X1Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y141_SLICE_X1Y141_CO5),
.O6(CLBLL_L_X2Y141_SLICE_X1Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y141_SLICE_X1Y141_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y141_SLICE_X1Y141_BO5),
.O6(CLBLL_L_X2Y141_SLICE_X1Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y141_SLICE_X1Y141_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y141_SLICE_X1Y141_AO5),
.O6(CLBLL_L_X2Y141_SLICE_X1Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y142_SLICE_X0Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y142_SLICE_X0Y142_AO6),
.Q(CLBLL_L_X2Y142_SLICE_X0Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y142_SLICE_X0Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y142_SLICE_X0Y142_BO6),
.Q(CLBLL_L_X2Y142_SLICE_X0Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y142_SLICE_X0Y142_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y142_SLICE_X0Y142_CO6),
.Q(CLBLL_L_X2Y142_SLICE_X0Y142_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y142_SLICE_X0Y142_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y142_SLICE_X0Y142_DO6),
.Q(CLBLL_L_X2Y142_SLICE_X0Y142_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0a0a0a08)
  ) CLBLL_L_X2Y142_SLICE_X0Y142_DLUT (
.I0(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I1(CLBLL_L_X2Y142_SLICE_X0Y142_AQ),
.I2(CLBLL_L_X2Y142_SLICE_X0Y142_DQ),
.I3(CLBLL_L_X2Y142_SLICE_X0Y142_BQ),
.I4(CLBLL_L_X2Y142_SLICE_X0Y142_CQ),
.I5(LIOB33_X0Y147_IOB_X0Y148_I),
.O5(CLBLL_L_X2Y142_SLICE_X0Y142_DO5),
.O6(CLBLL_L_X2Y142_SLICE_X0Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaaaa80000)
  ) CLBLL_L_X2Y142_SLICE_X0Y142_CLUT (
.I0(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I1(CLBLL_L_X2Y142_SLICE_X0Y142_AQ),
.I2(CLBLL_L_X2Y142_SLICE_X0Y142_DQ),
.I3(CLBLL_L_X2Y142_SLICE_X0Y142_BQ),
.I4(CLBLL_L_X2Y142_SLICE_X0Y142_CQ),
.I5(LIOB33_X0Y147_IOB_X0Y148_I),
.O5(CLBLL_L_X2Y142_SLICE_X0Y142_CO5),
.O6(CLBLL_L_X2Y142_SLICE_X0Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000c0c00000c020)
  ) CLBLL_L_X2Y142_SLICE_X0Y142_BLUT (
.I0(CLBLL_L_X2Y142_SLICE_X0Y142_CQ),
.I1(CLBLL_L_X2Y142_SLICE_X0Y142_BQ),
.I2(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I3(CLBLL_L_X2Y142_SLICE_X0Y142_AQ),
.I4(LIOB33_X0Y147_IOB_X0Y148_I),
.I5(CLBLL_L_X2Y142_SLICE_X0Y142_DQ),
.O5(CLBLL_L_X2Y142_SLICE_X0Y142_BO5),
.O6(CLBLL_L_X2Y142_SLICE_X0Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff00000f0fe0000)
  ) CLBLL_L_X2Y142_SLICE_X0Y142_ALUT (
.I0(CLBLL_L_X2Y142_SLICE_X0Y142_CQ),
.I1(CLBLL_L_X2Y142_SLICE_X0Y142_BQ),
.I2(LIOB33_X0Y147_IOB_X0Y148_I),
.I3(CLBLL_L_X2Y142_SLICE_X0Y142_AQ),
.I4(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I5(CLBLL_L_X2Y142_SLICE_X0Y142_DQ),
.O5(CLBLL_L_X2Y142_SLICE_X0Y142_AO5),
.O6(CLBLL_L_X2Y142_SLICE_X0Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y142_SLICE_X1Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y142_SLICE_X1Y142_DO5),
.O6(CLBLL_L_X2Y142_SLICE_X1Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y142_SLICE_X1Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y142_SLICE_X1Y142_CO5),
.O6(CLBLL_L_X2Y142_SLICE_X1Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y142_SLICE_X1Y142_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y142_SLICE_X1Y142_BO5),
.O6(CLBLL_L_X2Y142_SLICE_X1Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y142_SLICE_X1Y142_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y142_SLICE_X1Y142_AO5),
.O6(CLBLL_L_X2Y142_SLICE_X1Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y152_SLICE_X0Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y187_IOB_X0Y187_I),
.Q(CLBLL_L_X2Y152_SLICE_X0Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y152_SLICE_X0Y152_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y152_SLICE_X0Y152_DO5),
.O6(CLBLL_L_X2Y152_SLICE_X0Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y152_SLICE_X0Y152_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y152_SLICE_X0Y152_CO5),
.O6(CLBLL_L_X2Y152_SLICE_X0Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y152_SLICE_X0Y152_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y152_SLICE_X0Y152_BO5),
.O6(CLBLL_L_X2Y152_SLICE_X0Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y152_SLICE_X0Y152_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y152_SLICE_X0Y152_AO5),
.O6(CLBLL_L_X2Y152_SLICE_X0Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y152_SLICE_X1Y152_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y152_SLICE_X1Y152_DO5),
.O6(CLBLL_L_X2Y152_SLICE_X1Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y152_SLICE_X1Y152_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y152_SLICE_X1Y152_CO5),
.O6(CLBLL_L_X2Y152_SLICE_X1Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y152_SLICE_X1Y152_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y152_SLICE_X1Y152_BO5),
.O6(CLBLL_L_X2Y152_SLICE_X1Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y152_SLICE_X1Y152_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y152_SLICE_X1Y152_AO5),
.O6(CLBLL_L_X2Y152_SLICE_X1Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y155_SLICE_X0Y155_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_SING_X0Y199_IOB_X0Y199_I),
.Q(CLBLL_L_X2Y155_SLICE_X0Y155_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y155_SLICE_X0Y155_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_SING_X0Y200_IOB_X0Y200_I),
.Q(CLBLL_L_X2Y155_SLICE_X0Y155_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y155_SLICE_X0Y155_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y203_IOB_X0Y203_I),
.Q(CLBLL_L_X2Y155_SLICE_X0Y155_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y155_SLICE_X0Y155_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y213_IOB_X0Y213_I),
.Q(CLBLL_L_X2Y155_SLICE_X0Y155_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y155_SLICE_X0Y155_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y155_SLICE_X0Y155_DO5),
.O6(CLBLL_L_X2Y155_SLICE_X0Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y155_SLICE_X0Y155_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y155_SLICE_X0Y155_CO5),
.O6(CLBLL_L_X2Y155_SLICE_X0Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y155_SLICE_X0Y155_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y155_SLICE_X0Y155_BO5),
.O6(CLBLL_L_X2Y155_SLICE_X0Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y155_SLICE_X0Y155_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y155_SLICE_X0Y155_AO5),
.O6(CLBLL_L_X2Y155_SLICE_X0Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y155_SLICE_X1Y155_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y195_IOB_X0Y195_I),
.Q(CLBLL_L_X2Y155_SLICE_X1Y155_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y155_SLICE_X1Y155_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y197_IOB_X0Y197_I),
.Q(CLBLL_L_X2Y155_SLICE_X1Y155_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y155_SLICE_X1Y155_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y155_SLICE_X1Y155_DO5),
.O6(CLBLL_L_X2Y155_SLICE_X1Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y155_SLICE_X1Y155_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y155_SLICE_X1Y155_CO5),
.O6(CLBLL_L_X2Y155_SLICE_X1Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y155_SLICE_X1Y155_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y155_SLICE_X1Y155_BO5),
.O6(CLBLL_L_X2Y155_SLICE_X1Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y155_SLICE_X1Y155_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y155_SLICE_X1Y155_AO5),
.O6(CLBLL_L_X2Y155_SLICE_X1Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y157_SLICE_X0Y157_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y209_IOB_X0Y210_I),
.Q(CLBLL_L_X2Y157_SLICE_X0Y157_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y157_SLICE_X0Y157_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y211_IOB_X0Y211_I),
.Q(CLBLL_L_X2Y157_SLICE_X0Y157_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y157_SLICE_X0Y157_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y211_IOB_X0Y212_I),
.Q(CLBLL_L_X2Y157_SLICE_X0Y157_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y157_SLICE_X0Y157_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y219_IOB_X0Y219_I),
.Q(CLBLL_L_X2Y157_SLICE_X0Y157_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y157_SLICE_X0Y157_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y157_SLICE_X0Y157_DO5),
.O6(CLBLL_L_X2Y157_SLICE_X0Y157_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y157_SLICE_X0Y157_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y157_SLICE_X0Y157_CO5),
.O6(CLBLL_L_X2Y157_SLICE_X0Y157_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y157_SLICE_X0Y157_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y157_SLICE_X0Y157_BO5),
.O6(CLBLL_L_X2Y157_SLICE_X0Y157_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y157_SLICE_X0Y157_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y157_SLICE_X0Y157_AO5),
.O6(CLBLL_L_X2Y157_SLICE_X0Y157_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y157_SLICE_X1Y157_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y203_IOB_X0Y204_I),
.Q(CLBLL_L_X2Y157_SLICE_X1Y157_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y157_SLICE_X1Y157_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y209_IOB_X0Y209_I),
.Q(CLBLL_L_X2Y157_SLICE_X1Y157_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y157_SLICE_X1Y157_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y157_SLICE_X1Y157_DO5),
.O6(CLBLL_L_X2Y157_SLICE_X1Y157_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y157_SLICE_X1Y157_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y157_SLICE_X1Y157_CO5),
.O6(CLBLL_L_X2Y157_SLICE_X1Y157_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y157_SLICE_X1Y157_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y157_SLICE_X1Y157_BO5),
.O6(CLBLL_L_X2Y157_SLICE_X1Y157_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y157_SLICE_X1Y157_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y157_SLICE_X1Y157_AO5),
.O6(CLBLL_L_X2Y157_SLICE_X1Y157_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y158_SLICE_X0Y158_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y207_IOB_X0Y208_I),
.Q(CLBLL_L_X2Y158_SLICE_X0Y158_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y158_SLICE_X0Y158_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y227_IOB_X0Y228_I),
.Q(CLBLL_L_X2Y158_SLICE_X0Y158_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y158_SLICE_X0Y158_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y229_IOB_X0Y229_I),
.Q(CLBLL_L_X2Y158_SLICE_X0Y158_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y158_SLICE_X0Y158_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y235_IOB_X0Y235_I),
.Q(CLBLL_L_X2Y158_SLICE_X0Y158_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y158_SLICE_X0Y158_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y158_SLICE_X0Y158_DO5),
.O6(CLBLL_L_X2Y158_SLICE_X0Y158_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y158_SLICE_X0Y158_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y158_SLICE_X0Y158_CO5),
.O6(CLBLL_L_X2Y158_SLICE_X0Y158_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y158_SLICE_X0Y158_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y158_SLICE_X0Y158_BO5),
.O6(CLBLL_L_X2Y158_SLICE_X0Y158_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y158_SLICE_X0Y158_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y158_SLICE_X0Y158_AO5),
.O6(CLBLL_L_X2Y158_SLICE_X0Y158_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y158_SLICE_X1Y158_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y158_SLICE_X1Y158_DO5),
.O6(CLBLL_L_X2Y158_SLICE_X1Y158_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y158_SLICE_X1Y158_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y158_SLICE_X1Y158_CO5),
.O6(CLBLL_L_X2Y158_SLICE_X1Y158_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y158_SLICE_X1Y158_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y158_SLICE_X1Y158_BO5),
.O6(CLBLL_L_X2Y158_SLICE_X1Y158_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y158_SLICE_X1Y158_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y158_SLICE_X1Y158_AO5),
.O6(CLBLL_L_X2Y158_SLICE_X1Y158_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y127_SLICE_X4Y127_DO5),
.O6(CLBLL_L_X4Y127_SLICE_X4Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y127_SLICE_X4Y127_CO5),
.O6(CLBLL_L_X4Y127_SLICE_X4Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y127_SLICE_X4Y127_BO5),
.O6(CLBLL_L_X4Y127_SLICE_X4Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y127_SLICE_X4Y127_AO5),
.O6(CLBLL_L_X4Y127_SLICE_X4Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y127_SLICE_X5Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y127_SLICE_X5Y127_AO6),
.Q(CLBLL_L_X4Y127_SLICE_X5Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y127_SLICE_X5Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y127_SLICE_X5Y127_DO5),
.O6(CLBLL_L_X4Y127_SLICE_X5Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y127_SLICE_X5Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y127_SLICE_X5Y127_CO5),
.O6(CLBLL_L_X4Y127_SLICE_X5Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3acaca3aca3a3ac)
  ) CLBLL_L_X4Y127_SLICE_X5Y127_BLUT (
.I0(LIOB33_SING_X0Y50_IOB_X0Y50_I),
.I1(CLBLL_L_X4Y128_SLICE_X5Y128_BQ),
.I2(LIOB33_X0Y147_IOB_X0Y148_I),
.I3(BRAM_L_X6Y125_RAMB18_X0Y50_DO7),
.I4(CLBLM_R_X5Y127_SLICE_X7Y127_DQ),
.I5(CLBLL_L_X4Y128_SLICE_X5Y128_AO5),
.O5(CLBLL_L_X4Y127_SLICE_X5Y127_BO5),
.O6(CLBLL_L_X4Y127_SLICE_X5Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdeed1221edde2112)
  ) CLBLL_L_X4Y127_SLICE_X5Y127_ALUT (
.I0(CLBLL_L_X4Y127_SLICE_X5Y127_AQ),
.I1(LIOB33_X0Y147_IOB_X0Y148_I),
.I2(CLBLM_R_X7Y129_SLICE_X9Y129_B5Q),
.I3(BRAM_L_X6Y125_RAMB18_X0Y50_DO6),
.I4(LIOB33_X0Y19_IOB_X0Y20_I),
.I5(CLBLM_R_X5Y127_SLICE_X6Y127_B5Q),
.O5(CLBLL_L_X4Y127_SLICE_X5Y127_AO5),
.O6(CLBLL_L_X4Y127_SLICE_X5Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y128_SLICE_X4Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y128_SLICE_X4Y128_DO5),
.O6(CLBLL_L_X4Y128_SLICE_X4Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y128_SLICE_X4Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y128_SLICE_X4Y128_CO5),
.O6(CLBLL_L_X4Y128_SLICE_X4Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y128_SLICE_X4Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y128_SLICE_X4Y128_BO5),
.O6(CLBLL_L_X4Y128_SLICE_X4Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y128_SLICE_X4Y128_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y128_SLICE_X4Y128_AO5),
.O6(CLBLL_L_X4Y128_SLICE_X4Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y128_SLICE_X5Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y128_SLICE_X5Y128_AO6),
.Q(CLBLL_L_X4Y128_SLICE_X5Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y128_SLICE_X5Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y128_SLICE_X5Y128_BO6),
.Q(CLBLL_L_X4Y128_SLICE_X5Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y128_SLICE_X5Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y128_SLICE_X5Y128_DO5),
.O6(CLBLL_L_X4Y128_SLICE_X5Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y128_SLICE_X5Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y128_SLICE_X5Y128_CO5),
.O6(CLBLL_L_X4Y128_SLICE_X5Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa3cc3aaaac33c)
  ) CLBLL_L_X4Y128_SLICE_X5Y128_BLUT (
.I0(LIOB33_X0Y21_IOB_X0Y21_I),
.I1(CLBLL_L_X4Y128_SLICE_X5Y128_BQ),
.I2(CLBLL_L_X4Y128_SLICE_X5Y128_AQ),
.I3(CLBLM_L_X8Y130_SLICE_X10Y130_A5Q),
.I4(LIOB33_X0Y147_IOB_X0Y148_I),
.I5(BRAM_L_X6Y125_RAMB18_X0Y50_DO7),
.O5(CLBLL_L_X4Y128_SLICE_X5Y128_BO5),
.O6(CLBLL_L_X4Y128_SLICE_X5Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff9600963c3c3c3c)
  ) CLBLL_L_X4Y128_SLICE_X5Y128_ALUT (
.I0(BRAM_L_X6Y125_RAMB18_X0Y50_DO7),
.I1(CLBLM_L_X8Y130_SLICE_X10Y130_A5Q),
.I2(CLBLL_L_X4Y128_SLICE_X5Y128_AQ),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(LIOB33_X0Y71_IOB_X0Y71_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y128_SLICE_X5Y128_AO5),
.O6(CLBLL_L_X4Y128_SLICE_X5Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y129_SLICE_X5Y129_BO6),
.Q(CLBLL_L_X4Y129_SLICE_X4Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y129_SLICE_X4Y129_DO5),
.O6(CLBLL_L_X4Y129_SLICE_X4Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y129_SLICE_X4Y129_CO5),
.O6(CLBLL_L_X4Y129_SLICE_X4Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y129_SLICE_X4Y129_BO5),
.O6(CLBLL_L_X4Y129_SLICE_X4Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y129_SLICE_X4Y129_AO5),
.O6(CLBLL_L_X4Y129_SLICE_X4Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y129_SLICE_X5Y129_AO6),
.Q(CLBLL_L_X4Y129_SLICE_X5Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y129_SLICE_X5Y129_CO6),
.Q(CLBLL_L_X4Y129_SLICE_X5Y129_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf6f9f9f606090906)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_DLUT (
.I0(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.I1(BRAM_L_X6Y125_RAMB18_X0Y50_DO18),
.I2(LIOB33_X0Y147_IOB_X0Y148_I),
.I3(CLBLL_L_X4Y129_SLICE_X5Y129_AO5),
.I4(CLBLL_L_X4Y129_SLICE_X5Y129_CQ),
.I5(LIOB33_X0Y9_IOB_X0Y9_I),
.O5(CLBLL_L_X4Y129_SLICE_X5Y129_DO5),
.O6(CLBLL_L_X4Y129_SLICE_X5Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb1e4e4b1e4b1b1e4)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_CLUT (
.I0(LIOB33_X0Y147_IOB_X0Y148_I),
.I1(BRAM_L_X6Y125_RAMB18_X0Y50_DO18),
.I2(LIOB33_X0Y23_IOB_X0Y24_I),
.I3(CLBLL_L_X4Y129_SLICE_X5Y129_AQ),
.I4(CLBLL_L_X4Y129_SLICE_X5Y129_CQ),
.I5(CLBLM_R_X7Y129_SLICE_X8Y129_B5Q),
.O5(CLBLL_L_X4Y129_SLICE_X5Y129_CO5),
.O6(CLBLL_L_X4Y129_SLICE_X5Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he2d1d1e25555aaaa)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_BLUT (
.I0(CLBLM_R_X7Y136_SLICE_X8Y136_A5Q),
.I1(LIOB33_X0Y147_IOB_X0Y148_I),
.I2(LIOB33_X0Y73_IOB_X0Y73_I),
.I3(BRAM_L_X6Y125_RAMB18_X0Y50_DO17),
.I4(CLBLL_L_X4Y129_SLICE_X4Y129_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y129_SLICE_X5Y129_BO5),
.O6(CLBLL_L_X4Y129_SLICE_X5Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haac3aa3c0f0ff0f0)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_ALUT (
.I0(LIOB33_X0Y73_IOB_X0Y74_I),
.I1(BRAM_L_X6Y125_RAMB18_X0Y50_DO18),
.I2(CLBLL_L_X4Y129_SLICE_X5Y129_AQ),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(CLBLM_R_X7Y129_SLICE_X8Y129_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y129_SLICE_X5Y129_AO5),
.O6(CLBLL_L_X4Y129_SLICE_X5Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y130_SLICE_X4Y130_BO6),
.Q(CLBLL_L_X4Y130_SLICE_X4Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf066f099f099f066)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_DLUT (
.I0(CLBLM_R_X3Y130_SLICE_X3Y130_BQ),
.I1(CLBLL_L_X4Y130_SLICE_X5Y130_A5Q),
.I2(LIOB33_X0Y11_IOB_X0Y12_I),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(CLBLM_R_X3Y130_SLICE_X3Y130_AO5),
.I5(BRAM_L_X6Y125_RAMB18_X0Y50_DO21),
.O5(CLBLL_L_X4Y130_SLICE_X4Y130_DO5),
.O6(CLBLL_L_X4Y130_SLICE_X4Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa3cc3c33c)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_CLUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(BRAM_L_X6Y130_RAMB18_X0Y52_DO2),
.I2(CLBLL_L_X4Y131_SLICE_X4Y131_BO5),
.I3(CLBLM_R_X5Y130_SLICE_X6Y130_DQ),
.I4(CLBLL_L_X4Y131_SLICE_X4Y131_DQ),
.I5(LIOB33_X0Y147_IOB_X0Y148_I),
.O5(CLBLL_L_X4Y130_SLICE_X4Y130_CO5),
.O6(CLBLL_L_X4Y130_SLICE_X4Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff699600006996)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_BLUT (
.I0(CLBLM_L_X8Y135_SLICE_X10Y135_A5Q),
.I1(CLBLL_L_X4Y130_SLICE_X4Y130_BQ),
.I2(CLBLL_L_X4Y131_SLICE_X4Y131_AQ),
.I3(BRAM_L_X6Y130_RAMB18_X0Y52_DO1),
.I4(LIOB33_X0Y147_IOB_X0Y148_I),
.I5(LIOB33_X0Y31_IOB_X0Y31_I),
.O5(CLBLL_L_X4Y130_SLICE_X4Y130_BO5),
.O6(CLBLL_L_X4Y130_SLICE_X4Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haca3a3ac3333cccc)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_ALUT (
.I0(LIOB33_X0Y81_IOB_X0Y81_I),
.I1(CLBLM_L_X8Y135_SLICE_X10Y135_A5Q),
.I2(LIOB33_X0Y147_IOB_X0Y148_I),
.I3(BRAM_L_X6Y130_RAMB18_X0Y52_DO1),
.I4(CLBLL_L_X4Y131_SLICE_X4Y131_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y130_SLICE_X4Y130_AO5),
.O6(CLBLL_L_X4Y130_SLICE_X4Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y130_SLICE_X4Y130_DO6),
.Q(CLBLL_L_X4Y130_SLICE_X5Y130_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y130_SLICE_X5Y130_AO6),
.Q(CLBLL_L_X4Y130_SLICE_X5Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y130_SLICE_X5Y130_DO6),
.Q(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf066f099f099f066)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_DLUT (
.I0(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I1(CLBLM_R_X3Y131_SLICE_X3Y131_AO5),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(CLBLL_L_X4Y130_SLICE_X5Y130_AQ),
.I5(CLBLM_R_X3Y131_SLICE_X3Y131_CQ),
.O5(CLBLL_L_X4Y130_SLICE_X5Y130_DO5),
.O6(CLBLL_L_X4Y130_SLICE_X5Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbeeb1441ebbe4114)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_CLUT (
.I0(LIOB33_X0Y147_IOB_X0Y148_I),
.I1(CLBLL_L_X4Y131_SLICE_X5Y131_CQ),
.I2(CLBLL_L_X4Y131_SLICE_X5Y131_AO5),
.I3(BRAM_L_X6Y125_RAMB18_X0Y50_DO22),
.I4(LIOB33_X0Y13_IOB_X0Y13_I),
.I5(CLBLM_R_X5Y130_SLICE_X6Y130_B5Q),
.O5(CLBLL_L_X4Y130_SLICE_X5Y130_CO5),
.O6(CLBLL_L_X4Y130_SLICE_X5Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf6f9f9f606090906)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_BLUT (
.I0(CLBLL_L_X4Y130_SLICE_X4Y130_AO5),
.I1(BRAM_L_X6Y130_RAMB18_X0Y52_DO1),
.I2(LIOB33_X0Y147_IOB_X0Y148_I),
.I3(CLBLL_L_X4Y130_SLICE_X4Y130_BQ),
.I4(CLBLM_R_X7Y130_SLICE_X8Y130_B5Q),
.I5(LIOB33_X0Y15_IOB_X0Y16_I),
.O5(CLBLL_L_X4Y130_SLICE_X5Y130_BO5),
.O6(CLBLL_L_X4Y130_SLICE_X5Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haac3aac3aa3caa3c)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_ALUT (
.I0(LIOB33_X0Y57_IOB_X0Y58_I),
.I1(CLBLM_R_X3Y131_SLICE_X3Y131_CQ),
.I2(CLBLL_L_X4Y130_SLICE_X5Y130_AQ),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(1'b1),
.I5(CLBLM_R_X3Y131_SLICE_X3Y131_AO5),
.O5(CLBLL_L_X4Y130_SLICE_X5Y130_AO5),
.O6(CLBLL_L_X4Y130_SLICE_X5Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y130_SLICE_X4Y130_AO6),
.Q(CLBLL_L_X4Y131_SLICE_X4Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.Q(CLBLL_L_X4Y131_SLICE_X4Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y131_SLICE_X4Y131_CO6),
.Q(CLBLL_L_X4Y131_SLICE_X4Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y131_SLICE_X4Y131_DO6),
.Q(CLBLL_L_X4Y131_SLICE_X4Y131_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc5acca5cca5cc5a)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_DLUT (
.I0(BRAM_L_X6Y130_RAMB18_X0Y52_DO2),
.I1(LIOB33_X0Y53_IOB_X0Y53_I),
.I2(CLBLL_L_X4Y131_SLICE_X4Y131_DQ),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(CLBLM_R_X7Y134_SLICE_X9Y134_A5Q),
.I5(CLBLL_L_X4Y131_SLICE_X4Y131_BQ),
.O5(CLBLL_L_X4Y131_SLICE_X4Y131_DO5),
.O6(CLBLL_L_X4Y131_SLICE_X4Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f06699f0f09966)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_CLUT (
.I0(CLBLL_L_X4Y132_SLICE_X4Y132_AQ),
.I1(CLBLL_L_X4Y131_SLICE_X4Y131_CQ),
.I2(LIOB33_X0Y89_IOB_X0Y89_I),
.I3(BRAM_L_X6Y130_RAMB18_X0Y52_DO17),
.I4(LIOB33_X0Y147_IOB_X0Y148_I),
.I5(CLBLM_R_X3Y131_SLICE_X2Y131_AQ),
.O5(CLBLL_L_X4Y131_SLICE_X4Y131_CO5),
.O6(CLBLL_L_X4Y131_SLICE_X4Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf909f60666666666)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_BLUT (
.I0(CLBLM_R_X7Y134_SLICE_X9Y134_A5Q),
.I1(CLBLL_L_X4Y131_SLICE_X4Y131_BQ),
.I2(LIOB33_X0Y147_IOB_X0Y148_I),
.I3(LIOB33_X0Y81_IOB_X0Y82_I),
.I4(BRAM_L_X6Y130_RAMB18_X0Y52_DO2),
.I5(1'b1),
.O5(CLBLL_L_X4Y131_SLICE_X4Y131_BO5),
.O6(CLBLL_L_X4Y131_SLICE_X4Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haac3aa3c0f0ff0f0)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_ALUT (
.I0(LIOB33_X0Y75_IOB_X0Y76_I),
.I1(BRAM_L_X6Y125_RAMB18_X0Y50_DO20),
.I2(CLBLM_R_X7Y132_SLICE_X8Y132_A5Q),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(CLBLL_L_X4Y131_SLICE_X5Y131_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y131_SLICE_X4Y131_AO5),
.O6(CLBLL_L_X4Y131_SLICE_X4Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y131_SLICE_X5Y131_AO6),
.Q(CLBLL_L_X4Y131_SLICE_X5Y131_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y131_SLICE_X4Y131_AO6),
.Q(CLBLL_L_X4Y131_SLICE_X5Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y131_SLICE_X5Y131_BO6),
.Q(CLBLL_L_X4Y131_SLICE_X5Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y131_SLICE_X5Y131_CO6),
.Q(CLBLL_L_X4Y131_SLICE_X5Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5aff005a5aff00)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_DLUT (
.I0(CLBLL_L_X4Y128_SLICE_X5Y128_AQ),
.I1(1'b1),
.I2(CLBLM_R_X3Y157_SLICE_X3Y157_DQ),
.I3(CLBLM_R_X5Y131_SLICE_X7Y131_DO6),
.I4(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y131_SLICE_X5Y131_DO5),
.O6(CLBLL_L_X4Y131_SLICE_X5Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa3caac3aac3aa3c)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_CLUT (
.I0(LIOB33_X0Y27_IOB_X0Y28_I),
.I1(CLBLL_L_X4Y131_SLICE_X5Y131_CQ),
.I2(BRAM_L_X6Y125_RAMB18_X0Y50_DO22),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(CLBLL_L_X4Y131_SLICE_X5Y131_B5Q),
.I5(CLBLM_R_X7Y137_SLICE_X8Y137_A5Q),
.O5(CLBLL_L_X4Y131_SLICE_X5Y131_CO5),
.O6(CLBLL_L_X4Y131_SLICE_X5Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa3cc3c33c)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_BLUT (
.I0(LIOB33_X0Y25_IOB_X0Y26_I),
.I1(CLBLL_L_X4Y131_SLICE_X5Y131_BQ),
.I2(CLBLL_L_X4Y131_SLICE_X5Y131_AQ),
.I3(BRAM_L_X6Y125_RAMB18_X0Y50_DO20),
.I4(CLBLM_R_X7Y132_SLICE_X8Y132_A5Q),
.I5(LIOB33_X0Y147_IOB_X0Y148_I),
.O5(CLBLL_L_X4Y131_SLICE_X5Y131_BO5),
.O6(CLBLL_L_X4Y131_SLICE_X5Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf9f6090666666666)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_ALUT (
.I0(CLBLL_L_X4Y131_SLICE_X5Y131_B5Q),
.I1(CLBLM_R_X7Y137_SLICE_X8Y137_A5Q),
.I2(LIOB33_X0Y147_IOB_X0Y148_I),
.I3(BRAM_L_X6Y125_RAMB18_X0Y50_DO22),
.I4(LIOB33_X0Y77_IOB_X0Y78_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y131_SLICE_X5Y131_AO5),
.O6(CLBLL_L_X4Y131_SLICE_X5Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y132_SLICE_X4Y132_AO6),
.Q(CLBLL_L_X4Y132_SLICE_X4Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y132_SLICE_X4Y132_BO6),
.Q(CLBLL_L_X4Y132_SLICE_X4Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y132_SLICE_X4Y132_CO6),
.Q(CLBLL_L_X4Y132_SLICE_X4Y132_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3acaca3aca3a3ac)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_DLUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(CLBLL_L_X4Y132_SLICE_X4Y132_BO5),
.I2(LIOB33_X0Y147_IOB_X0Y148_I),
.I3(CLBLL_L_X4Y133_SLICE_X4Y133_AQ),
.I4(BRAM_L_X6Y130_RAMB18_X0Y52_DO6),
.I5(CLBLM_R_X5Y132_SLICE_X7Y132_A5Q),
.O5(CLBLL_L_X4Y132_SLICE_X4Y132_DO5),
.O6(CLBLL_L_X4Y132_SLICE_X4Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haca3aca3a3aca3ac)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_CLUT (
.I0(LIOB33_X0Y57_IOB_X0Y57_I),
.I1(CLBLL_L_X4Y132_SLICE_X4Y132_CQ),
.I2(LIOB33_X0Y147_IOB_X0Y148_I),
.I3(CLBLL_L_X4Y132_SLICE_X4Y132_AO5),
.I4(1'b1),
.I5(CLBLL_L_X4Y131_SLICE_X4Y131_CQ),
.O5(CLBLL_L_X4Y132_SLICE_X4Y132_CO5),
.O6(CLBLL_L_X4Y132_SLICE_X4Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0996633cc33cc)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_BLUT (
.I0(BRAM_L_X6Y130_RAMB18_X0Y52_DO6),
.I1(CLBLL_L_X4Y132_SLICE_X4Y132_BQ),
.I2(LIOB33_X0Y85_IOB_X0Y86_I),
.I3(CLBLM_L_X8Y137_SLICE_X10Y137_A5Q),
.I4(LIOB33_X0Y147_IOB_X0Y148_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y132_SLICE_X4Y132_BO5),
.O6(CLBLL_L_X4Y132_SLICE_X4Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaac33cc33cc33c)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_ALUT (
.I0(LIOB33_X0Y141_IOB_X0Y141_I),
.I1(BRAM_L_X6Y130_RAMB18_X0Y52_DO17),
.I2(CLBLL_L_X4Y132_SLICE_X4Y132_AQ),
.I3(CLBLM_R_X3Y131_SLICE_X2Y131_AQ),
.I4(LIOB33_X0Y147_IOB_X0Y148_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y132_SLICE_X4Y132_AO5),
.O6(CLBLL_L_X4Y132_SLICE_X4Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y133_SLICE_X5Y133_CO6),
.Q(CLBLL_L_X4Y132_SLICE_X5Y132_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y132_SLICE_X5Y132_AO6),
.Q(CLBLL_L_X4Y132_SLICE_X5Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y132_SLICE_X5Y132_BO6),
.Q(CLBLL_L_X4Y132_SLICE_X5Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000069966996)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_DLUT (
.I0(CLBLL_L_X4Y131_SLICE_X4Y131_CQ),
.I1(CLBLL_L_X4Y132_SLICE_X4Y132_AO5),
.I2(CLBLM_R_X5Y132_SLICE_X6Y132_B5Q),
.I3(CLBLL_L_X4Y132_SLICE_X4Y132_CQ),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(LIOB33_X0Y147_IOB_X0Y148_I),
.O5(CLBLL_L_X4Y132_SLICE_X5Y132_DO5),
.O6(CLBLL_L_X4Y132_SLICE_X5Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff690069ff960096)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_CLUT (
.I0(CLBLL_L_X2Y132_SLICE_X1Y132_AQ),
.I1(CLBLM_R_X5Y132_SLICE_X7Y132_B5Q),
.I2(CLBLM_R_X3Y132_SLICE_X2Y132_CQ),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(CLBLM_R_X3Y132_SLICE_X2Y132_AO5),
.O5(CLBLL_L_X4Y132_SLICE_X5Y132_CO5),
.O6(CLBLL_L_X4Y132_SLICE_X5Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb1e4e4b1e4b1b1e4)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_BLUT (
.I0(LIOB33_X0Y147_IOB_X0Y148_I),
.I1(CLBLL_L_X4Y132_SLICE_X5Y132_BQ),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(CLBLM_R_X3Y132_SLICE_X2Y132_DQ),
.I4(CLBLM_R_X3Y132_SLICE_X3Y132_CQ),
.I5(CLBLM_R_X3Y132_SLICE_X2Y132_BO5),
.O5(CLBLL_L_X4Y132_SLICE_X5Y132_BO5),
.O6(CLBLL_L_X4Y132_SLICE_X5Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000069966996)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_ALUT (
.I0(BRAM_L_X6Y130_RAMB18_X0Y52_DO5),
.I1(CLBLM_R_X5Y132_SLICE_X6Y132_AQ),
.I2(CLBLL_L_X4Y132_SLICE_X5Y132_AQ),
.I3(CLBLM_L_X10Y135_SLICE_X12Y135_A5Q),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(LIOB33_X0Y147_IOB_X0Y148_I),
.O5(CLBLL_L_X4Y132_SLICE_X5Y132_AO5),
.O6(CLBLL_L_X4Y132_SLICE_X5Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y133_SLICE_X4Y133_CO6),
.Q(CLBLL_L_X4Y133_SLICE_X4Y133_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y133_SLICE_X4Y133_AO6),
.Q(CLBLL_L_X4Y133_SLICE_X4Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y133_SLICE_X4Y133_BO6),
.Q(CLBLL_L_X4Y133_SLICE_X4Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y133_SLICE_X4Y133_DO5),
.O6(CLBLL_L_X4Y133_SLICE_X4Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdeededde12212112)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_CLUT (
.I0(CLBLL_L_X4Y133_SLICE_X4Y133_BQ),
.I1(LIOB33_X0Y147_IOB_X0Y148_I),
.I2(CLBLM_R_X3Y132_SLICE_X3Y132_BQ),
.I3(CLBLL_L_X4Y133_SLICE_X4Y133_A5Q),
.I4(CLBLM_R_X3Y133_SLICE_X3Y133_AO5),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLL_L_X4Y133_SLICE_X4Y133_CO5),
.O6(CLBLL_L_X4Y133_SLICE_X4Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf099f099f066f066)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_BLUT (
.I0(CLBLM_R_X3Y133_SLICE_X3Y133_AO5),
.I1(CLBLL_L_X4Y133_SLICE_X4Y133_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y61_I),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(1'b1),
.I5(CLBLM_R_X3Y132_SLICE_X3Y132_BQ),
.O5(CLBLL_L_X4Y133_SLICE_X4Y133_BO5),
.O6(CLBLL_L_X4Y133_SLICE_X4Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc5aa5a55a)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_ALUT (
.I0(CLBLM_L_X8Y137_SLICE_X10Y137_A5Q),
.I1(LIOB33_X0Y117_IOB_X0Y118_I),
.I2(CLBLL_L_X4Y133_SLICE_X4Y133_AQ),
.I3(CLBLL_L_X4Y132_SLICE_X4Y132_BQ),
.I4(BRAM_L_X6Y130_RAMB18_X0Y52_DO6),
.I5(LIOB33_X0Y147_IOB_X0Y148_I),
.O5(CLBLL_L_X4Y133_SLICE_X4Y133_AO5),
.O6(CLBLL_L_X4Y133_SLICE_X4Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y133_SLICE_X5Y133_AO6),
.Q(CLBLL_L_X4Y133_SLICE_X5Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y133_SLICE_X5Y133_BO6),
.Q(CLBLL_L_X4Y133_SLICE_X5Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff69ff9600690096)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_DLUT (
.I0(CLBLM_R_X5Y133_SLICE_X6Y133_BQ),
.I1(CLBLM_R_X3Y132_SLICE_X3Y132_AO5),
.I2(CLBLM_R_X3Y131_SLICE_X3Y131_DQ),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(CLBLM_R_X3Y133_SLICE_X3Y133_BQ),
.I5(LIOB33_X0Y111_IOB_X0Y111_I),
.O5(CLBLL_L_X4Y133_SLICE_X5Y133_DO5),
.O6(CLBLL_L_X4Y133_SLICE_X5Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdeed1221edde2112)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_CLUT (
.I0(BRAM_L_X6Y130_RAMB18_X0Y52_DO7),
.I1(LIOB33_X0Y147_IOB_X0Y148_I),
.I2(CLBLL_L_X4Y133_SLICE_X5Y133_BQ),
.I3(CLBLL_L_X4Y133_SLICE_X5Y133_AO5),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLL_L_X4Y132_SLICE_X5Y132_A5Q),
.O5(CLBLL_L_X4Y133_SLICE_X5Y133_CO5),
.O6(CLBLL_L_X4Y133_SLICE_X5Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa3cc3c33c)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_BLUT (
.I0(LIOB33_X0Y55_IOB_X0Y55_I),
.I1(CLBLL_L_X4Y133_SLICE_X5Y133_BQ),
.I2(CLBLL_L_X4Y133_SLICE_X5Y133_AQ),
.I3(CLBLM_L_X8Y137_SLICE_X10Y137_B5Q),
.I4(BRAM_L_X6Y130_RAMB18_X0Y52_DO7),
.I5(LIOB33_X0Y147_IOB_X0Y148_I),
.O5(CLBLL_L_X4Y133_SLICE_X5Y133_BO5),
.O6(CLBLL_L_X4Y133_SLICE_X5Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hebbe41143c3c3c3c)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_ALUT (
.I0(LIOB33_X0Y147_IOB_X0Y148_I),
.I1(CLBLM_L_X8Y137_SLICE_X10Y137_B5Q),
.I2(CLBLL_L_X4Y133_SLICE_X5Y133_AQ),
.I3(BRAM_L_X6Y130_RAMB18_X0Y52_DO7),
.I4(LIOB33_X0Y87_IOB_X0Y87_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y133_SLICE_X5Y133_AO5),
.O6(CLBLL_L_X4Y133_SLICE_X5Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y134_SLICE_X3Y134_AO6),
.Q(CLBLL_L_X4Y134_SLICE_X4Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y134_SLICE_X4Y134_DO5),
.O6(CLBLL_L_X4Y134_SLICE_X4Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y134_SLICE_X4Y134_CO5),
.O6(CLBLL_L_X4Y134_SLICE_X4Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y134_SLICE_X4Y134_BO5),
.O6(CLBLL_L_X4Y134_SLICE_X4Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y134_SLICE_X4Y134_AO5),
.O6(CLBLL_L_X4Y134_SLICE_X4Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y134_SLICE_X5Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y134_SLICE_X5Y134_AO6),
.Q(CLBLL_L_X4Y134_SLICE_X5Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y134_SLICE_X5Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y134_SLICE_X5Y134_BO6),
.Q(CLBLL_L_X4Y134_SLICE_X5Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f0c0cf3f3c0c0)
  ) CLBLL_L_X4Y134_SLICE_X5Y134_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I2(CLBLM_R_X3Y147_SLICE_X2Y147_DQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y134_SLICE_X6Y134_CO6),
.I5(CLBLL_L_X4Y132_SLICE_X5Y132_A5Q),
.O5(CLBLL_L_X4Y134_SLICE_X5Y134_DO5),
.O6(CLBLL_L_X4Y134_SLICE_X5Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h553caac355c3aa3c)
  ) CLBLL_L_X4Y134_SLICE_X5Y134_CLUT (
.I0(CLBLL_L_X4Y145_SLICE_X4Y145_AQ),
.I1(CLBLL_L_X4Y135_SLICE_X5Y135_AO6),
.I2(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO0),
.I3(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I4(CLBLM_R_X5Y130_SLICE_X6Y130_CQ),
.I5(CLBLM_R_X5Y134_SLICE_X6Y134_AO6),
.O5(CLBLL_L_X4Y134_SLICE_X5Y134_CO5),
.O6(CLBLL_L_X4Y134_SLICE_X5Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0ff0f00f0ff0f0)
  ) CLBLL_L_X4Y134_SLICE_X5Y134_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X2Y132_SLICE_X1Y132_AQ),
.I3(1'b1),
.I4(BRAM_L_X6Y140_RAMB18_X0Y56_DO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y134_SLICE_X5Y134_BO5),
.O6(CLBLL_L_X4Y134_SLICE_X5Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff00ff00ff00ff0)
  ) CLBLL_L_X4Y134_SLICE_X5Y134_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X4Y133_SLICE_X5Y133_BQ),
.I3(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO7),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y134_SLICE_X5Y134_AO5),
.O6(CLBLL_L_X4Y134_SLICE_X5Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7b7b7b7b48484848)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_DLUT (
.I0(CLBLL_L_X4Y133_SLICE_X4Y133_AQ),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I2(CLBLL_L_X2Y157_SLICE_X1Y157_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X4Y135_SLICE_X4Y135_BO6),
.O5(CLBLL_L_X4Y135_SLICE_X4Y135_DO5),
.O6(CLBLL_L_X4Y135_SLICE_X4Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h09f9f90906f6f606)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_CLUT (
.I0(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO7),
.I1(CLBLL_L_X4Y135_SLICE_X5Y135_CO6),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I3(CLBLM_R_X5Y131_SLICE_X7Y131_CQ),
.I4(CLBLM_R_X3Y155_SLICE_X3Y155_CQ),
.I5(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO7),
.O5(CLBLL_L_X4Y135_SLICE_X4Y135_CO5),
.O6(CLBLL_L_X4Y135_SLICE_X4Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_BLUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y56_DO6),
.I1(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO5),
.I2(CLBLL_L_X4Y133_SLICE_X4Y133_AQ),
.I3(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO5),
.I4(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO6),
.I5(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO6),
.O5(CLBLL_L_X4Y135_SLICE_X4Y135_BO5),
.O6(CLBLL_L_X4Y135_SLICE_X4Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5a5555aaaa)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_ALUT (
.I0(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO0),
.I1(1'b1),
.I2(BRAM_L_X6Y140_RAMB18_X0Y56_DO0),
.I3(1'b1),
.I4(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y135_SLICE_X4Y135_AO5),
.O6(CLBLL_L_X4Y135_SLICE_X4Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y135_SLICE_X5Y135_BO6),
.Q(CLBLL_L_X4Y135_SLICE_X5Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c663c993c993c66)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_DLUT (
.I0(CLBLL_L_X4Y135_SLICE_X5Y135_AO6),
.I1(CLBLM_R_X5Y130_SLICE_X7Y130_CQ),
.I2(CLBLM_R_X3Y141_SLICE_X2Y141_CQ),
.I3(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I4(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO0),
.I5(CLBLM_R_X5Y134_SLICE_X6Y134_BO6),
.O5(CLBLL_L_X4Y135_SLICE_X5Y135_DO5),
.O6(CLBLL_L_X4Y135_SLICE_X5Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_CLUT (
.I0(CLBLM_R_X5Y131_SLICE_X7Y131_CQ),
.I1(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO3),
.I2(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO4),
.I3(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO3),
.I4(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO4),
.I5(BRAM_L_X6Y140_RAMB18_X0Y56_DO4),
.O5(CLBLL_L_X4Y135_SLICE_X5Y135_CO5),
.O6(CLBLL_L_X4Y135_SLICE_X5Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3c3c3c3c3c)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y133_SLICE_X4Y133_BQ),
.I2(BRAM_L_X6Y140_RAMB18_X0Y56_DO5),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y135_SLICE_X5Y135_BO5),
.O6(CLBLL_L_X4Y135_SLICE_X5Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6666666655aa55aa)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_ALUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO0),
.I1(BRAM_L_X6Y140_RAMB18_X0Y56_DO16),
.I2(1'b1),
.I3(CLBLM_R_X5Y127_SLICE_X6Y127_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y135_SLICE_X5Y135_AO5),
.O6(CLBLL_L_X4Y135_SLICE_X5Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y136_SLICE_X4Y136_DO5),
.O6(CLBLL_L_X4Y136_SLICE_X4Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa55aac3c33c3c)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_CLUT (
.I0(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.I1(CLBLL_L_X4Y136_SLICE_X4Y136_BO6),
.I2(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO7),
.I3(CLBLM_R_X3Y153_SLICE_X2Y153_DQ),
.I4(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO7),
.I5(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.O5(CLBLL_L_X4Y136_SLICE_X4Y136_CO5),
.O6(CLBLL_L_X4Y136_SLICE_X4Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_BLUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y56_DO3),
.I1(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO3),
.I2(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO2),
.I3(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.I4(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO3),
.I5(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO2),
.O5(CLBLL_L_X4Y136_SLICE_X4Y136_BO5),
.O6(CLBLL_L_X4Y136_SLICE_X4Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_ALUT (
.I0(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO6),
.I1(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO6),
.I2(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO5),
.I3(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO6),
.I4(CLBLL_L_X2Y132_SLICE_X1Y132_AQ),
.I5(BRAM_L_X6Y140_RAMB18_X0Y56_DO5),
.O5(CLBLL_L_X4Y136_SLICE_X4Y136_AO5),
.O6(CLBLL_L_X4Y136_SLICE_X4Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h77bb77bb44884488)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_DLUT (
.I0(CLBLM_R_X3Y153_SLICE_X2Y153_CQ),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y129_SLICE_X5Y129_CQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y136_SLICE_X5Y136_BO6),
.O5(CLBLL_L_X4Y136_SLICE_X5Y136_DO5),
.O6(CLBLL_L_X4Y136_SLICE_X5Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33aa33aaccaaccaa)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_CLUT (
.I0(CLBLM_R_X5Y136_SLICE_X6Y136_CO6),
.I1(CLBLM_R_X3Y141_SLICE_X2Y141_BQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.O5(CLBLL_L_X4Y136_SLICE_X5Y136_CO5),
.O6(CLBLL_L_X4Y136_SLICE_X5Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_BLUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y56_DO2),
.I1(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO2),
.I2(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO1),
.I3(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO1),
.I4(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO2),
.I5(CLBLL_L_X4Y129_SLICE_X5Y129_CQ),
.O5(CLBLL_L_X4Y136_SLICE_X5Y136_BO5),
.O6(CLBLL_L_X4Y136_SLICE_X5Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_ALUT (
.I0(CLBLM_R_X5Y129_SLICE_X6Y129_AQ),
.I1(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO2),
.I2(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO3),
.I3(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO3),
.I4(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO3),
.I5(BRAM_L_X6Y140_RAMB18_X0Y56_DO2),
.O5(CLBLL_L_X4Y136_SLICE_X5Y136_AO5),
.O6(CLBLL_L_X4Y136_SLICE_X5Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLL_L_X4Y137_SLICE_X4Y137_DLUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y56_DO0),
.I1(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO0),
.I2(BRAM_L_X6Y140_RAMB18_X0Y56_DO1),
.I3(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO1),
.I4(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO1),
.I5(CLBLM_R_X5Y125_SLICE_X7Y125_CQ),
.O5(CLBLL_L_X4Y137_SLICE_X4Y137_DO5),
.O6(CLBLL_L_X4Y137_SLICE_X4Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h35ca3ac53ac535ca)
  ) CLBLL_L_X4Y137_SLICE_X4Y137_CLUT (
.I0(CLBLL_L_X4Y135_SLICE_X4Y135_AO6),
.I1(CLBLM_R_X3Y155_SLICE_X3Y155_BQ),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I3(CLBLM_R_X5Y131_SLICE_X6Y131_CQ),
.I4(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO0),
.I5(CLBLM_R_X3Y137_SLICE_X3Y137_AO6),
.O5(CLBLL_L_X4Y137_SLICE_X4Y137_CO5),
.O6(CLBLL_L_X4Y137_SLICE_X4Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLL_L_X4Y137_SLICE_X4Y137_BLUT (
.I0(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO1),
.I1(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO2),
.I2(CLBLL_L_X4Y131_SLICE_X4Y131_DQ),
.I3(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO1),
.I4(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO2),
.I5(BRAM_L_X6Y140_RAMB18_X0Y56_DO2),
.O5(CLBLL_L_X4Y137_SLICE_X4Y137_BO5),
.O6(CLBLL_L_X4Y137_SLICE_X4Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLL_L_X4Y137_SLICE_X4Y137_ALUT (
.I0(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO1),
.I1(BRAM_L_X6Y140_RAMB18_X0Y56_DO0),
.I2(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO0),
.I3(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO1),
.I4(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO1),
.I5(CLBLL_L_X4Y132_SLICE_X4Y132_CQ),
.O5(CLBLL_L_X4Y137_SLICE_X4Y137_AO5),
.O6(CLBLL_L_X4Y137_SLICE_X4Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cc33cc69699696)
  ) CLBLL_L_X4Y137_SLICE_X5Y137_DLUT (
.I0(CLBLL_L_X4Y137_SLICE_X5Y137_AO6),
.I1(CLBLM_R_X5Y129_SLICE_X7Y129_BQ),
.I2(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO0),
.I3(CLBLM_R_X3Y153_SLICE_X2Y153_AQ),
.I4(CLBLL_L_X4Y135_SLICE_X4Y135_AO6),
.I5(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.O5(CLBLL_L_X4Y137_SLICE_X5Y137_DO5),
.O6(CLBLL_L_X4Y137_SLICE_X5Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5acc3333cc)
  ) CLBLL_L_X4Y137_SLICE_X5Y137_CLUT (
.I0(CLBLL_L_X4Y155_SLICE_X4Y155_AQ),
.I1(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO7),
.I2(CLBLL_L_X4Y131_SLICE_X5Y131_BQ),
.I3(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO7),
.I4(CLBLL_L_X4Y137_SLICE_X5Y137_BO6),
.I5(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.O5(CLBLL_L_X4Y137_SLICE_X5Y137_CO5),
.O6(CLBLL_L_X4Y137_SLICE_X5Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLL_L_X4Y137_SLICE_X5Y137_BLUT (
.I0(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO3),
.I1(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO3),
.I2(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO4),
.I3(BRAM_L_X6Y140_RAMB18_X0Y56_DO4),
.I4(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO4),
.I5(CLBLL_L_X4Y131_SLICE_X5Y131_BQ),
.O5(CLBLL_L_X4Y137_SLICE_X5Y137_BO5),
.O6(CLBLL_L_X4Y137_SLICE_X5Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa55aa0ff00ff0)
  ) CLBLL_L_X4Y137_SLICE_X5Y137_ALUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO7),
.I1(1'b1),
.I2(CLBLL_L_X4Y128_SLICE_X5Y128_BQ),
.I3(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO7),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y137_SLICE_X5Y137_AO5),
.O6(CLBLL_L_X4Y137_SLICE_X5Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLL_L_X4Y138_SLICE_X4Y138_DLUT (
.I0(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO1),
.I1(BRAM_L_X6Y140_RAMB18_X0Y56_DO2),
.I2(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.I3(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO2),
.I4(BRAM_L_X6Y140_RAMB18_X0Y56_DO1),
.I5(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO2),
.O5(CLBLL_L_X4Y138_SLICE_X4Y138_DO5),
.O6(CLBLL_L_X4Y138_SLICE_X4Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLL_L_X4Y138_SLICE_X4Y138_CLUT (
.I0(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO2),
.I1(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO3),
.I2(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO3),
.I3(BRAM_L_X6Y140_RAMB18_X0Y56_DO2),
.I4(BRAM_L_X6Y140_RAMB18_X0Y56_DO3),
.I5(CLBLM_R_X5Y126_SLICE_X6Y126_BQ),
.O5(CLBLL_L_X4Y138_SLICE_X4Y138_CO5),
.O6(CLBLL_L_X4Y138_SLICE_X4Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff00ff099996666)
  ) CLBLL_L_X4Y138_SLICE_X4Y138_BLUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO7),
.I1(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO7),
.I2(CLBLL_L_X2Y155_SLICE_X0Y155_AQ),
.I3(CLBLL_L_X4Y130_SLICE_X4Y130_BQ),
.I4(CLBLL_L_X4Y138_SLICE_X4Y138_AO6),
.I5(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.O5(CLBLL_L_X4Y138_SLICE_X4Y138_BO5),
.O6(CLBLL_L_X4Y138_SLICE_X4Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLL_L_X4Y138_SLICE_X4Y138_ALUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y56_DO1),
.I1(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO1),
.I2(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO1),
.I3(CLBLL_L_X4Y130_SLICE_X4Y130_BQ),
.I4(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO0),
.I5(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO0),
.O5(CLBLL_L_X4Y138_SLICE_X4Y138_AO5),
.O6(CLBLL_L_X4Y138_SLICE_X4Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_DLUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO5),
.I1(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO4),
.I2(CLBLM_R_X5Y127_SLICE_X7Y127_BQ),
.I3(BRAM_L_X6Y140_RAMB18_X0Y56_DO4),
.I4(BRAM_L_X6Y140_RAMB18_X0Y56_DO5),
.I5(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO5),
.O5(CLBLL_L_X4Y138_SLICE_X5Y138_DO5),
.O6(CLBLL_L_X4Y138_SLICE_X5Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_CLUT (
.I0(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO2),
.I1(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO2),
.I2(BRAM_L_X6Y140_RAMB18_X0Y56_DO1),
.I3(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO1),
.I4(CLBLL_L_X4Y130_SLICE_X5Y130_AQ),
.I5(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO2),
.O5(CLBLL_L_X4Y138_SLICE_X5Y138_CO5),
.O6(CLBLL_L_X4Y138_SLICE_X5Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_BLUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO4),
.I1(BRAM_L_X6Y140_RAMB18_X0Y56_DO3),
.I2(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO4),
.I3(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO3),
.I4(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO4),
.I5(CLBLM_R_X3Y133_SLICE_X3Y133_BQ),
.O5(CLBLL_L_X4Y138_SLICE_X5Y138_BO5),
.O6(CLBLL_L_X4Y138_SLICE_X5Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_ALUT (
.I0(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO5),
.I1(CLBLL_L_X4Y133_SLICE_X4Y133_BQ),
.I2(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO4),
.I3(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO5),
.I4(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO5),
.I5(BRAM_L_X6Y140_RAMB18_X0Y56_DO4),
.O5(CLBLL_L_X4Y138_SLICE_X5Y138_AO5),
.O6(CLBLL_L_X4Y138_SLICE_X5Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f0cf3c03f0cf3c0)
  ) CLBLL_L_X4Y139_SLICE_X4Y139_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I2(CLBLM_R_X5Y127_SLICE_X6Y127_CQ),
.I3(CLBLL_L_X4Y139_SLICE_X5Y139_BO6),
.I4(CLBLM_R_X3Y141_SLICE_X2Y141_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y139_SLICE_X4Y139_DO5),
.O6(CLBLL_L_X4Y139_SLICE_X4Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLL_L_X4Y139_SLICE_X4Y139_CLUT (
.I0(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO7),
.I1(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO0),
.I2(BRAM_L_X6Y140_RAMB18_X0Y56_DO7),
.I3(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO0),
.I4(BRAM_L_X6Y140_RAMB18_X0Y56_DO0),
.I5(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.O5(CLBLL_L_X4Y139_SLICE_X4Y139_CO5),
.O6(CLBLL_L_X4Y139_SLICE_X4Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h72d8278d278d72d8)
  ) CLBLL_L_X4Y139_SLICE_X4Y139_BLUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I1(CLBLL_L_X4Y132_SLICE_X4Y132_CQ),
.I2(CLBLL_L_X4Y137_SLICE_X4Y137_AO6),
.I3(CLBLL_L_X4Y156_SLICE_X4Y156_AQ),
.I4(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO7),
.I5(BRAM_L_X6Y140_RAMB18_X0Y56_DO7),
.O5(CLBLL_L_X4Y139_SLICE_X4Y139_BO5),
.O6(CLBLL_L_X4Y139_SLICE_X4Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h41eb14beeb41be14)
  ) CLBLL_L_X4Y139_SLICE_X4Y139_ALUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I1(CLBLL_L_X4Y136_SLICE_X5Y136_AO6),
.I2(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO7),
.I3(CLBLL_L_X2Y157_SLICE_X1Y157_BQ),
.I4(BRAM_L_X6Y140_RAMB18_X0Y56_DO7),
.I5(CLBLM_R_X5Y129_SLICE_X6Y129_AQ),
.O5(CLBLL_L_X4Y139_SLICE_X4Y139_AO5),
.O6(CLBLL_L_X4Y139_SLICE_X4Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55cc55ccaaccaacc)
  ) CLBLL_L_X4Y139_SLICE_X5Y139_DLUT (
.I0(CLBLM_R_X5Y127_SLICE_X7Y127_BQ),
.I1(CLBLL_L_X4Y138_SLICE_X5Y138_DO6),
.I2(1'b1),
.I3(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I4(1'b1),
.I5(CLBLL_L_X2Y152_SLICE_X0Y152_AQ),
.O5(CLBLL_L_X4Y139_SLICE_X5Y139_DO5),
.O6(CLBLL_L_X4Y139_SLICE_X5Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5acccc5a5acccc)
  ) CLBLL_L_X4Y139_SLICE_X5Y139_CLUT (
.I0(CLBLL_L_X2Y158_SLICE_X0Y158_AQ),
.I1(CLBLL_L_X4Y138_SLICE_X5Y138_CO6),
.I2(CLBLL_L_X4Y130_SLICE_X5Y130_AQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y139_SLICE_X5Y139_CO5),
.O6(CLBLL_L_X4Y139_SLICE_X5Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLL_L_X4Y139_SLICE_X5Y139_BLUT (
.I0(CLBLM_R_X5Y127_SLICE_X6Y127_CQ),
.I1(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO7),
.I2(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO0),
.I3(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO0),
.I4(BRAM_L_X6Y140_RAMB18_X0Y56_DO16),
.I5(BRAM_L_X6Y140_RAMB18_X0Y56_DO23),
.O5(CLBLL_L_X4Y139_SLICE_X5Y139_BO5),
.O6(CLBLL_L_X4Y139_SLICE_X5Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLL_L_X4Y139_SLICE_X5Y139_ALUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO0),
.I1(CLBLM_R_X5Y130_SLICE_X7Y130_BQ),
.I2(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO0),
.I3(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO7),
.I4(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO0),
.I5(BRAM_L_X6Y140_RAMB18_X0Y56_DO23),
.O5(CLBLL_L_X4Y139_SLICE_X5Y139_AO5),
.O6(CLBLL_L_X4Y139_SLICE_X5Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y140_SLICE_X4Y140_DO5),
.O6(CLBLL_L_X4Y140_SLICE_X4Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y140_SLICE_X4Y140_CO5),
.O6(CLBLL_L_X4Y140_SLICE_X4Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fcc0fccf0ccf0cc)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y139_SLICE_X4Y139_CO6),
.I2(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.I3(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y151_SLICE_X2Y151_BQ),
.O5(CLBLL_L_X4Y140_SLICE_X4Y140_BO5),
.O6(CLBLL_L_X4Y140_SLICE_X4Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33aaccaa33aaccaa)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_ALUT (
.I0(CLBLL_L_X4Y138_SLICE_X4Y138_DO6),
.I1(CLBLM_R_X3Y151_SLICE_X2Y151_DQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I4(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y140_SLICE_X4Y140_AO5),
.O6(CLBLL_L_X4Y140_SLICE_X4Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y140_SLICE_X5Y140_DO5),
.O6(CLBLL_L_X4Y140_SLICE_X5Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y140_SLICE_X5Y140_CO5),
.O6(CLBLL_L_X4Y140_SLICE_X5Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h30fc30fcfc30fc30)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I2(CLBLL_L_X4Y138_SLICE_X5Y138_AO6),
.I3(CLBLL_L_X4Y133_SLICE_X4Y133_BQ),
.I4(1'b1),
.I5(CLBLL_L_X2Y157_SLICE_X0Y157_BQ),
.O5(CLBLL_L_X4Y140_SLICE_X5Y140_BO5),
.O6(CLBLL_L_X4Y140_SLICE_X5Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff00ccff33cc00)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I2(1'b1),
.I3(CLBLM_R_X3Y149_SLICE_X3Y149_AQ),
.I4(CLBLL_L_X4Y139_SLICE_X5Y139_AO6),
.I5(CLBLM_R_X5Y130_SLICE_X7Y130_BQ),
.O5(CLBLL_L_X4Y140_SLICE_X5Y140_AO5),
.O6(CLBLL_L_X4Y140_SLICE_X5Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y165_IOB_X0Y166_I),
.Q(CLBLL_L_X4Y145_SLICE_X4Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y167_IOB_X0Y167_I),
.Q(CLBLL_L_X4Y145_SLICE_X4Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y145_SLICE_X4Y145_DO5),
.O6(CLBLL_L_X4Y145_SLICE_X4Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y145_SLICE_X4Y145_CO5),
.O6(CLBLL_L_X4Y145_SLICE_X4Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y145_SLICE_X4Y145_BO5),
.O6(CLBLL_L_X4Y145_SLICE_X4Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y145_SLICE_X4Y145_AO5),
.O6(CLBLL_L_X4Y145_SLICE_X4Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y145_SLICE_X5Y145_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y145_SLICE_X5Y145_DO5),
.O6(CLBLL_L_X4Y145_SLICE_X5Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y145_SLICE_X5Y145_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y145_SLICE_X5Y145_CO5),
.O6(CLBLL_L_X4Y145_SLICE_X5Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y145_SLICE_X5Y145_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y145_SLICE_X5Y145_BO5),
.O6(CLBLL_L_X4Y145_SLICE_X5Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y145_SLICE_X5Y145_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y145_SLICE_X5Y145_AO5),
.O6(CLBLL_L_X4Y145_SLICE_X5Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y169_IOB_X0Y169_I),
.Q(CLBLL_L_X4Y146_SLICE_X4Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y146_SLICE_X4Y146_DO5),
.O6(CLBLL_L_X4Y146_SLICE_X4Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y146_SLICE_X4Y146_CO5),
.O6(CLBLL_L_X4Y146_SLICE_X4Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y146_SLICE_X4Y146_BO5),
.O6(CLBLL_L_X4Y146_SLICE_X4Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y146_SLICE_X4Y146_AO5),
.O6(CLBLL_L_X4Y146_SLICE_X4Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y146_SLICE_X5Y146_DO5),
.O6(CLBLL_L_X4Y146_SLICE_X5Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y146_SLICE_X5Y146_CO5),
.O6(CLBLL_L_X4Y146_SLICE_X5Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y146_SLICE_X5Y146_BO5),
.O6(CLBLL_L_X4Y146_SLICE_X5Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y146_SLICE_X5Y146_AO5),
.O6(CLBLL_L_X4Y146_SLICE_X5Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y155_SLICE_X4Y155_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y193_IOB_X0Y194_I),
.Q(CLBLL_L_X4Y155_SLICE_X4Y155_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y155_SLICE_X4Y155_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y201_IOB_X0Y201_I),
.Q(CLBLL_L_X4Y155_SLICE_X4Y155_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y155_SLICE_X4Y155_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y231_IOB_X0Y232_I),
.Q(CLBLL_L_X4Y155_SLICE_X4Y155_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y155_SLICE_X4Y155_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y243_IOB_X0Y244_I),
.Q(CLBLL_L_X4Y155_SLICE_X4Y155_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y155_SLICE_X4Y155_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y155_SLICE_X4Y155_DO5),
.O6(CLBLL_L_X4Y155_SLICE_X4Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y155_SLICE_X4Y155_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y155_SLICE_X4Y155_CO5),
.O6(CLBLL_L_X4Y155_SLICE_X4Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y155_SLICE_X4Y155_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y155_SLICE_X4Y155_BO5),
.O6(CLBLL_L_X4Y155_SLICE_X4Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y155_SLICE_X4Y155_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y155_SLICE_X4Y155_AO5),
.O6(CLBLL_L_X4Y155_SLICE_X4Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y155_SLICE_X5Y155_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y155_SLICE_X5Y155_DO5),
.O6(CLBLL_L_X4Y155_SLICE_X5Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y155_SLICE_X5Y155_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y155_SLICE_X5Y155_CO5),
.O6(CLBLL_L_X4Y155_SLICE_X5Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y155_SLICE_X5Y155_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y155_SLICE_X5Y155_BO5),
.O6(CLBLL_L_X4Y155_SLICE_X5Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y155_SLICE_X5Y155_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y155_SLICE_X5Y155_AO5),
.O6(CLBLL_L_X4Y155_SLICE_X5Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y156_SLICE_X4Y156_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y207_IOB_X0Y207_I),
.Q(CLBLL_L_X4Y156_SLICE_X4Y156_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y156_SLICE_X4Y156_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y215_IOB_X0Y215_I),
.Q(CLBLL_L_X4Y156_SLICE_X4Y156_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y156_SLICE_X4Y156_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y215_IOB_X0Y216_I),
.Q(CLBLL_L_X4Y156_SLICE_X4Y156_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y156_SLICE_X4Y156_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y217_IOB_X0Y217_I),
.Q(CLBLL_L_X4Y156_SLICE_X4Y156_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y156_SLICE_X4Y156_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y156_SLICE_X4Y156_DO5),
.O6(CLBLL_L_X4Y156_SLICE_X4Y156_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y156_SLICE_X4Y156_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y156_SLICE_X4Y156_CO5),
.O6(CLBLL_L_X4Y156_SLICE_X4Y156_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y156_SLICE_X4Y156_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y156_SLICE_X4Y156_BO5),
.O6(CLBLL_L_X4Y156_SLICE_X4Y156_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y156_SLICE_X4Y156_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y156_SLICE_X4Y156_AO5),
.O6(CLBLL_L_X4Y156_SLICE_X4Y156_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y156_SLICE_X5Y156_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y247_IOB_X0Y247_I),
.Q(CLBLL_L_X4Y156_SLICE_X5Y156_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y156_SLICE_X5Y156_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(CLBLL_L_X4Y156_SLICE_X5Y156_AO6),
.Q(CLBLL_L_X4Y156_SLICE_X5Y156_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y156_SLICE_X5Y156_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y241_IOB_X0Y242_I),
.Q(CLBLL_L_X4Y156_SLICE_X5Y156_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y156_SLICE_X5Y156_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y245_IOB_X0Y245_I),
.Q(CLBLL_L_X4Y156_SLICE_X5Y156_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y156_SLICE_X5Y156_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y245_IOB_X0Y246_I),
.Q(CLBLL_L_X4Y156_SLICE_X5Y156_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y156_SLICE_X5Y156_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y156_SLICE_X5Y156_DO5),
.O6(CLBLL_L_X4Y156_SLICE_X5Y156_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y156_SLICE_X5Y156_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y156_SLICE_X5Y156_CO5),
.O6(CLBLL_L_X4Y156_SLICE_X5Y156_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y156_SLICE_X5Y156_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y156_SLICE_X5Y156_BO5),
.O6(CLBLL_L_X4Y156_SLICE_X5Y156_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLL_L_X4Y156_SLICE_X5Y156_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y237_IOB_X0Y237_I),
.O5(CLBLL_L_X4Y156_SLICE_X5Y156_AO5),
.O6(CLBLL_L_X4Y156_SLICE_X5Y156_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X54Y96_SLICE_X82Y96_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X0Y20_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X11Y130_AO5),
.Q(CLBLL_L_X54Y96_SLICE_X82Y96_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y96_SLICE_X82Y96_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y96_SLICE_X82Y96_DO5),
.O6(CLBLL_L_X54Y96_SLICE_X82Y96_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y96_SLICE_X82Y96_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y96_SLICE_X82Y96_CO5),
.O6(CLBLL_L_X54Y96_SLICE_X82Y96_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y96_SLICE_X82Y96_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y96_SLICE_X82Y96_BO5),
.O6(CLBLL_L_X54Y96_SLICE_X82Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y96_SLICE_X82Y96_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y96_SLICE_X82Y96_AO5),
.O6(CLBLL_L_X54Y96_SLICE_X82Y96_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y96_SLICE_X83Y96_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y96_SLICE_X83Y96_DO5),
.O6(CLBLL_L_X54Y96_SLICE_X83Y96_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y96_SLICE_X83Y96_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y96_SLICE_X83Y96_CO5),
.O6(CLBLL_L_X54Y96_SLICE_X83Y96_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y96_SLICE_X83Y96_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y96_SLICE_X83Y96_BO5),
.O6(CLBLL_L_X54Y96_SLICE_X83Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y96_SLICE_X83Y96_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y96_SLICE_X83Y96_AO5),
.O6(CLBLL_L_X54Y96_SLICE_X83Y96_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X54Y101_SLICE_X82Y101_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X8Y130_AO5),
.Q(CLBLL_L_X54Y101_SLICE_X82Y101_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y101_SLICE_X82Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y101_SLICE_X82Y101_DO5),
.O6(CLBLL_L_X54Y101_SLICE_X82Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y101_SLICE_X82Y101_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y101_SLICE_X82Y101_CO5),
.O6(CLBLL_L_X54Y101_SLICE_X82Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y101_SLICE_X82Y101_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y101_SLICE_X82Y101_BO5),
.O6(CLBLL_L_X54Y101_SLICE_X82Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y101_SLICE_X82Y101_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y101_SLICE_X82Y101_AO5),
.O6(CLBLL_L_X54Y101_SLICE_X82Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y101_SLICE_X83Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y101_SLICE_X83Y101_DO5),
.O6(CLBLL_L_X54Y101_SLICE_X83Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y101_SLICE_X83Y101_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y101_SLICE_X83Y101_CO5),
.O6(CLBLL_L_X54Y101_SLICE_X83Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y101_SLICE_X83Y101_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y101_SLICE_X83Y101_BO5),
.O6(CLBLL_L_X54Y101_SLICE_X83Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y101_SLICE_X83Y101_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y101_SLICE_X83Y101_AO5),
.O6(CLBLL_L_X54Y101_SLICE_X83Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X54Y105_SLICE_X82Y105_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y133_SLICE_X11Y133_AO5),
.Q(CLBLL_L_X54Y105_SLICE_X82Y105_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y105_SLICE_X82Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y105_SLICE_X82Y105_DO5),
.O6(CLBLL_L_X54Y105_SLICE_X82Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y105_SLICE_X82Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y105_SLICE_X82Y105_CO5),
.O6(CLBLL_L_X54Y105_SLICE_X82Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y105_SLICE_X82Y105_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y105_SLICE_X82Y105_BO5),
.O6(CLBLL_L_X54Y105_SLICE_X82Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y105_SLICE_X82Y105_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y105_SLICE_X82Y105_AO5),
.O6(CLBLL_L_X54Y105_SLICE_X82Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y105_SLICE_X83Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y105_SLICE_X83Y105_DO5),
.O6(CLBLL_L_X54Y105_SLICE_X83Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y105_SLICE_X83Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y105_SLICE_X83Y105_CO5),
.O6(CLBLL_L_X54Y105_SLICE_X83Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y105_SLICE_X83Y105_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y105_SLICE_X83Y105_BO5),
.O6(CLBLL_L_X54Y105_SLICE_X83Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y105_SLICE_X83Y105_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y105_SLICE_X83Y105_AO5),
.O6(CLBLL_L_X54Y105_SLICE_X83Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X54Y116_SLICE_X82Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y135_SLICE_X5Y135_AO5),
.Q(CLBLL_L_X54Y116_SLICE_X82Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y116_SLICE_X82Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y116_SLICE_X82Y116_DO5),
.O6(CLBLL_L_X54Y116_SLICE_X82Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y116_SLICE_X82Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y116_SLICE_X82Y116_CO5),
.O6(CLBLL_L_X54Y116_SLICE_X82Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y116_SLICE_X82Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y116_SLICE_X82Y116_BO5),
.O6(CLBLL_L_X54Y116_SLICE_X82Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y116_SLICE_X82Y116_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y116_SLICE_X82Y116_AO5),
.O6(CLBLL_L_X54Y116_SLICE_X82Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y116_SLICE_X83Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y116_SLICE_X83Y116_DO5),
.O6(CLBLL_L_X54Y116_SLICE_X83Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y116_SLICE_X83Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y116_SLICE_X83Y116_CO5),
.O6(CLBLL_L_X54Y116_SLICE_X83Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y116_SLICE_X83Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y116_SLICE_X83Y116_BO5),
.O6(CLBLL_L_X54Y116_SLICE_X83Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y116_SLICE_X83Y116_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y116_SLICE_X83Y116_AO5),
.O6(CLBLL_L_X54Y116_SLICE_X83Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X54Y119_SLICE_X82Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X6Y134_BO5),
.Q(CLBLL_L_X54Y119_SLICE_X82Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y119_SLICE_X82Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y119_SLICE_X82Y119_DO5),
.O6(CLBLL_L_X54Y119_SLICE_X82Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y119_SLICE_X82Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y119_SLICE_X82Y119_CO5),
.O6(CLBLL_L_X54Y119_SLICE_X82Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y119_SLICE_X82Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y119_SLICE_X82Y119_BO5),
.O6(CLBLL_L_X54Y119_SLICE_X82Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y119_SLICE_X82Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y119_SLICE_X82Y119_AO5),
.O6(CLBLL_L_X54Y119_SLICE_X82Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y119_SLICE_X83Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y119_SLICE_X83Y119_DO5),
.O6(CLBLL_L_X54Y119_SLICE_X83Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y119_SLICE_X83Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y119_SLICE_X83Y119_CO5),
.O6(CLBLL_L_X54Y119_SLICE_X83Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y119_SLICE_X83Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y119_SLICE_X83Y119_BO5),
.O6(CLBLL_L_X54Y119_SLICE_X83Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y119_SLICE_X83Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y119_SLICE_X83Y119_AO5),
.O6(CLBLL_L_X54Y119_SLICE_X83Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X54Y123_SLICE_X82Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X6Y134_AO5),
.Q(CLBLL_L_X54Y123_SLICE_X82Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y123_SLICE_X82Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y123_SLICE_X82Y123_DO5),
.O6(CLBLL_L_X54Y123_SLICE_X82Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y123_SLICE_X82Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y123_SLICE_X82Y123_CO5),
.O6(CLBLL_L_X54Y123_SLICE_X82Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y123_SLICE_X82Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y123_SLICE_X82Y123_BO5),
.O6(CLBLL_L_X54Y123_SLICE_X82Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y123_SLICE_X82Y123_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y123_SLICE_X82Y123_AO5),
.O6(CLBLL_L_X54Y123_SLICE_X82Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y123_SLICE_X83Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y123_SLICE_X83Y123_DO5),
.O6(CLBLL_L_X54Y123_SLICE_X83Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y123_SLICE_X83Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y123_SLICE_X83Y123_CO5),
.O6(CLBLL_L_X54Y123_SLICE_X83Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y123_SLICE_X83Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y123_SLICE_X83Y123_BO5),
.O6(CLBLL_L_X54Y123_SLICE_X83Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y123_SLICE_X83Y123_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y123_SLICE_X83Y123_AO5),
.O6(CLBLL_L_X54Y123_SLICE_X83Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X54Y133_SLICE_X82Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y135_SLICE_X4Y135_AO5),
.Q(CLBLL_L_X54Y133_SLICE_X82Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y133_SLICE_X82Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y133_SLICE_X82Y133_DO5),
.O6(CLBLL_L_X54Y133_SLICE_X82Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y133_SLICE_X82Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y133_SLICE_X82Y133_CO5),
.O6(CLBLL_L_X54Y133_SLICE_X82Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y133_SLICE_X82Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y133_SLICE_X82Y133_BO5),
.O6(CLBLL_L_X54Y133_SLICE_X82Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y133_SLICE_X82Y133_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y133_SLICE_X82Y133_AO5),
.O6(CLBLL_L_X54Y133_SLICE_X82Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y133_SLICE_X83Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y133_SLICE_X83Y133_DO5),
.O6(CLBLL_L_X54Y133_SLICE_X83Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y133_SLICE_X83Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y133_SLICE_X83Y133_CO5),
.O6(CLBLL_L_X54Y133_SLICE_X83Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y133_SLICE_X83Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y133_SLICE_X83Y133_BO5),
.O6(CLBLL_L_X54Y133_SLICE_X83Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y133_SLICE_X83Y133_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y133_SLICE_X83Y133_AO5),
.O6(CLBLL_L_X54Y133_SLICE_X83Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X54Y138_SLICE_X82Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y137_SLICE_X5Y137_AO5),
.Q(CLBLL_L_X54Y138_SLICE_X82Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y138_SLICE_X82Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y138_SLICE_X82Y138_DO5),
.O6(CLBLL_L_X54Y138_SLICE_X82Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y138_SLICE_X82Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y138_SLICE_X82Y138_CO5),
.O6(CLBLL_L_X54Y138_SLICE_X82Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y138_SLICE_X82Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y138_SLICE_X82Y138_BO5),
.O6(CLBLL_L_X54Y138_SLICE_X82Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y138_SLICE_X82Y138_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y138_SLICE_X82Y138_AO5),
.O6(CLBLL_L_X54Y138_SLICE_X82Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y138_SLICE_X83Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y138_SLICE_X83Y138_DO5),
.O6(CLBLL_L_X54Y138_SLICE_X83Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y138_SLICE_X83Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y138_SLICE_X83Y138_CO5),
.O6(CLBLL_L_X54Y138_SLICE_X83Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y138_SLICE_X83Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y138_SLICE_X83Y138_BO5),
.O6(CLBLL_L_X54Y138_SLICE_X83Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y138_SLICE_X83Y138_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y138_SLICE_X83Y138_AO5),
.O6(CLBLL_L_X54Y138_SLICE_X83Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X54Y141_SLICE_X82Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y137_SLICE_X3Y137_AO5),
.Q(CLBLL_L_X54Y141_SLICE_X82Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y141_SLICE_X82Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y141_SLICE_X82Y141_DO5),
.O6(CLBLL_L_X54Y141_SLICE_X82Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y141_SLICE_X82Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y141_SLICE_X82Y141_CO5),
.O6(CLBLL_L_X54Y141_SLICE_X82Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y141_SLICE_X82Y141_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y141_SLICE_X82Y141_BO5),
.O6(CLBLL_L_X54Y141_SLICE_X82Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y141_SLICE_X82Y141_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y141_SLICE_X82Y141_AO5),
.O6(CLBLL_L_X54Y141_SLICE_X82Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y141_SLICE_X83Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y141_SLICE_X83Y141_DO5),
.O6(CLBLL_L_X54Y141_SLICE_X83Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y141_SLICE_X83Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y141_SLICE_X83Y141_CO5),
.O6(CLBLL_L_X54Y141_SLICE_X83Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y141_SLICE_X83Y141_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y141_SLICE_X83Y141_BO5),
.O6(CLBLL_L_X54Y141_SLICE_X83Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y141_SLICE_X83Y141_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y141_SLICE_X83Y141_AO5),
.O6(CLBLL_L_X54Y141_SLICE_X83Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y127_SLICE_X10Y127_AO6),
.Q(CLBLM_L_X8Y127_SLICE_X10Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y127_SLICE_X10Y127_BO6),
.Q(CLBLM_L_X8Y127_SLICE_X10Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y127_SLICE_X10Y127_DO5),
.O6(CLBLM_L_X8Y127_SLICE_X10Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y127_SLICE_X10Y127_CO5),
.O6(CLBLM_L_X8Y127_SLICE_X10Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3c3c3c3c3c)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_BLUT (
.I0(1'b1),
.I1(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO3),
.I2(CLBLM_R_X5Y126_SLICE_X6Y126_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y127_SLICE_X10Y127_BO5),
.O6(CLBLM_L_X8Y127_SLICE_X10Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0ff0f0f0f0)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X5Y125_SLICE_X7Y125_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO1),
.O5(CLBLM_L_X8Y127_SLICE_X10Y127_AO5),
.O6(CLBLM_L_X8Y127_SLICE_X10Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y127_SLICE_X11Y127_DO5),
.O6(CLBLM_L_X8Y127_SLICE_X11Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y127_SLICE_X11Y127_CO5),
.O6(CLBLM_L_X8Y127_SLICE_X11Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y127_SLICE_X11Y127_BO5),
.O6(CLBLM_L_X8Y127_SLICE_X11Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y127_SLICE_X11Y127_AO5),
.O6(CLBLM_L_X8Y127_SLICE_X11Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y129_SLICE_X10Y129_AO6),
.Q(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y129_SLICE_X10Y129_BO6),
.Q(CLBLM_L_X8Y129_SLICE_X10Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y129_SLICE_X10Y129_CO6),
.Q(CLBLM_L_X8Y129_SLICE_X10Y129_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y129_SLICE_X10Y129_DO5),
.O6(CLBLM_L_X8Y129_SLICE_X10Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ffff00ff00)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO6),
.I4(1'b1),
.I5(CLBLM_R_X5Y127_SLICE_X6Y127_B5Q),
.O5(CLBLM_L_X8Y129_SLICE_X10Y129_CO5),
.O6(CLBLM_L_X8Y129_SLICE_X10Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3c3c3c3c3c)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_BLUT (
.I0(1'b1),
.I1(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO5),
.I2(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y129_SLICE_X10Y129_BO5),
.O6(CLBLM_L_X8Y129_SLICE_X10Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5a5a5a5a5a)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_ALUT (
.I0(CLBLM_R_X5Y126_SLICE_X7Y126_AQ),
.I1(1'b1),
.I2(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO4),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y129_SLICE_X10Y129_AO5),
.O6(CLBLM_L_X8Y129_SLICE_X10Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y129_SLICE_X11Y129_DO5),
.O6(CLBLM_L_X8Y129_SLICE_X11Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y129_SLICE_X11Y129_CO5),
.O6(CLBLM_L_X8Y129_SLICE_X11Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y129_SLICE_X11Y129_BO5),
.O6(CLBLM_L_X8Y129_SLICE_X11Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y129_SLICE_X11Y129_AO5),
.O6(CLBLM_L_X8Y129_SLICE_X11Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X10Y130_AO5),
.Q(CLBLM_L_X8Y130_SLICE_X10Y130_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X10Y130_BO5),
.Q(CLBLM_L_X8Y130_SLICE_X10Y130_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X10Y130_AO6),
.Q(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X10Y130_BO6),
.Q(CLBLM_L_X8Y130_SLICE_X10Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X10Y130_CO6),
.Q(CLBLM_L_X8Y130_SLICE_X10Y130_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X10Y130_DO6),
.Q(CLBLM_L_X8Y130_SLICE_X10Y130_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5a5a5a5a5a)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_DLUT (
.I0(CLBLM_R_X5Y128_SLICE_X6Y128_AQ),
.I1(1'b1),
.I2(BRAM_L_X6Y135_RAMB18_X0Y54_DO19),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y130_SLICE_X10Y130_DO5),
.O6(CLBLM_L_X8Y130_SLICE_X10Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa55aa55aa55aa)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_CLUT (
.I0(CLBLL_L_X4Y130_SLICE_X5Y130_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(BRAM_L_X6Y140_RAMB18_X0Y56_DO2),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y130_SLICE_X10Y130_CO5),
.O6(CLBLM_L_X8Y130_SLICE_X10Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa55aaf0f06666)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_BLUT (
.I0(CLBLM_L_X8Y130_SLICE_X10Y130_B5Q),
.I1(BRAM_L_X6Y125_RAMB18_X0Y50_DO19),
.I2(LIOB33_X0Y125_IOB_X0Y126_I),
.I3(BRAM_L_X6Y135_RAMB18_X0Y54_DO3),
.I4(LIOB33_X0Y147_IOB_X0Y148_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y130_SLICE_X10Y130_BO5),
.O6(CLBLM_L_X8Y130_SLICE_X10Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h66666666ff3c003c)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_ALUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO7),
.I1(CLBLM_L_X8Y130_SLICE_X10Y130_A5Q),
.I2(BRAM_L_X6Y125_RAMB18_X0Y50_DO7),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(LIOB33_X0Y121_IOB_X0Y122_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y130_SLICE_X10Y130_AO5),
.O6(CLBLM_L_X8Y130_SLICE_X10Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X11Y130_BO6),
.Q(CLBLM_L_X8Y130_SLICE_X11Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X11Y130_CO6),
.Q(CLBLM_L_X8Y130_SLICE_X11Y130_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X11Y130_DO6),
.Q(CLBLM_L_X8Y130_SLICE_X11Y130_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555555aaaaaaaa)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_DLUT (
.I0(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO2),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X4Y131_SLICE_X4Y131_BQ),
.O5(CLBLM_L_X8Y130_SLICE_X11Y130_DO5),
.O6(CLBLM_L_X8Y130_SLICE_X11Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333333cccccccc)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_CLUT (
.I0(1'b1),
.I1(BRAM_L_X6Y135_RAMB18_X0Y54_DO21),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X3Y130_SLICE_X3Y130_AQ),
.O5(CLBLM_L_X8Y130_SLICE_X11Y130_CO5),
.O6(CLBLM_L_X8Y130_SLICE_X11Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333cccc3333cccc)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_BLUT (
.I0(1'b1),
.I1(BRAM_L_X6Y135_RAMB18_X0Y54_DO17),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X4Y129_SLICE_X4Y129_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y130_SLICE_X11Y130_BO5),
.O6(CLBLM_L_X8Y130_SLICE_X11Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa55aa5a5a5a5a)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_ALUT (
.I0(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO0),
.I1(1'b1),
.I2(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.I3(BRAM_R_X17Y135_RAMB18_X1Y54_DO16),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y130_SLICE_X11Y130_AO5),
.O6(CLBLM_L_X8Y130_SLICE_X11Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X10Y131_AO6),
.Q(CLBLM_L_X8Y131_SLICE_X10Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X10Y131_BO6),
.Q(CLBLM_L_X8Y131_SLICE_X10Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_DLUT (
.I0(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO1),
.I1(BRAM_R_X17Y135_RAMB18_X1Y54_DO17),
.I2(CLBLM_R_X5Y125_SLICE_X7Y125_AQ),
.I3(BRAM_L_X6Y135_RAMB18_X0Y54_DO17),
.I4(BRAM_R_X17Y135_RAMB18_X1Y54_DO16),
.I5(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO0),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_DO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_CLUT (
.I0(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO2),
.I1(BRAM_R_X17Y135_RAMB18_X1Y54_DO19),
.I2(CLBLM_R_X5Y126_SLICE_X6Y126_AQ),
.I3(BRAM_R_X17Y135_RAMB18_X1Y54_DO18),
.I4(BRAM_L_X6Y135_RAMB18_X0Y54_DO19),
.I5(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO3),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_CO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555555aaaaaaaa)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_BLUT (
.I0(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO3),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y133_SLICE_X6Y133_AQ),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_BO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ffff00ff00)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO5),
.I4(1'b1),
.I5(CLBLL_L_X4Y132_SLICE_X5Y132_AQ),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_AO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X11Y131_AO6),
.Q(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X11Y131_BO6),
.Q(CLBLM_L_X8Y131_SLICE_X11Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X11Y131_CO6),
.Q(CLBLM_L_X8Y131_SLICE_X11Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_DLUT (
.I0(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO0),
.I1(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO0),
.I2(BRAM_R_X17Y135_RAMB18_X1Y54_DO23),
.I3(CLBLM_R_X3Y131_SLICE_X3Y131_BQ),
.I4(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO7),
.I5(BRAM_L_X6Y135_RAMB18_X0Y54_DO16),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_DO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa55aa55aa55aa)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_CLUT (
.I0(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_L_X4Y131_SLICE_X4Y131_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_CO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333333cccccccc)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y131_SLICE_X7Y131_A5Q),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO0),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_BO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555555aaaaaaaa)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_ALUT (
.I0(CLBLL_L_X4Y131_SLICE_X5Y131_B5Q),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(BRAM_L_X6Y135_RAMB18_X0Y54_DO22),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_AO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_DLUT (
.I0(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO1),
.I1(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO1),
.I2(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO0),
.I3(CLBLL_L_X4Y131_SLICE_X4Y131_CQ),
.I4(BRAM_L_X6Y135_RAMB18_X0Y54_DO17),
.I5(BRAM_R_X17Y135_RAMB18_X1Y54_DO16),
.O5(CLBLM_L_X8Y132_SLICE_X10Y132_DO5),
.O6(CLBLM_L_X8Y132_SLICE_X10Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_CLUT (
.I0(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO2),
.I1(BRAM_R_X17Y135_RAMB18_X1Y54_DO18),
.I2(BRAM_L_X6Y135_RAMB18_X0Y54_DO19),
.I3(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO3),
.I4(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO3),
.I5(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.O5(CLBLM_L_X8Y132_SLICE_X10Y132_CO5),
.O6(CLBLM_L_X8Y132_SLICE_X10Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffff0096969696)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_BLUT (
.I0(CLBLM_L_X8Y132_SLICE_X10Y132_DO6),
.I1(BRAM_R_X17Y135_RAMB18_X1Y54_DO23),
.I2(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO7),
.I3(CLBLM_R_X5Y158_SLICE_X6Y158_CQ),
.I4(CLBLL_L_X4Y131_SLICE_X4Y131_CQ),
.I5(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.O5(CLBLM_L_X8Y132_SLICE_X10Y132_BO5),
.O6(CLBLM_L_X8Y132_SLICE_X10Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3a35cac5353ac5ca)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_ALUT (
.I0(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO7),
.I1(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I3(BRAM_R_X17Y135_RAMB18_X1Y54_DO23),
.I4(CLBLM_R_X5Y158_SLICE_X6Y158_DQ),
.I5(CLBLM_L_X8Y132_SLICE_X10Y132_CO6),
.O5(CLBLM_L_X8Y132_SLICE_X10Y132_AO5),
.O6(CLBLM_L_X8Y132_SLICE_X10Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y132_SLICE_X11Y132_AO5),
.Q(CLBLM_L_X8Y132_SLICE_X11Y132_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y132_SLICE_X11Y132_AO6),
.Q(CLBLM_L_X8Y132_SLICE_X11Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y132_SLICE_X11Y132_BO6),
.Q(CLBLM_L_X8Y132_SLICE_X11Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y132_SLICE_X11Y132_CO6),
.Q(CLBLM_L_X8Y132_SLICE_X11Y132_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_DLUT (
.I0(CLBLL_L_X4Y131_SLICE_X4Y131_AQ),
.I1(BRAM_R_X17Y135_RAMB18_X1Y54_DO17),
.I2(BRAM_L_X6Y135_RAMB18_X0Y54_DO17),
.I3(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO1),
.I4(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO0),
.I5(BRAM_L_X6Y135_RAMB18_X0Y54_DO16),
.O5(CLBLM_L_X8Y132_SLICE_X11Y132_DO5),
.O6(CLBLM_L_X8Y132_SLICE_X11Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0ff0f0f0f0)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO6),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X4Y132_SLICE_X4Y132_BQ),
.O5(CLBLM_L_X8Y132_SLICE_X11Y132_CO5),
.O6(CLBLM_L_X8Y132_SLICE_X11Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555555aaaaaaaa)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_BLUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y56_DO22),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y132_SLICE_X7Y132_B5Q),
.O5(CLBLM_L_X8Y132_SLICE_X11Y132_BO5),
.O6(CLBLM_L_X8Y132_SLICE_X11Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffff00b1b1e4e4)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_ALUT (
.I0(LIOB33_X0Y147_IOB_X0Y148_I),
.I1(BRAM_L_X6Y130_RAMB18_X0Y52_DO0),
.I2(LIOB33_X0Y131_IOB_X0Y132_I),
.I3(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO0),
.I4(CLBLM_L_X8Y132_SLICE_X11Y132_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y132_SLICE_X11Y132_AO5),
.O6(CLBLM_L_X8Y132_SLICE_X11Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_DLUT (
.I0(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO2),
.I1(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO3),
.I2(BRAM_R_X17Y135_RAMB18_X1Y54_DO19),
.I3(BRAM_L_X6Y135_RAMB18_X0Y54_DO18),
.I4(BRAM_L_X6Y135_RAMB18_X0Y54_DO19),
.I5(CLBLM_R_X5Y133_SLICE_X6Y133_AQ),
.O5(CLBLM_L_X8Y133_SLICE_X10Y133_DO5),
.O6(CLBLM_L_X8Y133_SLICE_X10Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_CLUT (
.I0(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.I1(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO4),
.I2(BRAM_L_X6Y135_RAMB18_X0Y54_DO19),
.I3(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO3),
.I4(BRAM_R_X17Y135_RAMB18_X1Y54_DO20),
.I5(BRAM_L_X6Y135_RAMB18_X0Y54_DO20),
.O5(CLBLM_L_X8Y133_SLICE_X10Y133_CO5),
.O6(CLBLM_L_X8Y133_SLICE_X10Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h72d8278d278d72d8)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_BLUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I1(CLBLM_R_X5Y158_SLICE_X6Y158_BQ),
.I2(CLBLM_L_X8Y133_SLICE_X10Y133_DO6),
.I3(CLBLM_R_X5Y133_SLICE_X6Y133_AQ),
.I4(BRAM_L_X6Y135_RAMB18_X0Y54_DO23),
.I5(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO7),
.O5(CLBLM_L_X8Y133_SLICE_X10Y133_BO5),
.O6(CLBLM_L_X8Y133_SLICE_X10Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7227d88d27728dd8)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_ALUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I1(CLBLM_R_X3Y158_SLICE_X2Y158_BQ),
.I2(BRAM_L_X6Y135_RAMB18_X0Y54_DO23),
.I3(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO7),
.I4(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.I5(CLBLM_L_X8Y133_SLICE_X10Y133_CO6),
.O5(CLBLM_L_X8Y133_SLICE_X10Y133_AO5),
.O6(CLBLM_L_X8Y133_SLICE_X10Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5050afafa0a0)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_DLUT (
.I0(CLBLM_R_X3Y158_SLICE_X2Y158_DQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y131_SLICE_X11Y131_DO6),
.I5(CLBLM_R_X3Y131_SLICE_X3Y131_BQ),
.O5(CLBLM_L_X8Y133_SLICE_X11Y133_DO5),
.O6(CLBLM_L_X8Y133_SLICE_X11Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff066990ff09966)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_CLUT (
.I0(CLBLM_L_X8Y133_SLICE_X11Y133_AO6),
.I1(BRAM_L_X6Y135_RAMB18_X0Y54_DO16),
.I2(CLBLM_R_X5Y158_SLICE_X6Y158_AQ),
.I3(CLBLM_R_X5Y131_SLICE_X7Y131_A5Q),
.I4(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I5(CLBLM_L_X8Y130_SLICE_X11Y130_AO6),
.O5(CLBLM_L_X8Y133_SLICE_X11Y133_CO5),
.O6(CLBLM_L_X8Y133_SLICE_X11Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_BLUT (
.I0(BRAM_R_X17Y135_RAMB18_X1Y54_DO19),
.I1(BRAM_L_X6Y135_RAMB18_X0Y54_DO20),
.I2(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO4),
.I3(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO3),
.I4(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO4),
.I5(CLBLM_R_X3Y131_SLICE_X3Y131_DQ),
.O5(CLBLM_L_X8Y133_SLICE_X11Y133_BO5),
.O6(CLBLM_L_X8Y133_SLICE_X11Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333cccc0f0ff0f0)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_ALUT (
.I0(1'b1),
.I1(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO7),
.I2(CLBLM_R_X3Y134_SLICE_X2Y134_AQ),
.I3(1'b1),
.I4(BRAM_L_X6Y135_RAMB18_X0Y54_DO23),
.I5(1'b1),
.O5(CLBLM_L_X8Y133_SLICE_X11Y133_AO5),
.O6(CLBLM_L_X8Y133_SLICE_X11Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y134_SLICE_X10Y134_AO6),
.Q(CLBLM_L_X8Y134_SLICE_X10Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_DLUT (
.I0(CLBLM_R_X7Y125_SLICE_X8Y125_C5Q),
.I1(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO2),
.I2(BRAM_R_X17Y135_RAMB18_X1Y54_DO1),
.I3(BRAM_L_X6Y135_RAMB18_X0Y54_DO2),
.I4(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO1),
.I5(BRAM_R_X17Y135_RAMB18_X1Y54_DO2),
.O5(CLBLM_L_X8Y134_SLICE_X10Y134_DO5),
.O6(CLBLM_L_X8Y134_SLICE_X10Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_CLUT (
.I0(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO1),
.I1(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO2),
.I2(BRAM_L_X6Y135_RAMB18_X0Y54_DO17),
.I3(BRAM_R_X17Y135_RAMB18_X1Y54_DO18),
.I4(BRAM_L_X6Y135_RAMB18_X0Y54_DO18),
.I5(CLBLL_L_X4Y131_SLICE_X4Y131_BQ),
.O5(CLBLM_L_X8Y134_SLICE_X10Y134_CO5),
.O6(CLBLM_L_X8Y134_SLICE_X10Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_BLUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y54_DO18),
.I1(BRAM_R_X17Y135_RAMB18_X1Y54_DO17),
.I2(CLBLM_R_X3Y131_SLICE_X3Y131_CQ),
.I3(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO2),
.I4(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO1),
.I5(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO2),
.O5(CLBLM_L_X8Y134_SLICE_X10Y134_BO5),
.O6(CLBLM_L_X8Y134_SLICE_X10Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cc33cc33cc33cc)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_ALUT (
.I0(1'b1),
.I1(BRAM_L_X6Y140_RAMB18_X0Y56_DO20),
.I2(1'b1),
.I3(CLBLM_R_X5Y133_SLICE_X6Y133_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y134_SLICE_X10Y134_AO5),
.O6(CLBLM_L_X8Y134_SLICE_X10Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33aa33aaccaaccaa)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_DLUT (
.I0(CLBLM_L_X8Y134_SLICE_X11Y134_AO6),
.I1(CLBLM_R_X3Y132_SLICE_X3Y132_BQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y157_SLICE_X2Y157_BQ),
.O5(CLBLM_L_X8Y134_SLICE_X11Y134_DO5),
.O6(CLBLM_L_X8Y134_SLICE_X11Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_CLUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y54_DO21),
.I1(CLBLM_R_X5Y132_SLICE_X6Y132_AQ),
.I2(BRAM_L_X6Y135_RAMB18_X0Y54_DO20),
.I3(BRAM_R_X17Y135_RAMB18_X1Y54_DO21),
.I4(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO4),
.I5(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO5),
.O5(CLBLM_L_X8Y134_SLICE_X11Y134_CO5),
.O6(CLBLM_L_X8Y134_SLICE_X11Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff00ff099996666)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_BLUT (
.I0(CLBLM_L_X8Y132_SLICE_X11Y132_DO6),
.I1(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO7),
.I2(CLBLL_L_X4Y131_SLICE_X4Y131_AQ),
.I3(CLBLM_R_X3Y155_SLICE_X2Y155_CQ),
.I4(BRAM_L_X6Y135_RAMB18_X0Y54_DO23),
.I5(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.O5(CLBLM_L_X8Y134_SLICE_X11Y134_BO5),
.O6(CLBLM_L_X8Y134_SLICE_X11Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_ALUT (
.I0(BRAM_R_X17Y135_RAMB18_X1Y54_DO20),
.I1(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO5),
.I2(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO5),
.I3(BRAM_L_X6Y135_RAMB18_X0Y54_DO21),
.I4(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO4),
.I5(CLBLM_R_X3Y132_SLICE_X3Y132_BQ),
.O5(CLBLM_L_X8Y134_SLICE_X11Y134_AO5),
.O6(CLBLM_L_X8Y134_SLICE_X11Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y135_SLICE_X10Y135_AO5),
.Q(CLBLM_L_X8Y135_SLICE_X10Y135_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y135_SLICE_X10Y135_AO6),
.Q(CLBLM_L_X8Y135_SLICE_X10Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55cc55ccaaccaacc)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_DLUT (
.I0(CLBLL_L_X4Y155_SLICE_X4Y155_CQ),
.I1(CLBLM_L_X8Y134_SLICE_X10Y134_CO6),
.I2(1'b1),
.I3(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y131_SLICE_X4Y131_BQ),
.O5(CLBLM_L_X8Y135_SLICE_X10Y135_DO5),
.O6(CLBLM_L_X8Y135_SLICE_X10Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff3300ccffcc00)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y158_SLICE_X2Y158_CQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I4(CLBLM_L_X8Y135_SLICE_X10Y135_BO6),
.I5(CLBLL_L_X4Y132_SLICE_X4Y132_BQ),
.O5(CLBLM_L_X8Y135_SLICE_X10Y135_CO5),
.O6(CLBLM_L_X8Y135_SLICE_X10Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_BLUT (
.I0(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO5),
.I1(CLBLL_L_X4Y132_SLICE_X4Y132_BQ),
.I2(BRAM_R_X17Y135_RAMB18_X1Y54_DO22),
.I3(BRAM_L_X6Y135_RAMB18_X0Y54_DO21),
.I4(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO6),
.I5(BRAM_L_X6Y135_RAMB18_X0Y54_DO22),
.O5(CLBLM_L_X8Y135_SLICE_X10Y135_BO5),
.O6(CLBLM_L_X8Y135_SLICE_X10Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h66666666f033f0cc)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_ALUT (
.I0(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO1),
.I1(CLBLM_L_X8Y135_SLICE_X10Y135_A5Q),
.I2(LIOB33_X0Y133_IOB_X0Y133_I),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(BRAM_L_X6Y130_RAMB18_X0Y52_DO1),
.I5(1'b1),
.O5(CLBLM_L_X8Y135_SLICE_X10Y135_AO5),
.O6(CLBLM_L_X8Y135_SLICE_X10Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7b7b7b7b48484848)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_DLUT (
.I0(CLBLM_R_X5Y132_SLICE_X6Y132_AQ),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I2(CLBLL_L_X2Y158_SLICE_X0Y158_DQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X8Y134_SLICE_X11Y134_CO6),
.O5(CLBLM_L_X8Y135_SLICE_X11Y135_DO5),
.O6(CLBLM_L_X8Y135_SLICE_X11Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h77bb77bb44884488)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_CLUT (
.I0(CLBLL_L_X4Y155_SLICE_X4Y155_DQ),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I2(1'b1),
.I3(CLBLM_R_X3Y132_SLICE_X2Y132_CQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y135_SLICE_X11Y135_BO6),
.O5(CLBLM_L_X8Y135_SLICE_X11Y135_CO5),
.O6(CLBLM_L_X8Y135_SLICE_X11Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_BLUT (
.I0(BRAM_R_X17Y135_RAMB18_X1Y54_DO21),
.I1(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO6),
.I2(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO6),
.I3(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO5),
.I4(CLBLM_R_X3Y132_SLICE_X2Y132_CQ),
.I5(BRAM_L_X6Y135_RAMB18_X0Y54_DO22),
.O5(CLBLM_L_X8Y135_SLICE_X11Y135_BO5),
.O6(CLBLM_L_X8Y135_SLICE_X11Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7447b88b47748bb8)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_ALUT (
.I0(CLBLM_R_X3Y131_SLICE_X3Y131_DQ),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I2(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO7),
.I3(CLBLM_L_X8Y133_SLICE_X11Y133_BO6),
.I4(CLBLL_L_X4Y156_SLICE_X5Y156_BQ),
.I5(BRAM_R_X17Y135_RAMB18_X1Y54_DO23),
.O5(CLBLM_L_X8Y135_SLICE_X11Y135_AO5),
.O6(CLBLM_L_X8Y135_SLICE_X11Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y136_SLICE_X10Y136_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y136_SLICE_X10Y136_AO5),
.Q(CLBLM_L_X8Y136_SLICE_X10Y136_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y136_SLICE_X10Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y136_SLICE_X10Y136_AO6),
.Q(CLBLM_L_X8Y136_SLICE_X10Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X8Y136_SLICE_X10Y136_DLUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y54_DO1),
.I1(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO1),
.I2(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO0),
.I3(BRAM_R_X17Y135_RAMB18_X1Y54_DO0),
.I4(CLBLM_R_X7Y125_SLICE_X8Y125_B5Q),
.I5(BRAM_R_X17Y135_RAMB18_X1Y54_DO1),
.O5(CLBLM_L_X8Y136_SLICE_X10Y136_DO5),
.O6(CLBLM_L_X8Y136_SLICE_X10Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55c3553caac3aa3c)
  ) CLBLM_L_X8Y136_SLICE_X10Y136_CLUT (
.I0(CLBLM_L_X8Y130_SLICE_X10Y130_B5Q),
.I1(BRAM_L_X6Y135_RAMB18_X0Y54_DO7),
.I2(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO7),
.I3(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I4(CLBLM_L_X8Y136_SLICE_X10Y136_BO6),
.I5(CLBLM_L_X16Y151_SLICE_X22Y151_AQ),
.O5(CLBLM_L_X8Y136_SLICE_X10Y136_CO5),
.O6(CLBLM_L_X8Y136_SLICE_X10Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X8Y136_SLICE_X10Y136_BLUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO2),
.I1(BRAM_L_X6Y135_RAMB18_X0Y54_DO2),
.I2(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO3),
.I3(BRAM_R_X17Y135_RAMB18_X1Y54_DO3),
.I4(CLBLM_L_X8Y130_SLICE_X10Y130_B5Q),
.I5(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO3),
.O5(CLBLM_L_X8Y136_SLICE_X10Y136_BO5),
.O6(CLBLM_L_X8Y136_SLICE_X10Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5aff006666)
  ) CLBLM_L_X8Y136_SLICE_X10Y136_ALUT (
.I0(CLBLM_L_X8Y136_SLICE_X10Y136_A5Q),
.I1(BRAM_L_X6Y130_RAMB18_X0Y52_DO4),
.I2(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO4),
.I3(LIOB33_X0Y135_IOB_X0Y136_I),
.I4(LIOB33_X0Y147_IOB_X0Y148_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y136_SLICE_X10Y136_AO5),
.O6(CLBLM_L_X8Y136_SLICE_X10Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3300ffccffcc3300)
  ) CLBLM_L_X8Y136_SLICE_X11Y136_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y136_SLICE_X11Y136_CO6),
.I4(CLBLM_R_X7Y129_SLICE_X9Y129_B5Q),
.I5(CLBLM_R_X25Y149_SLICE_X36Y149_BQ),
.O5(CLBLM_L_X8Y136_SLICE_X11Y136_DO5),
.O6(CLBLM_L_X8Y136_SLICE_X11Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X8Y136_SLICE_X11Y136_CLUT (
.I0(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO6),
.I1(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO5),
.I2(BRAM_R_X17Y135_RAMB18_X1Y54_DO6),
.I3(BRAM_R_X17Y135_RAMB18_X1Y54_DO5),
.I4(CLBLM_R_X7Y129_SLICE_X9Y129_B5Q),
.I5(BRAM_L_X6Y135_RAMB18_X0Y54_DO6),
.O5(CLBLM_L_X8Y136_SLICE_X11Y136_CO5),
.O6(CLBLM_L_X8Y136_SLICE_X11Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h74474774b88b8bb8)
  ) CLBLM_L_X8Y136_SLICE_X11Y136_BLUT (
.I0(CLBLM_R_X7Y132_SLICE_X8Y132_A5Q),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I2(BRAM_L_X6Y135_RAMB18_X0Y54_DO7),
.I3(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO7),
.I4(CLBLM_L_X8Y136_SLICE_X11Y136_AO6),
.I5(CLBLM_L_X16Y151_SLICE_X22Y151_BQ),
.O5(CLBLM_L_X8Y136_SLICE_X11Y136_BO5),
.O6(CLBLM_L_X8Y136_SLICE_X11Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X8Y136_SLICE_X11Y136_ALUT (
.I0(CLBLM_R_X7Y132_SLICE_X8Y132_A5Q),
.I1(BRAM_L_X6Y135_RAMB18_X0Y54_DO3),
.I2(BRAM_R_X17Y135_RAMB18_X1Y54_DO4),
.I3(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO4),
.I4(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO4),
.I5(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO3),
.O5(CLBLM_L_X8Y136_SLICE_X11Y136_AO5),
.O6(CLBLM_L_X8Y136_SLICE_X11Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y137_SLICE_X10Y137_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y137_SLICE_X10Y137_AO5),
.Q(CLBLM_L_X8Y137_SLICE_X10Y137_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y137_SLICE_X10Y137_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y137_SLICE_X10Y137_BO5),
.Q(CLBLM_L_X8Y137_SLICE_X10Y137_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y137_SLICE_X10Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y137_SLICE_X10Y137_AO6),
.Q(CLBLM_L_X8Y137_SLICE_X10Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y137_SLICE_X10Y137_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y137_SLICE_X10Y137_BO6),
.Q(CLBLM_L_X8Y137_SLICE_X10Y137_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2112eddeedde2112)
  ) CLBLM_L_X8Y137_SLICE_X10Y137_DLUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y54_DO7),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I2(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO7),
.I3(CLBLM_L_X8Y137_SLICE_X10Y137_CO6),
.I4(CLBLM_L_X16Y151_SLICE_X23Y151_AQ),
.I5(CLBLM_R_X7Y136_SLICE_X8Y136_A5Q),
.O5(CLBLM_L_X8Y137_SLICE_X10Y137_DO5),
.O6(CLBLM_L_X8Y137_SLICE_X10Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X8Y137_SLICE_X10Y137_CLUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y54_DO0),
.I1(BRAM_R_X17Y135_RAMB18_X1Y54_DO1),
.I2(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO1),
.I3(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO1),
.I4(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO0),
.I5(CLBLM_R_X7Y136_SLICE_X8Y136_A5Q),
.O5(CLBLM_L_X8Y137_SLICE_X10Y137_CO5),
.O6(CLBLM_L_X8Y137_SLICE_X10Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555aaaacc5acc5a)
  ) CLBLM_L_X8Y137_SLICE_X10Y137_BLUT (
.I0(CLBLM_L_X8Y137_SLICE_X10Y137_B5Q),
.I1(LIOB33_X0Y139_IOB_X0Y139_I),
.I2(BRAM_L_X6Y130_RAMB18_X0Y52_DO7),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO7),
.I5(1'b1),
.O5(CLBLM_L_X8Y137_SLICE_X10Y137_BO5),
.O6(CLBLM_L_X8Y137_SLICE_X10Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ccccf066f066)
  ) CLBLM_L_X8Y137_SLICE_X10Y137_ALUT (
.I0(BRAM_L_X6Y130_RAMB18_X0Y52_DO6),
.I1(CLBLM_L_X8Y137_SLICE_X10Y137_A5Q),
.I2(LIOB33_X0Y137_IOB_X0Y138_I),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y137_SLICE_X10Y137_AO5),
.O6(CLBLM_L_X8Y137_SLICE_X10Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h77dd77dd22882288)
  ) CLBLM_L_X8Y137_SLICE_X11Y137_DLUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I1(CLBLM_L_X16Y149_SLICE_X22Y149_BQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y130_SLICE_X10Y130_A5Q),
.I4(1'b1),
.I5(CLBLM_L_X8Y137_SLICE_X11Y137_BO6),
.O5(CLBLM_L_X8Y137_SLICE_X11Y137_DO5),
.O6(CLBLM_L_X8Y137_SLICE_X11Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3caaaaaaaa)
  ) CLBLM_L_X8Y137_SLICE_X11Y137_CLUT (
.I0(CLBLM_L_X8Y137_SLICE_X11Y137_AO6),
.I1(CLBLM_R_X5Y134_SLICE_X7Y134_A5Q),
.I2(CLBLM_R_X25Y151_SLICE_X36Y151_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.O5(CLBLM_L_X8Y137_SLICE_X11Y137_CO5),
.O6(CLBLM_L_X8Y137_SLICE_X11Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X8Y137_SLICE_X11Y137_BLUT (
.I0(BRAM_R_X17Y135_RAMB18_X1Y54_DO6),
.I1(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO6),
.I2(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO7),
.I3(BRAM_R_X17Y135_RAMB18_X1Y54_DO7),
.I4(BRAM_L_X6Y135_RAMB18_X0Y54_DO7),
.I5(CLBLM_L_X8Y130_SLICE_X10Y130_A5Q),
.O5(CLBLM_L_X8Y137_SLICE_X11Y137_BO5),
.O6(CLBLM_L_X8Y137_SLICE_X11Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X8Y137_SLICE_X11Y137_ALUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO7),
.I1(BRAM_L_X6Y135_RAMB18_X0Y54_DO6),
.I2(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO7),
.I3(BRAM_R_X17Y135_RAMB18_X1Y54_DO7),
.I4(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO6),
.I5(CLBLM_R_X5Y134_SLICE_X7Y134_A5Q),
.O5(CLBLM_L_X8Y137_SLICE_X11Y137_AO5),
.O6(CLBLM_L_X8Y137_SLICE_X11Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y138_SLICE_X10Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.Q(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y138_SLICE_X10Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y138_SLICE_X10Y138_DO5),
.O6(CLBLM_L_X8Y138_SLICE_X10Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y138_SLICE_X10Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y138_SLICE_X10Y138_CO5),
.O6(CLBLM_L_X8Y138_SLICE_X10Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y138_SLICE_X10Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y138_SLICE_X10Y138_BO5),
.O6(CLBLM_L_X8Y138_SLICE_X10Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0ff0f0f0f0)
  ) CLBLM_L_X8Y138_SLICE_X10Y138_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO3),
.O5(CLBLM_L_X8Y138_SLICE_X10Y138_AO5),
.O6(CLBLM_L_X8Y138_SLICE_X10Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y138_SLICE_X11Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y138_SLICE_X11Y138_DO5),
.O6(CLBLM_L_X8Y138_SLICE_X11Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y138_SLICE_X11Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y138_SLICE_X11Y138_CO5),
.O6(CLBLM_L_X8Y138_SLICE_X11Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y138_SLICE_X11Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y138_SLICE_X11Y138_BO5),
.O6(CLBLM_L_X8Y138_SLICE_X11Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y138_SLICE_X11Y138_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y138_SLICE_X11Y138_AO5),
.O6(CLBLM_L_X8Y138_SLICE_X11Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y130_SLICE_X12Y130_AO6),
.Q(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y130_SLICE_X12Y130_BO6),
.Q(CLBLM_L_X10Y130_SLICE_X12Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X12Y130_DO5),
.O6(CLBLM_L_X10Y130_SLICE_X12Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X12Y130_CO5),
.O6(CLBLM_L_X10Y130_SLICE_X12Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3c3c3c3c3c)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y131_SLICE_X3Y131_CQ),
.I2(BRAM_R_X17Y135_RAMB18_X1Y54_DO18),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X12Y130_BO5),
.O6(CLBLM_L_X10Y130_SLICE_X12Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa55aa55aa55aa)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_ALUT (
.I0(BRAM_R_X17Y135_RAMB18_X1Y54_DO16),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X3Y131_SLICE_X3Y131_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X12Y130_AO5),
.O6(CLBLM_L_X10Y130_SLICE_X12Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X13Y130_DO5),
.O6(CLBLM_L_X10Y130_SLICE_X13Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X13Y130_CO5),
.O6(CLBLM_L_X10Y130_SLICE_X13Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X13Y130_BO5),
.O6(CLBLM_L_X10Y130_SLICE_X13Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X13Y130_AO5),
.O6(CLBLM_L_X10Y130_SLICE_X13Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y131_SLICE_X12Y131_AO6),
.Q(CLBLM_L_X10Y131_SLICE_X12Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y131_SLICE_X12Y131_DO5),
.O6(CLBLM_L_X10Y131_SLICE_X12Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y131_SLICE_X12Y131_CO5),
.O6(CLBLM_L_X10Y131_SLICE_X12Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y131_SLICE_X12Y131_BO5),
.O6(CLBLM_L_X10Y131_SLICE_X12Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff00ff00ff00ff0)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X5Y130_SLICE_X6Y130_DQ),
.I3(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO2),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y131_SLICE_X12Y131_AO5),
.O6(CLBLM_L_X10Y131_SLICE_X12Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y131_SLICE_X13Y131_AO6),
.Q(CLBLM_L_X10Y131_SLICE_X13Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y131_SLICE_X13Y131_DO5),
.O6(CLBLM_L_X10Y131_SLICE_X13Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y131_SLICE_X13Y131_CO5),
.O6(CLBLM_L_X10Y131_SLICE_X13Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y131_SLICE_X13Y131_BO5),
.O6(CLBLM_L_X10Y131_SLICE_X13Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ffff00ff00)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(BRAM_R_X17Y135_RAMB18_X1Y54_DO22),
.I4(1'b1),
.I5(CLBLM_R_X3Y132_SLICE_X2Y132_CQ),
.O5(CLBLM_L_X10Y131_SLICE_X13Y131_AO5),
.O6(CLBLM_L_X10Y131_SLICE_X13Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y132_SLICE_X12Y132_AO6),
.Q(CLBLM_L_X10Y132_SLICE_X12Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y132_SLICE_X12Y132_BO6),
.Q(CLBLM_L_X10Y132_SLICE_X12Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y132_SLICE_X12Y132_CO6),
.Q(CLBLM_L_X10Y132_SLICE_X12Y132_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y132_SLICE_X12Y132_DO6),
.Q(CLBLM_L_X10Y132_SLICE_X12Y132_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5a5a5a5a5a)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_DLUT (
.I0(CLBLL_L_X4Y133_SLICE_X5Y133_AQ),
.I1(1'b1),
.I2(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO7),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_DO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555555aaaaaaaa)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_CLUT (
.I0(CLBLM_R_X5Y132_SLICE_X6Y132_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO5),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_CO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3c3c3c3c3c)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.I2(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO4),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_BO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555555aaaaaaaa)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_ALUT (
.I0(CLBLL_L_X4Y131_SLICE_X5Y131_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(BRAM_L_X6Y135_RAMB18_X0Y54_DO20),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_AO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_DO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_CO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_BO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_AO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y133_SLICE_X12Y133_DO5),
.O6(CLBLM_L_X10Y133_SLICE_X12Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y133_SLICE_X12Y133_CO5),
.O6(CLBLM_L_X10Y133_SLICE_X12Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y133_SLICE_X12Y133_BO5),
.O6(CLBLM_L_X10Y133_SLICE_X12Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y133_SLICE_X12Y133_AO5),
.O6(CLBLM_L_X10Y133_SLICE_X12Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y133_SLICE_X13Y133_AO6),
.Q(CLBLM_L_X10Y133_SLICE_X13Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y133_SLICE_X13Y133_BO6),
.Q(CLBLM_L_X10Y133_SLICE_X13Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y133_SLICE_X13Y133_CO6),
.Q(CLBLM_L_X10Y133_SLICE_X13Y133_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y133_SLICE_X13Y133_DO5),
.O6(CLBLM_L_X10Y133_SLICE_X13Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cc33cc33cc33cc)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y132_SLICE_X7Y132_A5Q),
.I2(1'b1),
.I3(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y133_SLICE_X13Y133_CO5),
.O6(CLBLM_L_X10Y133_SLICE_X13Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ffff00ff00)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO4),
.I4(1'b1),
.I5(CLBLM_R_X5Y131_SLICE_X6Y131_A5Q),
.O5(CLBLM_L_X10Y133_SLICE_X13Y133_BO5),
.O6(CLBLM_L_X10Y133_SLICE_X13Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555555aaaaaaaa)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_ALUT (
.I0(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO0),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y130_SLICE_X6Y130_CQ),
.O5(CLBLM_L_X10Y133_SLICE_X13Y133_AO5),
.O6(CLBLM_L_X10Y133_SLICE_X13Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y134_SLICE_X12Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y134_SLICE_X12Y134_DO5),
.O6(CLBLM_L_X10Y134_SLICE_X12Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7b7b7b7b48484848)
  ) CLBLM_L_X10Y134_SLICE_X12Y134_CLUT (
.I0(CLBLM_R_X3Y131_SLICE_X3Y131_CQ),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I2(CLBLM_R_X3Y155_SLICE_X2Y155_DQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X8Y134_SLICE_X10Y134_BO6),
.O5(CLBLM_L_X10Y134_SLICE_X12Y134_CO5),
.O6(CLBLM_L_X10Y134_SLICE_X12Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff00ff099996666)
  ) CLBLM_L_X10Y134_SLICE_X12Y134_BLUT (
.I0(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO7),
.I1(BRAM_L_X6Y135_RAMB18_X0Y54_DO7),
.I2(CLBLM_L_X16Y153_SLICE_X22Y153_AQ),
.I3(CLBLM_R_X7Y134_SLICE_X9Y134_B5Q),
.I4(CLBLM_L_X10Y134_SLICE_X12Y134_AO6),
.I5(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.O5(CLBLM_L_X10Y134_SLICE_X12Y134_BO5),
.O6(CLBLM_L_X10Y134_SLICE_X12Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X10Y134_SLICE_X12Y134_ALUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO3),
.I1(BRAM_L_X6Y135_RAMB18_X0Y54_DO3),
.I2(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO2),
.I3(BRAM_R_X17Y135_RAMB18_X1Y54_DO3),
.I4(BRAM_L_X6Y135_RAMB18_X0Y54_DO2),
.I5(CLBLM_R_X7Y134_SLICE_X9Y134_B5Q),
.O5(CLBLM_L_X10Y134_SLICE_X12Y134_AO5),
.O6(CLBLM_L_X10Y134_SLICE_X12Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y134_SLICE_X13Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y134_SLICE_X13Y134_DO5),
.O6(CLBLM_L_X10Y134_SLICE_X13Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y134_SLICE_X13Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y134_SLICE_X13Y134_CO5),
.O6(CLBLM_L_X10Y134_SLICE_X13Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h74474774b88b8bb8)
  ) CLBLM_L_X10Y134_SLICE_X13Y134_BLUT (
.I0(CLBLM_L_X16Y149_SLICE_X22Y149_AQ),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I2(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO7),
.I3(BRAM_R_X17Y135_RAMB18_X1Y54_DO7),
.I4(CLBLM_L_X10Y134_SLICE_X13Y134_AO6),
.I5(CLBLM_R_X7Y129_SLICE_X9Y129_A5Q),
.O5(CLBLM_L_X10Y134_SLICE_X13Y134_BO5),
.O6(CLBLM_L_X10Y134_SLICE_X13Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X10Y134_SLICE_X13Y134_ALUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO3),
.I1(BRAM_R_X17Y135_RAMB18_X1Y54_DO3),
.I2(BRAM_R_X17Y135_RAMB18_X1Y54_DO4),
.I3(BRAM_L_X6Y135_RAMB18_X0Y54_DO4),
.I4(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO4),
.I5(CLBLM_R_X7Y129_SLICE_X9Y129_A5Q),
.O5(CLBLM_L_X10Y134_SLICE_X13Y134_AO5),
.O6(CLBLM_L_X10Y134_SLICE_X13Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y135_SLICE_X12Y135_AO5),
.Q(CLBLM_L_X10Y135_SLICE_X12Y135_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y135_SLICE_X12Y135_AO6),
.Q(CLBLM_L_X10Y135_SLICE_X12Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_DLUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y54_DO4),
.I1(BRAM_L_X6Y135_RAMB18_X0Y54_DO5),
.I2(BRAM_R_X17Y135_RAMB18_X1Y54_DO5),
.I3(CLBLM_L_X10Y135_SLICE_X12Y135_A5Q),
.I4(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO5),
.I5(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO4),
.O5(CLBLM_L_X10Y135_SLICE_X12Y135_DO5),
.O6(CLBLM_L_X10Y135_SLICE_X12Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_CLUT (
.I0(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO2),
.I1(CLBLM_R_X5Y130_SLICE_X6Y130_AQ),
.I2(BRAM_R_X17Y135_RAMB18_X1Y54_DO2),
.I3(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO3),
.I4(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO3),
.I5(BRAM_L_X6Y135_RAMB18_X0Y54_DO3),
.O5(CLBLM_L_X10Y135_SLICE_X12Y135_CO5),
.O6(CLBLM_L_X10Y135_SLICE_X12Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_BLUT (
.I0(BRAM_R_X17Y135_RAMB18_X1Y54_DO4),
.I1(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO5),
.I2(CLBLM_R_X3Y133_SLICE_X3Y133_AQ),
.I3(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO4),
.I4(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO5),
.I5(BRAM_L_X6Y135_RAMB18_X0Y54_DO5),
.O5(CLBLM_L_X10Y135_SLICE_X12Y135_BO5),
.O6(CLBLM_L_X10Y135_SLICE_X12Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffff008d8dd8d8)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_ALUT (
.I0(LIOB33_X0Y147_IOB_X0Y148_I),
.I1(LIOB33_X0Y137_IOB_X0Y137_I),
.I2(BRAM_L_X6Y130_RAMB18_X0Y52_DO5),
.I3(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO5),
.I4(CLBLM_L_X10Y135_SLICE_X12Y135_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y135_SLICE_X12Y135_AO5),
.O6(CLBLM_L_X10Y135_SLICE_X12Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_DLUT (
.I0(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO0),
.I1(BRAM_L_X6Y135_RAMB18_X0Y54_DO1),
.I2(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO1),
.I3(CLBLM_L_X8Y135_SLICE_X10Y135_A5Q),
.I4(BRAM_R_X17Y135_RAMB18_X1Y54_DO1),
.I5(BRAM_L_X6Y135_RAMB18_X0Y54_DO0),
.O5(CLBLM_L_X10Y135_SLICE_X13Y135_DO5),
.O6(CLBLM_L_X10Y135_SLICE_X13Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_CLUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y54_DO2),
.I1(BRAM_L_X6Y135_RAMB18_X0Y54_DO1),
.I2(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO1),
.I3(BRAM_R_X17Y135_RAMB18_X1Y54_DO2),
.I4(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO2),
.I5(CLBLM_R_X7Y134_SLICE_X9Y134_A5Q),
.O5(CLBLM_L_X10Y135_SLICE_X13Y135_CO5),
.O6(CLBLM_L_X10Y135_SLICE_X13Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_BLUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO1),
.I1(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO0),
.I2(CLBLL_L_X4Y132_SLICE_X4Y132_AQ),
.I3(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO1),
.I4(BRAM_R_X17Y135_RAMB18_X1Y54_DO0),
.I5(BRAM_L_X6Y135_RAMB18_X0Y54_DO1),
.O5(CLBLM_L_X10Y135_SLICE_X13Y135_BO5),
.O6(CLBLM_L_X10Y135_SLICE_X13Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_ALUT (
.I0(CLBLM_R_X3Y132_SLICE_X3Y132_AQ),
.I1(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO3),
.I2(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO4),
.I3(BRAM_L_X6Y135_RAMB18_X0Y54_DO4),
.I4(BRAM_R_X17Y135_RAMB18_X1Y54_DO3),
.I5(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO4),
.O5(CLBLM_L_X10Y135_SLICE_X13Y135_AO5),
.O6(CLBLM_L_X10Y135_SLICE_X13Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1441beebebbe4114)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_DLUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I1(CLBLM_L_X10Y136_SLICE_X13Y136_AO5),
.I2(CLBLM_L_X10Y136_SLICE_X13Y136_BO5),
.I3(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO0),
.I4(CLBLM_R_X25Y149_SLICE_X37Y149_AQ),
.I5(CLBLM_R_X7Y129_SLICE_X8Y129_A5Q),
.O5(CLBLM_L_X10Y136_SLICE_X12Y136_DO5),
.O6(CLBLM_L_X10Y136_SLICE_X12Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33a5cca5335acc5a)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_CLUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y54_DO7),
.I1(CLBLM_L_X8Y136_SLICE_X10Y136_A5Q),
.I2(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO7),
.I3(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I4(CLBLM_L_X16Y154_SLICE_X22Y154_AQ),
.I5(CLBLM_L_X10Y136_SLICE_X12Y136_BO6),
.O5(CLBLM_L_X10Y136_SLICE_X12Y136_CO5),
.O6(CLBLM_L_X10Y136_SLICE_X12Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_BLUT (
.I0(BRAM_R_X17Y135_RAMB18_X1Y54_DO4),
.I1(BRAM_L_X6Y135_RAMB18_X0Y54_DO3),
.I2(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO3),
.I3(BRAM_L_X6Y135_RAMB18_X0Y54_DO4),
.I4(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO4),
.I5(CLBLM_L_X8Y136_SLICE_X10Y136_A5Q),
.O5(CLBLM_L_X10Y136_SLICE_X12Y136_BO5),
.O6(CLBLM_L_X10Y136_SLICE_X12Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_ALUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y54_DO6),
.I1(CLBLM_L_X8Y137_SLICE_X10Y137_A5Q),
.I2(BRAM_R_X17Y135_RAMB18_X1Y54_DO6),
.I3(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO5),
.I4(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO6),
.I5(BRAM_L_X6Y135_RAMB18_X0Y54_DO5),
.O5(CLBLM_L_X10Y136_SLICE_X12Y136_AO5),
.O6(CLBLM_L_X10Y136_SLICE_X12Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h12ed21dede21ed12)
  ) CLBLM_L_X10Y136_SLICE_X13Y136_DLUT (
.I0(CLBLM_L_X10Y136_SLICE_X13Y136_AO6),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I2(BRAM_L_X6Y135_RAMB18_X0Y54_DO0),
.I3(CLBLM_L_X8Y132_SLICE_X11Y132_A5Q),
.I4(CLBLM_L_X10Y136_SLICE_X13Y136_BO5),
.I5(CLBLM_L_X16Y152_SLICE_X22Y152_AQ),
.O5(CLBLM_L_X10Y136_SLICE_X13Y136_DO5),
.O6(CLBLM_L_X10Y136_SLICE_X13Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X10Y136_SLICE_X13Y136_CLUT (
.I0(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO2),
.I1(BRAM_R_X17Y135_RAMB18_X1Y54_DO1),
.I2(CLBLM_R_X3Y131_SLICE_X3Y131_B5Q),
.I3(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO1),
.I4(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO2),
.I5(BRAM_L_X6Y135_RAMB18_X0Y54_DO2),
.O5(CLBLM_L_X10Y136_SLICE_X13Y136_CO5),
.O6(CLBLM_L_X10Y136_SLICE_X13Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3c66666666)
  ) CLBLM_L_X10Y136_SLICE_X13Y136_BLUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO0),
.I1(BRAM_R_X17Y135_RAMB18_X1Y54_DO0),
.I2(CLBLM_R_X3Y131_SLICE_X3Y131_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y136_SLICE_X13Y136_BO5),
.O6(CLBLM_L_X10Y136_SLICE_X13Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff00ff05a5a5a5a)
  ) CLBLM_L_X10Y136_SLICE_X13Y136_ALUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO7),
.I1(1'b1),
.I2(BRAM_L_X6Y135_RAMB18_X0Y54_DO7),
.I3(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO7),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y136_SLICE_X13Y136_AO5),
.O6(CLBLM_L_X10Y136_SLICE_X13Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777dddd22228888)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_DLUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I1(CLBLM_R_X7Y128_SLICE_X8Y128_A5Q),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X25Y149_SLICE_X36Y149_AQ),
.I5(CLBLM_L_X10Y137_SLICE_X12Y137_BO6),
.O5(CLBLM_L_X10Y137_SLICE_X12Y137_DO5),
.O6(CLBLM_L_X10Y137_SLICE_X12Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f0af5a05f0af5a0)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_CLUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I1(1'b1),
.I2(CLBLM_R_X25Y151_SLICE_X36Y151_BQ),
.I3(CLBLM_L_X10Y137_SLICE_X12Y137_AO6),
.I4(CLBLM_R_X7Y137_SLICE_X8Y137_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y137_SLICE_X12Y137_CO5),
.O6(CLBLM_L_X10Y137_SLICE_X12Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_BLUT (
.I0(CLBLM_R_X7Y128_SLICE_X8Y128_A5Q),
.I1(BRAM_R_X17Y135_RAMB18_X1Y54_DO5),
.I2(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO4),
.I3(BRAM_R_X17Y135_RAMB18_X1Y54_DO4),
.I4(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO5),
.I5(BRAM_L_X6Y135_RAMB18_X0Y54_DO5),
.O5(CLBLM_L_X10Y137_SLICE_X12Y137_BO5),
.O6(CLBLM_L_X10Y137_SLICE_X12Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_ALUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO6),
.I1(CLBLM_R_X7Y137_SLICE_X8Y137_A5Q),
.I2(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO5),
.I3(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO6),
.I4(BRAM_R_X17Y135_RAMB18_X1Y54_DO6),
.I5(BRAM_L_X6Y135_RAMB18_X0Y54_DO5),
.O5(CLBLM_L_X10Y137_SLICE_X12Y137_AO5),
.O6(CLBLM_L_X10Y137_SLICE_X12Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y137_SLICE_X13Y137_DO5),
.O6(CLBLM_L_X10Y137_SLICE_X13Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y137_SLICE_X13Y137_CO5),
.O6(CLBLM_L_X10Y137_SLICE_X13Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6f6f60606f6f6060)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_BLUT (
.I0(CLBLM_L_X16Y151_SLICE_X22Y151_CQ),
.I1(CLBLM_R_X7Y131_SLICE_X9Y131_A5Q),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y137_SLICE_X13Y137_AO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y137_SLICE_X13Y137_BO5),
.O6(CLBLM_L_X10Y137_SLICE_X13Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_ALUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO4),
.I1(CLBLM_R_X7Y131_SLICE_X9Y131_A5Q),
.I2(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO5),
.I3(BRAM_L_X6Y135_RAMB18_X0Y54_DO4),
.I4(BRAM_R_X17Y135_RAMB18_X1Y54_DO5),
.I5(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO5),
.O5(CLBLM_L_X10Y137_SLICE_X13Y137_AO5),
.O6(CLBLM_L_X10Y137_SLICE_X13Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y138_SLICE_X12Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(LIOB33_X0Y147_IOB_X0Y148_I),
.Q(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y138_SLICE_X12Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y138_SLICE_X12Y138_DO5),
.O6(CLBLM_L_X10Y138_SLICE_X12Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y138_SLICE_X12Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y138_SLICE_X12Y138_CO5),
.O6(CLBLM_L_X10Y138_SLICE_X12Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y138_SLICE_X12Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y138_SLICE_X12Y138_BO5),
.O6(CLBLM_L_X10Y138_SLICE_X12Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y138_SLICE_X12Y138_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y138_SLICE_X12Y138_AO5),
.O6(CLBLM_L_X10Y138_SLICE_X12Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y138_SLICE_X13Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y138_SLICE_X13Y138_DO5),
.O6(CLBLM_L_X10Y138_SLICE_X13Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y138_SLICE_X13Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y138_SLICE_X13Y138_CO5),
.O6(CLBLM_L_X10Y138_SLICE_X13Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y138_SLICE_X13Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y138_SLICE_X13Y138_BO5),
.O6(CLBLM_L_X10Y138_SLICE_X13Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y138_SLICE_X13Y138_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y138_SLICE_X13Y138_AO5),
.O6(CLBLM_L_X10Y138_SLICE_X13Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y130_SLICE_X16Y130_AO6),
.Q(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y130_SLICE_X16Y130_DO5),
.O6(CLBLM_L_X12Y130_SLICE_X16Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y130_SLICE_X16Y130_CO5),
.O6(CLBLM_L_X12Y130_SLICE_X16Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y130_SLICE_X16Y130_BO5),
.O6(CLBLM_L_X12Y130_SLICE_X16Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa55aa55aa55aa)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_ALUT (
.I0(BRAM_R_X17Y135_RAMB18_X1Y54_DO19),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y130_SLICE_X16Y130_AO5),
.O6(CLBLM_L_X12Y130_SLICE_X16Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y130_SLICE_X17Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y130_SLICE_X17Y130_DO5),
.O6(CLBLM_L_X12Y130_SLICE_X17Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y130_SLICE_X17Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y130_SLICE_X17Y130_CO5),
.O6(CLBLM_L_X12Y130_SLICE_X17Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y130_SLICE_X17Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y130_SLICE_X17Y130_BO5),
.O6(CLBLM_L_X12Y130_SLICE_X17Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y130_SLICE_X17Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y130_SLICE_X17Y130_AO5),
.O6(CLBLM_L_X12Y130_SLICE_X17Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y132_SLICE_X16Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y132_SLICE_X16Y132_AO6),
.Q(CLBLM_L_X12Y132_SLICE_X16Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y132_SLICE_X16Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y132_SLICE_X16Y132_BO6),
.Q(CLBLM_L_X12Y132_SLICE_X16Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y132_SLICE_X16Y132_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y132_SLICE_X16Y132_CO6),
.Q(CLBLM_L_X12Y132_SLICE_X16Y132_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y132_SLICE_X16Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y132_SLICE_X16Y132_DO5),
.O6(CLBLM_L_X12Y132_SLICE_X16Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff00ff00ff00ff0)
  ) CLBLM_L_X12Y132_SLICE_X16Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X3Y132_SLICE_X3Y132_BQ),
.I3(BRAM_R_X17Y135_RAMB18_X1Y54_DO21),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y132_SLICE_X16Y132_CO5),
.O6(CLBLM_L_X12Y132_SLICE_X16Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ffff00ff00)
  ) CLBLM_L_X12Y132_SLICE_X16Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO7),
.I4(1'b1),
.I5(CLBLL_L_X4Y132_SLICE_X5Y132_A5Q),
.O5(CLBLM_L_X12Y132_SLICE_X16Y132_BO5),
.O6(CLBLM_L_X12Y132_SLICE_X16Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0ff0f0f0f0)
  ) CLBLM_L_X12Y132_SLICE_X16Y132_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X7Y130_SLICE_X8Y130_B5Q),
.I3(1'b1),
.I4(1'b1),
.I5(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO1),
.O5(CLBLM_L_X12Y132_SLICE_X16Y132_AO5),
.O6(CLBLM_L_X12Y132_SLICE_X16Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y132_SLICE_X17Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y132_SLICE_X17Y132_DO5),
.O6(CLBLM_L_X12Y132_SLICE_X17Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y132_SLICE_X17Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y132_SLICE_X17Y132_CO5),
.O6(CLBLM_L_X12Y132_SLICE_X17Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y132_SLICE_X17Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y132_SLICE_X17Y132_BO5),
.O6(CLBLM_L_X12Y132_SLICE_X17Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y132_SLICE_X17Y132_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y132_SLICE_X17Y132_AO5),
.O6(CLBLM_L_X12Y132_SLICE_X17Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y135_SLICE_X16Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y135_SLICE_X16Y135_DO5),
.O6(CLBLM_L_X12Y135_SLICE_X16Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y135_SLICE_X16Y135_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y135_SLICE_X16Y135_CO5),
.O6(CLBLM_L_X12Y135_SLICE_X16Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5ff55ff50aa00aa0)
  ) CLBLM_L_X12Y135_SLICE_X16Y135_BLUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I1(1'b1),
.I2(CLBLM_L_X16Y152_SLICE_X22Y152_BQ),
.I3(CLBLM_R_X7Y134_SLICE_X9Y134_A5Q),
.I4(1'b1),
.I5(CLBLM_L_X10Y135_SLICE_X13Y135_CO6),
.O5(CLBLM_L_X12Y135_SLICE_X16Y135_BO5),
.O6(CLBLM_L_X12Y135_SLICE_X16Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h77dd77dd22882288)
  ) CLBLM_L_X12Y135_SLICE_X16Y135_ALUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I1(CLBLM_R_X25Y154_SLICE_X36Y154_AQ),
.I2(1'b1),
.I3(CLBLM_R_X3Y131_SLICE_X3Y131_AQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y135_SLICE_X14Y135_AO6),
.O5(CLBLM_L_X12Y135_SLICE_X16Y135_AO5),
.O6(CLBLM_L_X12Y135_SLICE_X16Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y135_SLICE_X17Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y135_SLICE_X17Y135_DO5),
.O6(CLBLM_L_X12Y135_SLICE_X17Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y135_SLICE_X17Y135_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y135_SLICE_X17Y135_CO5),
.O6(CLBLM_L_X12Y135_SLICE_X17Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y135_SLICE_X17Y135_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y135_SLICE_X17Y135_BO5),
.O6(CLBLM_L_X12Y135_SLICE_X17Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y135_SLICE_X17Y135_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y135_SLICE_X17Y135_AO5),
.O6(CLBLM_L_X12Y135_SLICE_X17Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y135_SLICE_X22Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X16Y135_SLICE_X22Y135_AO6),
.Q(CLBLM_L_X16Y135_SLICE_X22Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y135_SLICE_X22Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X16Y135_SLICE_X22Y135_BO6),
.Q(CLBLM_L_X16Y135_SLICE_X22Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5c53aca3535ca3ac)
  ) CLBLM_L_X16Y135_SLICE_X22Y135_DLUT (
.I0(CLBLM_R_X5Y130_SLICE_X6Y130_AQ),
.I1(BRAM_R_X17Y135_RAMB18_X1Y54_DO7),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I3(CLBLM_L_X10Y135_SLICE_X12Y135_CO6),
.I4(CLBLM_L_X16Y157_SLICE_X22Y157_AQ),
.I5(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO7),
.O5(CLBLM_L_X16Y135_SLICE_X22Y135_DO5),
.O6(CLBLM_L_X16Y135_SLICE_X22Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff099990ff06666)
  ) CLBLM_L_X16Y135_SLICE_X22Y135_CLUT (
.I0(CLBLM_L_X10Y135_SLICE_X13Y135_AO6),
.I1(BRAM_R_X17Y135_RAMB18_X1Y54_DO7),
.I2(CLBLM_R_X3Y132_SLICE_X3Y132_AQ),
.I3(CLBLM_R_X25Y157_SLICE_X36Y157_BQ),
.I4(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I5(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO7),
.O5(CLBLM_L_X16Y135_SLICE_X22Y135_CO5),
.O6(CLBLM_L_X16Y135_SLICE_X22Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa55aa55aa55aa)
  ) CLBLM_L_X16Y135_SLICE_X22Y135_BLUT (
.I0(CLBLM_R_X3Y132_SLICE_X3Y132_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(BRAM_R_X17Y135_RAMB18_X1Y54_DO4),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y135_SLICE_X22Y135_BO5),
.O6(CLBLM_L_X16Y135_SLICE_X22Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3c3c3c3c3c)
  ) CLBLM_L_X16Y135_SLICE_X22Y135_ALUT (
.I0(1'b1),
.I1(BRAM_R_X17Y135_RAMB18_X1Y54_DO3),
.I2(CLBLM_R_X5Y130_SLICE_X6Y130_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y135_SLICE_X22Y135_AO5),
.O6(CLBLM_L_X16Y135_SLICE_X22Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y135_SLICE_X23Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y135_SLICE_X23Y135_DO5),
.O6(CLBLM_L_X16Y135_SLICE_X23Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y135_SLICE_X23Y135_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y135_SLICE_X23Y135_CO5),
.O6(CLBLM_L_X16Y135_SLICE_X23Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y135_SLICE_X23Y135_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y135_SLICE_X23Y135_BO5),
.O6(CLBLM_L_X16Y135_SLICE_X23Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y135_SLICE_X23Y135_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y135_SLICE_X23Y135_AO5),
.O6(CLBLM_L_X16Y135_SLICE_X23Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y136_SLICE_X22Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X16Y136_SLICE_X22Y136_AO6),
.Q(CLBLM_L_X16Y136_SLICE_X22Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5c5cacac5c5cacac)
  ) CLBLM_L_X16Y136_SLICE_X22Y136_DLUT (
.I0(CLBLM_L_X16Y155_SLICE_X22Y155_AQ),
.I1(CLBLM_L_X10Y136_SLICE_X13Y136_CO6),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I3(1'b1),
.I4(CLBLM_R_X3Y131_SLICE_X3Y131_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X16Y136_SLICE_X22Y136_DO5),
.O6(CLBLM_L_X16Y136_SLICE_X22Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0afa0afafa0afa0a)
  ) CLBLM_L_X16Y136_SLICE_X22Y136_CLUT (
.I0(CLBLM_R_X11Y136_SLICE_X14Y136_BO6),
.I1(1'b1),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I3(CLBLM_R_X25Y154_SLICE_X36Y154_BQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y132_SLICE_X2Y132_AQ),
.O5(CLBLM_L_X16Y136_SLICE_X22Y136_CO5),
.O6(CLBLM_L_X16Y136_SLICE_X22Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5ff55ff50aa00aa0)
  ) CLBLM_L_X16Y136_SLICE_X22Y136_BLUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I1(1'b1),
.I2(CLBLM_R_X3Y132_SLICE_X2Y132_BQ),
.I3(CLBLM_R_X25Y154_SLICE_X36Y154_CQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y136_SLICE_X14Y136_AO6),
.O5(CLBLM_L_X16Y136_SLICE_X22Y136_BO5),
.O6(CLBLM_L_X16Y136_SLICE_X22Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa55aa55aa55aa)
  ) CLBLM_L_X16Y136_SLICE_X22Y136_ALUT (
.I0(CLBLM_R_X3Y131_SLICE_X3Y131_B5Q),
.I1(1'b1),
.I2(1'b1),
.I3(BRAM_R_X17Y135_RAMB18_X1Y54_DO2),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y136_SLICE_X22Y136_AO5),
.O6(CLBLM_L_X16Y136_SLICE_X22Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y136_SLICE_X23Y136_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y136_SLICE_X23Y136_DO5),
.O6(CLBLM_L_X16Y136_SLICE_X23Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y136_SLICE_X23Y136_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y136_SLICE_X23Y136_CO5),
.O6(CLBLM_L_X16Y136_SLICE_X23Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y136_SLICE_X23Y136_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y136_SLICE_X23Y136_BO5),
.O6(CLBLM_L_X16Y136_SLICE_X23Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y136_SLICE_X23Y136_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y136_SLICE_X23Y136_AO5),
.O6(CLBLM_L_X16Y136_SLICE_X23Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y137_SLICE_X22Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X16Y137_SLICE_X22Y137_AO6),
.Q(CLBLM_L_X16Y137_SLICE_X22Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y137_SLICE_X22Y137_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X16Y137_SLICE_X22Y137_BO6),
.Q(CLBLM_L_X16Y137_SLICE_X22Y137_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y137_SLICE_X22Y137_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y137_SLICE_X22Y137_DO5),
.O6(CLBLM_L_X16Y137_SLICE_X22Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y137_SLICE_X22Y137_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y137_SLICE_X22Y137_CO5),
.O6(CLBLM_L_X16Y137_SLICE_X22Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3c3c3c3c3c)
  ) CLBLM_L_X16Y137_SLICE_X22Y137_BLUT (
.I0(1'b1),
.I1(BRAM_R_X17Y135_RAMB18_X1Y54_DO7),
.I2(CLBLM_R_X3Y132_SLICE_X2Y132_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y137_SLICE_X22Y137_BO5),
.O6(CLBLM_L_X16Y137_SLICE_X22Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff00ff00ff00ff0)
  ) CLBLM_L_X16Y137_SLICE_X22Y137_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(BRAM_R_X17Y135_RAMB18_X1Y54_DO6),
.I3(CLBLM_R_X3Y132_SLICE_X2Y132_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y137_SLICE_X22Y137_AO5),
.O6(CLBLM_L_X16Y137_SLICE_X22Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y137_SLICE_X23Y137_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y137_SLICE_X23Y137_DO5),
.O6(CLBLM_L_X16Y137_SLICE_X23Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y137_SLICE_X23Y137_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y137_SLICE_X23Y137_CO5),
.O6(CLBLM_L_X16Y137_SLICE_X23Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y137_SLICE_X23Y137_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y137_SLICE_X23Y137_BO5),
.O6(CLBLM_L_X16Y137_SLICE_X23Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y137_SLICE_X23Y137_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y137_SLICE_X23Y137_AO5),
.O6(CLBLM_L_X16Y137_SLICE_X23Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y149_SLICE_X22Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(RIOB33_X105Y177_IOB_X1Y178_I),
.Q(CLBLM_L_X16Y149_SLICE_X22Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y149_SLICE_X22Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(RIOB33_X105Y181_IOB_X1Y181_I),
.Q(CLBLM_L_X16Y149_SLICE_X22Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y149_SLICE_X22Y149_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y149_SLICE_X22Y149_DO5),
.O6(CLBLM_L_X16Y149_SLICE_X22Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y149_SLICE_X22Y149_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y149_SLICE_X22Y149_CO5),
.O6(CLBLM_L_X16Y149_SLICE_X22Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y149_SLICE_X22Y149_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y149_SLICE_X22Y149_BO5),
.O6(CLBLM_L_X16Y149_SLICE_X22Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y149_SLICE_X22Y149_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y149_SLICE_X22Y149_AO5),
.O6(CLBLM_L_X16Y149_SLICE_X22Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y149_SLICE_X23Y149_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y149_SLICE_X23Y149_DO5),
.O6(CLBLM_L_X16Y149_SLICE_X23Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y149_SLICE_X23Y149_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y149_SLICE_X23Y149_CO5),
.O6(CLBLM_L_X16Y149_SLICE_X23Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y149_SLICE_X23Y149_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y149_SLICE_X23Y149_BO5),
.O6(CLBLM_L_X16Y149_SLICE_X23Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y149_SLICE_X23Y149_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y149_SLICE_X23Y149_AO5),
.O6(CLBLM_L_X16Y149_SLICE_X23Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y151_SLICE_X22Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(RIOB33_X105Y185_IOB_X1Y185_I),
.Q(CLBLM_L_X16Y151_SLICE_X22Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y151_SLICE_X22Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(RIOB33_X105Y185_IOB_X1Y186_I),
.Q(CLBLM_L_X16Y151_SLICE_X22Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y151_SLICE_X22Y151_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(RIOB33_X105Y187_IOB_X1Y187_I),
.Q(CLBLM_L_X16Y151_SLICE_X22Y151_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y151_SLICE_X22Y151_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(RIOB33_X105Y191_IOB_X1Y191_I),
.Q(CLBLM_L_X16Y151_SLICE_X22Y151_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y151_SLICE_X22Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y151_SLICE_X22Y151_DO5),
.O6(CLBLM_L_X16Y151_SLICE_X22Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y151_SLICE_X22Y151_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y151_SLICE_X22Y151_CO5),
.O6(CLBLM_L_X16Y151_SLICE_X22Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y151_SLICE_X22Y151_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y151_SLICE_X22Y151_BO5),
.O6(CLBLM_L_X16Y151_SLICE_X22Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y151_SLICE_X22Y151_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y151_SLICE_X22Y151_AO5),
.O6(CLBLM_L_X16Y151_SLICE_X22Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y151_SLICE_X23Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(RIOB33_X105Y183_IOB_X1Y183_I),
.Q(CLBLM_L_X16Y151_SLICE_X23Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y151_SLICE_X23Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y151_SLICE_X23Y151_DO5),
.O6(CLBLM_L_X16Y151_SLICE_X23Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y151_SLICE_X23Y151_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y151_SLICE_X23Y151_CO5),
.O6(CLBLM_L_X16Y151_SLICE_X23Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y151_SLICE_X23Y151_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y151_SLICE_X23Y151_BO5),
.O6(CLBLM_L_X16Y151_SLICE_X23Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y151_SLICE_X23Y151_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y151_SLICE_X23Y151_AO5),
.O6(CLBLM_L_X16Y151_SLICE_X23Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y152_SLICE_X22Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(RIOB33_X105Y189_IOB_X1Y190_I),
.Q(CLBLM_L_X16Y152_SLICE_X22Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y152_SLICE_X22Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(RIOB33_X105Y191_IOB_X1Y192_I),
.Q(CLBLM_L_X16Y152_SLICE_X22Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y152_SLICE_X22Y152_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y152_SLICE_X22Y152_DO5),
.O6(CLBLM_L_X16Y152_SLICE_X22Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y152_SLICE_X22Y152_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y152_SLICE_X22Y152_CO5),
.O6(CLBLM_L_X16Y152_SLICE_X22Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y152_SLICE_X22Y152_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y152_SLICE_X22Y152_BO5),
.O6(CLBLM_L_X16Y152_SLICE_X22Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y152_SLICE_X22Y152_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y152_SLICE_X22Y152_AO5),
.O6(CLBLM_L_X16Y152_SLICE_X22Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y152_SLICE_X23Y152_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y152_SLICE_X23Y152_DO5),
.O6(CLBLM_L_X16Y152_SLICE_X23Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y152_SLICE_X23Y152_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y152_SLICE_X23Y152_CO5),
.O6(CLBLM_L_X16Y152_SLICE_X23Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y152_SLICE_X23Y152_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y152_SLICE_X23Y152_BO5),
.O6(CLBLM_L_X16Y152_SLICE_X23Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y152_SLICE_X23Y152_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y152_SLICE_X23Y152_AO5),
.O6(CLBLM_L_X16Y152_SLICE_X23Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y153_SLICE_X22Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(RIOB33_X105Y193_IOB_X1Y193_I),
.Q(CLBLM_L_X16Y153_SLICE_X22Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y153_SLICE_X22Y153_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y153_SLICE_X22Y153_DO5),
.O6(CLBLM_L_X16Y153_SLICE_X22Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y153_SLICE_X22Y153_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y153_SLICE_X22Y153_CO5),
.O6(CLBLM_L_X16Y153_SLICE_X22Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y153_SLICE_X22Y153_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y153_SLICE_X22Y153_BO5),
.O6(CLBLM_L_X16Y153_SLICE_X22Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y153_SLICE_X22Y153_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y153_SLICE_X22Y153_AO5),
.O6(CLBLM_L_X16Y153_SLICE_X22Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y153_SLICE_X23Y153_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y153_SLICE_X23Y153_DO5),
.O6(CLBLM_L_X16Y153_SLICE_X23Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y153_SLICE_X23Y153_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y153_SLICE_X23Y153_CO5),
.O6(CLBLM_L_X16Y153_SLICE_X23Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y153_SLICE_X23Y153_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y153_SLICE_X23Y153_BO5),
.O6(CLBLM_L_X16Y153_SLICE_X23Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y153_SLICE_X23Y153_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y153_SLICE_X23Y153_AO5),
.O6(CLBLM_L_X16Y153_SLICE_X23Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y154_SLICE_X22Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(RIOB33_X105Y193_IOB_X1Y194_I),
.Q(CLBLM_L_X16Y154_SLICE_X22Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y154_SLICE_X22Y154_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(RIOB33_X105Y197_IOB_X1Y197_I),
.Q(CLBLM_L_X16Y154_SLICE_X22Y154_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y154_SLICE_X22Y154_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y154_SLICE_X22Y154_DO5),
.O6(CLBLM_L_X16Y154_SLICE_X22Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y154_SLICE_X22Y154_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y154_SLICE_X22Y154_CO5),
.O6(CLBLM_L_X16Y154_SLICE_X22Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y154_SLICE_X22Y154_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y154_SLICE_X22Y154_BO5),
.O6(CLBLM_L_X16Y154_SLICE_X22Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y154_SLICE_X22Y154_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y154_SLICE_X22Y154_AO5),
.O6(CLBLM_L_X16Y154_SLICE_X22Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y154_SLICE_X23Y154_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y154_SLICE_X23Y154_DO5),
.O6(CLBLM_L_X16Y154_SLICE_X23Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y154_SLICE_X23Y154_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y154_SLICE_X23Y154_CO5),
.O6(CLBLM_L_X16Y154_SLICE_X23Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y154_SLICE_X23Y154_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y154_SLICE_X23Y154_BO5),
.O6(CLBLM_L_X16Y154_SLICE_X23Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y154_SLICE_X23Y154_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y154_SLICE_X23Y154_AO5),
.O6(CLBLM_L_X16Y154_SLICE_X23Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y155_SLICE_X22Y155_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(RIOB33_X105Y201_IOB_X1Y202_I),
.Q(CLBLM_L_X16Y155_SLICE_X22Y155_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y155_SLICE_X22Y155_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y155_SLICE_X22Y155_DO5),
.O6(CLBLM_L_X16Y155_SLICE_X22Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y155_SLICE_X22Y155_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y155_SLICE_X22Y155_CO5),
.O6(CLBLM_L_X16Y155_SLICE_X22Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y155_SLICE_X22Y155_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y155_SLICE_X22Y155_BO5),
.O6(CLBLM_L_X16Y155_SLICE_X22Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y155_SLICE_X22Y155_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y155_SLICE_X22Y155_AO5),
.O6(CLBLM_L_X16Y155_SLICE_X22Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y155_SLICE_X23Y155_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y155_SLICE_X23Y155_DO5),
.O6(CLBLM_L_X16Y155_SLICE_X23Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y155_SLICE_X23Y155_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y155_SLICE_X23Y155_CO5),
.O6(CLBLM_L_X16Y155_SLICE_X23Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y155_SLICE_X23Y155_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y155_SLICE_X23Y155_BO5),
.O6(CLBLM_L_X16Y155_SLICE_X23Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y155_SLICE_X23Y155_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y155_SLICE_X23Y155_AO5),
.O6(CLBLM_L_X16Y155_SLICE_X23Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y157_SLICE_X22Y157_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(RIOB33_X105Y203_IOB_X1Y203_I),
.Q(CLBLM_L_X16Y157_SLICE_X22Y157_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y157_SLICE_X22Y157_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y157_SLICE_X22Y157_DO5),
.O6(CLBLM_L_X16Y157_SLICE_X22Y157_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y157_SLICE_X22Y157_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y157_SLICE_X22Y157_CO5),
.O6(CLBLM_L_X16Y157_SLICE_X22Y157_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y157_SLICE_X22Y157_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y157_SLICE_X22Y157_BO5),
.O6(CLBLM_L_X16Y157_SLICE_X22Y157_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y157_SLICE_X22Y157_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y157_SLICE_X22Y157_AO5),
.O6(CLBLM_L_X16Y157_SLICE_X22Y157_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y157_SLICE_X23Y157_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y157_SLICE_X23Y157_DO5),
.O6(CLBLM_L_X16Y157_SLICE_X23Y157_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y157_SLICE_X23Y157_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y157_SLICE_X23Y157_CO5),
.O6(CLBLM_L_X16Y157_SLICE_X23Y157_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y157_SLICE_X23Y157_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y157_SLICE_X23Y157_BO5),
.O6(CLBLM_L_X16Y157_SLICE_X23Y157_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y157_SLICE_X23Y157_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y157_SLICE_X23Y157_AO5),
.O6(CLBLM_L_X16Y157_SLICE_X23Y157_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X56Y151_SLICE_X84Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X1Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y136_SLICE_X13Y136_BO6),
.Q(CLBLM_L_X56Y151_SLICE_X84Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y151_SLICE_X84Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y151_SLICE_X84Y151_DO5),
.O6(CLBLM_L_X56Y151_SLICE_X84Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y151_SLICE_X84Y151_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y151_SLICE_X84Y151_CO5),
.O6(CLBLM_L_X56Y151_SLICE_X84Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y151_SLICE_X84Y151_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y151_SLICE_X84Y151_BO5),
.O6(CLBLM_L_X56Y151_SLICE_X84Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y151_SLICE_X84Y151_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y151_SLICE_X84Y151_AO5),
.O6(CLBLM_L_X56Y151_SLICE_X84Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y151_SLICE_X85Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y151_SLICE_X85Y151_DO5),
.O6(CLBLM_L_X56Y151_SLICE_X85Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y151_SLICE_X85Y151_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y151_SLICE_X85Y151_CO5),
.O6(CLBLM_L_X56Y151_SLICE_X85Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y151_SLICE_X85Y151_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y151_SLICE_X85Y151_BO5),
.O6(CLBLM_L_X56Y151_SLICE_X85Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y151_SLICE_X85Y151_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y151_SLICE_X85Y151_AO5),
.O6(CLBLM_L_X56Y151_SLICE_X85Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y129_SLICE_X2Y129_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y129_SLICE_X2Y129_AO5),
.Q(CLBLM_R_X3Y129_SLICE_X2Y129_A5Q),
.R(LIOB33_X0Y147_IOB_X0Y148_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y129_SLICE_X2Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y129_SLICE_X2Y129_AO6),
.Q(CLBLM_R_X3Y129_SLICE_X2Y129_AQ),
.R(LIOB33_X0Y147_IOB_X0Y148_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y129_SLICE_X2Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y129_SLICE_X2Y129_BO6),
.Q(CLBLM_R_X3Y129_SLICE_X2Y129_BQ),
.R(LIOB33_X0Y147_IOB_X0Y148_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y129_SLICE_X2Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y129_SLICE_X2Y129_DO5),
.O6(CLBLM_R_X3Y129_SLICE_X2Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y129_SLICE_X2Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y129_SLICE_X2Y129_CO5),
.O6(CLBLM_R_X3Y129_SLICE_X2Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333333333333)
  ) CLBLM_R_X3Y129_SLICE_X2Y129_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y129_SLICE_X2Y129_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y129_SLICE_X2Y129_BO5),
.O6(CLBLM_R_X3Y129_SLICE_X2Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3c3f3fc0c0)
  ) CLBLM_R_X3Y129_SLICE_X2Y129_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y129_SLICE_X2Y129_BQ),
.I2(CLBLM_R_X3Y129_SLICE_X2Y129_AQ),
.I3(1'b1),
.I4(CLBLM_R_X3Y129_SLICE_X2Y129_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y129_SLICE_X2Y129_AO5),
.O6(CLBLM_R_X3Y129_SLICE_X2Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y129_SLICE_X3Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y129_SLICE_X3Y129_DO5),
.O6(CLBLM_R_X3Y129_SLICE_X3Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y129_SLICE_X3Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y129_SLICE_X3Y129_CO5),
.O6(CLBLM_R_X3Y129_SLICE_X3Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y129_SLICE_X3Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y129_SLICE_X3Y129_BO5),
.O6(CLBLM_R_X3Y129_SLICE_X3Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y129_SLICE_X3Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y129_SLICE_X3Y129_AO5),
.O6(CLBLM_R_X3Y129_SLICE_X3Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y130_SLICE_X2Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y130_SLICE_X2Y130_AO6),
.Q(CLBLM_R_X3Y130_SLICE_X2Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y130_SLICE_X2Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y130_SLICE_X2Y130_DO5),
.O6(CLBLM_R_X3Y130_SLICE_X2Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y130_SLICE_X2Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y130_SLICE_X2Y130_CO5),
.O6(CLBLM_R_X3Y130_SLICE_X2Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y130_SLICE_X2Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y130_SLICE_X2Y130_BO5),
.O6(CLBLM_R_X3Y130_SLICE_X2Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff96ff9600960096)
  ) CLBLM_R_X3Y130_SLICE_X2Y130_ALUT (
.I0(CLBLM_R_X3Y131_SLICE_X2Y131_DO6),
.I1(CLBLM_R_X3Y131_SLICE_X3Y131_BQ),
.I2(CLBLM_R_X3Y130_SLICE_X2Y130_AQ),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(1'b1),
.I5(LIOB33_X0Y55_IOB_X0Y56_I),
.O5(CLBLM_R_X3Y130_SLICE_X2Y130_AO5),
.O6(CLBLM_R_X3Y130_SLICE_X2Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y130_SLICE_X3Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y130_SLICE_X3Y130_AO6),
.Q(CLBLM_R_X3Y130_SLICE_X3Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y130_SLICE_X3Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y130_SLICE_X3Y130_BO6),
.Q(CLBLM_R_X3Y130_SLICE_X3Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y130_SLICE_X3Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y130_SLICE_X3Y130_DO5),
.O6(CLBLM_R_X3Y130_SLICE_X3Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hde12ed21ed21de12)
  ) CLBLM_R_X3Y130_SLICE_X3Y130_CLUT (
.I0(CLBLM_R_X3Y130_SLICE_X2Y130_AQ),
.I1(LIOB33_X0Y147_IOB_X0Y148_I),
.I2(CLBLM_R_X3Y131_SLICE_X2Y131_DO6),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(CLBLM_R_X5Y130_SLICE_X7Y130_BQ),
.I5(CLBLM_R_X3Y131_SLICE_X3Y131_BQ),
.O5(CLBLM_R_X3Y130_SLICE_X3Y130_CO5),
.O6(CLBLM_R_X3Y130_SLICE_X3Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa3caac3aac3aa3c)
  ) CLBLM_R_X3Y130_SLICE_X3Y130_BLUT (
.I0(LIOB33_X0Y27_IOB_X0Y27_I),
.I1(CLBLM_R_X3Y130_SLICE_X3Y130_BQ),
.I2(CLBLM_R_X3Y130_SLICE_X3Y130_AQ),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(BRAM_L_X6Y125_RAMB18_X0Y50_DO21),
.I5(CLBLM_R_X7Y131_SLICE_X9Y131_A5Q),
.O5(CLBLM_R_X3Y130_SLICE_X3Y130_BO5),
.O6(CLBLM_R_X3Y130_SLICE_X3Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hedde21125a5a5a5a)
  ) CLBLM_R_X3Y130_SLICE_X3Y130_ALUT (
.I0(CLBLM_R_X7Y131_SLICE_X9Y131_A5Q),
.I1(LIOB33_X0Y147_IOB_X0Y148_I),
.I2(CLBLM_R_X3Y130_SLICE_X3Y130_AQ),
.I3(BRAM_L_X6Y125_RAMB18_X0Y50_DO21),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y130_SLICE_X3Y130_AO5),
.O6(CLBLM_R_X3Y130_SLICE_X3Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y131_SLICE_X2Y131_AO5),
.Q(CLBLM_R_X3Y131_SLICE_X2Y131_A5Q),
.R(LIOB33_X0Y147_IOB_X0Y148_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y131_SLICE_X2Y131_BO5),
.Q(CLBLM_R_X3Y131_SLICE_X2Y131_B5Q),
.R(LIOB33_X0Y147_IOB_X0Y148_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y131_SLICE_X2Y131_CO5),
.Q(CLBLM_R_X3Y131_SLICE_X2Y131_C5Q),
.R(LIOB33_X0Y147_IOB_X0Y148_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y131_SLICE_X2Y131_AO6),
.Q(CLBLM_R_X3Y131_SLICE_X2Y131_AQ),
.R(LIOB33_X0Y147_IOB_X0Y148_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y131_SLICE_X2Y131_BO6),
.Q(CLBLM_R_X3Y131_SLICE_X2Y131_BQ),
.R(LIOB33_X0Y147_IOB_X0Y148_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y131_SLICE_X2Y131_CO6),
.Q(CLBLM_R_X3Y131_SLICE_X2Y131_CQ),
.R(LIOB33_X0Y147_IOB_X0Y148_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha55aa55aedde2112)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_DLUT (
.I0(CLBLM_R_X3Y131_SLICE_X3Y131_AQ),
.I1(LIOB33_X0Y147_IOB_X0Y148_I),
.I2(BRAM_L_X6Y130_RAMB18_X0Y52_DO16),
.I3(CLBLL_L_X2Y131_SLICE_X1Y131_BQ),
.I4(LIOB33_X0Y139_IOB_X0Y140_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X2Y131_DO5),
.O6(CLBLM_R_X3Y131_SLICE_X2Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000440000002200)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_CLUT (
.I0(CLBLM_R_X3Y129_SLICE_X2Y129_AQ),
.I1(CLBLM_R_X3Y129_SLICE_X2Y129_BQ),
.I2(1'b1),
.I3(CLBLM_R_X3Y129_SLICE_X2Y129_A5Q),
.I4(CLBLL_L_X2Y131_SLICE_X1Y131_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X2Y131_CO5),
.O6(CLBLM_R_X3Y131_SLICE_X2Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0006000640104010)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_BLUT (
.I0(CLBLL_L_X2Y131_SLICE_X1Y131_A5Q),
.I1(CLBLM_R_X3Y129_SLICE_X2Y129_BQ),
.I2(CLBLM_R_X3Y129_SLICE_X2Y129_AQ),
.I3(CLBLM_R_X3Y129_SLICE_X2Y129_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X2Y131_BO5),
.O6(CLBLM_R_X3Y131_SLICE_X2Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3000000f3300000c)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y131_SLICE_X1Y131_A5Q),
.I2(CLBLM_R_X3Y129_SLICE_X2Y129_A5Q),
.I3(CLBLM_R_X3Y129_SLICE_X2Y129_BQ),
.I4(CLBLM_R_X3Y129_SLICE_X2Y129_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X2Y131_AO5),
.O6(CLBLM_R_X3Y131_SLICE_X2Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y131_SLICE_X3Y131_AO6),
.Q(CLBLM_R_X3Y131_SLICE_X3Y131_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y131_SLICE_X2Y131_DO5),
.Q(CLBLM_R_X3Y131_SLICE_X3Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y131_SLICE_X3Y131_BO6),
.Q(CLBLM_R_X3Y131_SLICE_X3Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y131_SLICE_X3Y131_CO6),
.Q(CLBLM_R_X3Y131_SLICE_X3Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y131_SLICE_X3Y131_DO6),
.Q(CLBLM_R_X3Y131_SLICE_X3Y131_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000069966996)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_DLUT (
.I0(CLBLM_R_X3Y132_SLICE_X3Y132_AQ),
.I1(CLBLM_R_X3Y131_SLICE_X2Y131_A5Q),
.I2(CLBLM_R_X3Y131_SLICE_X3Y131_DQ),
.I3(BRAM_L_X6Y130_RAMB18_X0Y52_DO20),
.I4(LIOB33_X0Y91_IOB_X0Y92_I),
.I5(LIOB33_X0Y147_IOB_X0Y148_I),
.O5(CLBLM_R_X3Y131_SLICE_X3Y131_DO5),
.O6(CLBLM_R_X3Y131_SLICE_X3Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf066f099f099f066)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_CLUT (
.I0(BRAM_L_X6Y130_RAMB18_X0Y52_DO18),
.I1(CLBLM_R_X3Y131_SLICE_X3Y131_CQ),
.I2(LIOB33_X0Y89_IOB_X0Y90_I),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(CLBLM_R_X3Y131_SLICE_X3Y131_B5Q),
.I5(CLBLM_R_X3Y131_SLICE_X2Y131_BQ),
.O5(CLBLM_R_X3Y131_SLICE_X3Y131_CO5),
.O6(CLBLM_R_X3Y131_SLICE_X3Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa3caac3aac3aa3c)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_BLUT (
.I0(LIOB33_X0Y87_IOB_X0Y88_I),
.I1(CLBLM_R_X3Y131_SLICE_X3Y131_BQ),
.I2(CLBLM_R_X3Y131_SLICE_X3Y131_AQ),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(BRAM_L_X6Y130_RAMB18_X0Y52_DO16),
.I5(CLBLL_L_X2Y131_SLICE_X1Y131_BQ),
.O5(CLBLM_R_X3Y131_SLICE_X3Y131_BO5),
.O6(CLBLM_R_X3Y131_SLICE_X3Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0996699669966)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_ALUT (
.I0(CLBLM_R_X3Y131_SLICE_X3Y131_B5Q),
.I1(BRAM_L_X6Y130_RAMB18_X0Y52_DO18),
.I2(LIOB33_X0Y141_IOB_X0Y142_I),
.I3(CLBLM_R_X3Y131_SLICE_X2Y131_BQ),
.I4(LIOB33_X0Y147_IOB_X0Y148_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X3Y131_AO5),
.O6(CLBLM_R_X3Y131_SLICE_X3Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y132_SLICE_X2Y132_AO6),
.Q(CLBLM_R_X3Y132_SLICE_X2Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y132_SLICE_X2Y132_BO6),
.Q(CLBLM_R_X3Y132_SLICE_X2Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y132_SLICE_X2Y132_CO6),
.Q(CLBLM_R_X3Y132_SLICE_X2Y132_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y132_SLICE_X2Y132_DO6),
.Q(CLBLM_R_X3Y132_SLICE_X2Y132_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000069966996)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_DLUT (
.I0(CLBLM_R_X3Y132_SLICE_X2Y132_BQ),
.I1(CLBLM_R_X3Y131_SLICE_X2Y131_C5Q),
.I2(CLBLM_R_X3Y132_SLICE_X2Y132_DQ),
.I3(BRAM_L_X6Y130_RAMB18_X0Y52_DO23),
.I4(LIOB33_X0Y95_IOB_X0Y95_I),
.I5(LIOB33_X0Y147_IOB_X0Y148_I),
.O5(CLBLM_R_X3Y132_SLICE_X2Y132_DO5),
.O6(CLBLM_R_X3Y132_SLICE_X2Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000069966996)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_CLUT (
.I0(CLBLM_R_X3Y132_SLICE_X2Y132_AQ),
.I1(CLBLM_R_X3Y132_SLICE_X2Y132_CQ),
.I2(BRAM_L_X6Y130_RAMB18_X0Y52_DO22),
.I3(CLBLM_R_X3Y131_SLICE_X2Y131_CQ),
.I4(LIOB33_X0Y93_IOB_X0Y94_I),
.I5(LIOB33_X0Y147_IOB_X0Y148_I),
.O5(CLBLM_R_X3Y132_SLICE_X2Y132_CO5),
.O6(CLBLM_R_X3Y132_SLICE_X2Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb88b8bb8f00f0ff0)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_BLUT (
.I0(LIOB33_X0Y147_IOB_X0Y147_I),
.I1(LIOB33_X0Y147_IOB_X0Y148_I),
.I2(CLBLM_R_X3Y131_SLICE_X2Y131_C5Q),
.I3(BRAM_L_X6Y130_RAMB18_X0Y52_DO23),
.I4(CLBLM_R_X3Y132_SLICE_X2Y132_BQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y132_SLICE_X2Y132_BO5),
.O6(CLBLM_R_X3Y132_SLICE_X2Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hed21de12a5a55a5a)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_ALUT (
.I0(BRAM_L_X6Y130_RAMB18_X0Y52_DO22),
.I1(LIOB33_X0Y147_IOB_X0Y148_I),
.I2(CLBLM_R_X3Y132_SLICE_X2Y132_AQ),
.I3(LIOB33_X0Y145_IOB_X0Y146_I),
.I4(CLBLM_R_X3Y131_SLICE_X2Y131_CQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y132_SLICE_X2Y132_AO5),
.O6(CLBLM_R_X3Y132_SLICE_X2Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y132_SLICE_X3Y132_AO6),
.Q(CLBLM_R_X3Y132_SLICE_X3Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y132_SLICE_X3Y132_BO6),
.Q(CLBLM_R_X3Y132_SLICE_X3Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y132_SLICE_X3Y132_CO6),
.Q(CLBLM_R_X3Y132_SLICE_X3Y132_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y132_SLICE_X3Y132_DO5),
.O6(CLBLM_R_X3Y132_SLICE_X3Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000096969696)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_CLUT (
.I0(CLBLM_R_X3Y132_SLICE_X2Y132_DQ),
.I1(CLBLM_R_X3Y132_SLICE_X3Y132_CQ),
.I2(CLBLM_R_X3Y132_SLICE_X2Y132_BO5),
.I3(1'b1),
.I4(LIOB33_X0Y63_IOB_X0Y63_I),
.I5(LIOB33_X0Y147_IOB_X0Y148_I),
.O5(CLBLM_R_X3Y132_SLICE_X3Y132_CO5),
.O6(CLBLM_R_X3Y132_SLICE_X3Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa3caac3aac3aa3c)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_BLUT (
.I0(LIOB33_X0Y93_IOB_X0Y93_I),
.I1(CLBLM_R_X3Y132_SLICE_X3Y132_BQ),
.I2(CLBLL_L_X2Y131_SLICE_X1Y131_AQ),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(CLBLM_R_X3Y133_SLICE_X3Y133_AQ),
.I5(BRAM_L_X6Y130_RAMB18_X0Y52_DO21),
.O5(CLBLM_R_X3Y132_SLICE_X3Y132_BO5),
.O6(CLBLM_R_X3Y132_SLICE_X3Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haac3aa3cc3c33c3c)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_ALUT (
.I0(1'b1),
.I1(BRAM_L_X6Y130_RAMB18_X0Y52_DO20),
.I2(CLBLM_R_X3Y132_SLICE_X3Y132_AQ),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(CLBLM_R_X3Y131_SLICE_X2Y131_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y132_SLICE_X3Y132_AO5),
.O6(CLBLM_R_X3Y132_SLICE_X3Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y133_SLICE_X2Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y133_SLICE_X2Y133_DO5),
.O6(CLBLM_R_X3Y133_SLICE_X2Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y133_SLICE_X2Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y133_SLICE_X2Y133_CO5),
.O6(CLBLM_R_X3Y133_SLICE_X2Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y133_SLICE_X2Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y133_SLICE_X2Y133_BO5),
.O6(CLBLM_R_X3Y133_SLICE_X2Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y133_SLICE_X2Y133_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y133_SLICE_X2Y133_AO5),
.O6(CLBLM_R_X3Y133_SLICE_X2Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y133_SLICE_X3Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y133_SLICE_X3Y133_AO6),
.Q(CLBLM_R_X3Y133_SLICE_X3Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y133_SLICE_X3Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y133_SLICE_X3Y133_BO6),
.Q(CLBLM_R_X3Y133_SLICE_X3Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y133_SLICE_X3Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y133_SLICE_X3Y133_DO5),
.O6(CLBLM_R_X3Y133_SLICE_X3Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y133_SLICE_X3Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y133_SLICE_X3Y133_CO5),
.O6(CLBLM_R_X3Y133_SLICE_X3Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff99ff6600990066)
  ) CLBLM_R_X3Y133_SLICE_X3Y133_BLUT (
.I0(CLBLM_R_X3Y131_SLICE_X3Y131_DQ),
.I1(CLBLM_R_X3Y133_SLICE_X3Y133_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(CLBLM_R_X3Y132_SLICE_X3Y132_AO5),
.I5(LIOB33_X0Y59_IOB_X0Y60_I),
.O5(CLBLM_R_X3Y133_SLICE_X3Y133_BO5),
.O6(CLBLM_R_X3Y133_SLICE_X3Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haac3aa3cc3c33c3c)
  ) CLBLM_R_X3Y133_SLICE_X3Y133_ALUT (
.I0(LIOB33_X0Y145_IOB_X0Y145_I),
.I1(BRAM_L_X6Y130_RAMB18_X0Y52_DO21),
.I2(CLBLM_R_X3Y133_SLICE_X3Y133_AQ),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(CLBLL_L_X2Y131_SLICE_X1Y131_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y133_SLICE_X3Y133_AO5),
.O6(CLBLM_R_X3Y133_SLICE_X3Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y134_SLICE_X2Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y134_SLICE_X2Y134_AO6),
.Q(CLBLM_R_X3Y134_SLICE_X2Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y134_SLICE_X2Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y134_SLICE_X2Y134_BO6),
.Q(CLBLM_R_X3Y134_SLICE_X2Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y134_SLICE_X2Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y134_SLICE_X2Y134_DO5),
.O6(CLBLM_R_X3Y134_SLICE_X2Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y134_SLICE_X2Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y134_SLICE_X2Y134_CO5),
.O6(CLBLM_R_X3Y134_SLICE_X2Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff69ff9600690096)
  ) CLBLM_R_X3Y134_SLICE_X2Y134_BLUT (
.I0(CLBLM_R_X5Y134_SLICE_X7Y134_A5Q),
.I1(CLBLM_R_X3Y134_SLICE_X2Y134_BQ),
.I2(CLBLM_R_X3Y134_SLICE_X2Y134_AQ),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(BRAM_L_X6Y125_RAMB18_X0Y50_DO23),
.I5(LIOB33_X0Y29_IOB_X0Y29_I),
.O5(CLBLM_R_X3Y134_SLICE_X2Y134_BO5),
.O6(CLBLM_R_X3Y134_SLICE_X2Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haac3aa3c3c3c3c3c)
  ) CLBLM_R_X3Y134_SLICE_X2Y134_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_R_X5Y134_SLICE_X7Y134_A5Q),
.I2(CLBLM_R_X3Y134_SLICE_X2Y134_AQ),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(BRAM_L_X6Y125_RAMB18_X0Y50_DO23),
.I5(1'b1),
.O5(CLBLM_R_X3Y134_SLICE_X2Y134_AO5),
.O6(CLBLM_R_X3Y134_SLICE_X2Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y134_SLICE_X3Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y134_SLICE_X3Y134_DO5),
.O6(CLBLM_R_X3Y134_SLICE_X3Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y134_SLICE_X3Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y134_SLICE_X3Y134_CO5),
.O6(CLBLM_R_X3Y134_SLICE_X3Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y134_SLICE_X3Y134_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y134_SLICE_X3Y134_BO5),
.O6(CLBLM_R_X3Y134_SLICE_X3Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa3cc3c33c)
  ) CLBLM_R_X3Y134_SLICE_X3Y134_ALUT (
.I0(LIOB33_X0Y13_IOB_X0Y14_I),
.I1(CLBLL_L_X4Y134_SLICE_X4Y134_AQ),
.I2(CLBLM_R_X3Y134_SLICE_X2Y134_AO5),
.I3(CLBLM_R_X3Y134_SLICE_X2Y134_BQ),
.I4(BRAM_L_X6Y125_RAMB18_X0Y50_DO23),
.I5(LIOB33_X0Y147_IOB_X0Y148_I),
.O5(CLBLM_R_X3Y134_SLICE_X3Y134_AO5),
.O6(CLBLM_R_X3Y134_SLICE_X3Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y135_SLICE_X2Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y135_SLICE_X2Y135_DO5),
.O6(CLBLM_R_X3Y135_SLICE_X2Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y135_SLICE_X2Y135_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y135_SLICE_X2Y135_CO5),
.O6(CLBLM_R_X3Y135_SLICE_X2Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y135_SLICE_X2Y135_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y135_SLICE_X2Y135_BO5),
.O6(CLBLM_R_X3Y135_SLICE_X2Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y135_SLICE_X2Y135_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y135_SLICE_X2Y135_AO5),
.O6(CLBLM_R_X3Y135_SLICE_X2Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa55aaf0f0f0f0)
  ) CLBLM_R_X3Y135_SLICE_X3Y135_DLUT (
.I0(CLBLM_R_X5Y130_SLICE_X6Y130_B5Q),
.I1(1'b1),
.I2(CLBLM_R_X5Y135_SLICE_X6Y135_DO6),
.I3(CLBLM_R_X3Y147_SLICE_X3Y147_CQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.O5(CLBLM_R_X3Y135_SLICE_X3Y135_DO5),
.O6(CLBLM_R_X3Y135_SLICE_X3Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h77bb448877bb4488)
  ) CLBLM_R_X3Y135_SLICE_X3Y135_CLUT (
.I0(CLBLM_R_X3Y134_SLICE_X2Y134_AQ),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I2(1'b1),
.I3(CLBLL_L_X2Y158_SLICE_X0Y158_CQ),
.I4(CLBLM_R_X5Y135_SLICE_X6Y135_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y135_SLICE_X3Y135_CO5),
.O6(CLBLM_R_X3Y135_SLICE_X3Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fcc0fccf0ccf0cc)
  ) CLBLM_R_X3Y135_SLICE_X3Y135_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y135_SLICE_X7Y135_BO6),
.I2(CLBLL_L_X2Y158_SLICE_X0Y158_BQ),
.I3(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y131_SLICE_X5Y131_B5Q),
.O5(CLBLM_R_X3Y135_SLICE_X3Y135_BO5),
.O6(CLBLM_R_X3Y135_SLICE_X3Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h22ee22eeee22ee22)
  ) CLBLM_R_X3Y135_SLICE_X3Y135_ALUT (
.I0(CLBLM_R_X5Y135_SLICE_X6Y135_BO6),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y132_SLICE_X7Y132_A5Q),
.I4(1'b1),
.I5(CLBLM_R_X3Y147_SLICE_X2Y147_CQ),
.O5(CLBLM_R_X3Y135_SLICE_X3Y135_AO5),
.O6(CLBLM_R_X3Y135_SLICE_X3Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aff5aff5a005a00)
  ) CLBLM_R_X3Y137_SLICE_X2Y137_DLUT (
.I0(CLBLM_R_X3Y134_SLICE_X2Y134_BQ),
.I1(1'b1),
.I2(CLBLL_L_X2Y155_SLICE_X1Y155_BQ),
.I3(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y137_SLICE_X2Y137_BO6),
.O5(CLBLM_R_X3Y137_SLICE_X2Y137_DO5),
.O6(CLBLM_R_X3Y137_SLICE_X2Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cc33ccf0f0f0f0)
  ) CLBLM_R_X3Y137_SLICE_X2Y137_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y155_SLICE_X0Y155_BQ),
.I2(CLBLL_L_X4Y137_SLICE_X4Y137_BO6),
.I3(CLBLL_L_X4Y131_SLICE_X4Y131_DQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.O5(CLBLM_R_X3Y137_SLICE_X2Y137_CO5),
.O6(CLBLM_R_X3Y137_SLICE_X2Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X3Y137_SLICE_X2Y137_BLUT (
.I0(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO7),
.I1(BRAM_L_X6Y140_RAMB18_X0Y56_DO7),
.I2(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO6),
.I3(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO7),
.I4(CLBLM_R_X3Y134_SLICE_X2Y134_BQ),
.I5(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO6),
.O5(CLBLM_R_X3Y137_SLICE_X2Y137_BO5),
.O6(CLBLM_R_X3Y137_SLICE_X2Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X3Y137_SLICE_X2Y137_ALUT (
.I0(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO7),
.I1(CLBLM_R_X3Y130_SLICE_X2Y130_AQ),
.I2(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO0),
.I3(BRAM_L_X6Y140_RAMB18_X0Y56_DO7),
.I4(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO0),
.I5(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO0),
.O5(CLBLM_R_X3Y137_SLICE_X2Y137_AO5),
.O6(CLBLM_R_X3Y137_SLICE_X2Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h77bb77bb44884488)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_DLUT (
.I0(CLBLM_R_X3Y157_SLICE_X3Y157_AQ),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y133_SLICE_X5Y133_BQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y137_SLICE_X3Y137_BO6),
.O5(CLBLM_R_X3Y137_SLICE_X3Y137_DO5),
.O6(CLBLM_R_X3Y137_SLICE_X3Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_CLUT (
.I0(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO6),
.I1(BRAM_L_X6Y140_RAMB18_X0Y56_DO7),
.I2(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO7),
.I3(BRAM_L_X6Y140_RAMB18_X0Y56_DO6),
.I4(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO7),
.I5(CLBLL_L_X4Y128_SLICE_X5Y128_BQ),
.O5(CLBLM_R_X3Y137_SLICE_X3Y137_CO5),
.O6(CLBLM_R_X3Y137_SLICE_X3Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_BLUT (
.I0(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO7),
.I1(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO6),
.I2(CLBLL_L_X4Y133_SLICE_X5Y133_BQ),
.I3(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO7),
.I4(BRAM_L_X6Y140_RAMB18_X0Y56_DO7),
.I5(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO6),
.O5(CLBLM_R_X3Y137_SLICE_X3Y137_BO5),
.O6(CLBLM_R_X3Y137_SLICE_X3Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cc33cc0ff00ff0)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_ALUT (
.I0(1'b1),
.I1(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO7),
.I2(CLBLM_R_X3Y134_SLICE_X2Y134_BQ),
.I3(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO7),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y137_SLICE_X3Y137_AO5),
.O6(CLBLM_R_X3Y137_SLICE_X3Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y138_SLICE_X2Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y138_SLICE_X2Y138_DO5),
.O6(CLBLM_R_X3Y138_SLICE_X2Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y138_SLICE_X2Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y138_SLICE_X2Y138_CO5),
.O6(CLBLM_R_X3Y138_SLICE_X2Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y138_SLICE_X2Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y138_SLICE_X2Y138_BO5),
.O6(CLBLM_R_X3Y138_SLICE_X2Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff00f0ff0ff000)
  ) CLBLM_R_X3Y138_SLICE_X2Y138_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I3(CLBLL_L_X2Y132_SLICE_X1Y132_AQ),
.I4(CLBLL_L_X4Y136_SLICE_X4Y136_AO6),
.I5(CLBLL_L_X2Y157_SLICE_X0Y157_CQ),
.O5(CLBLM_R_X3Y138_SLICE_X2Y138_AO5),
.O6(CLBLM_R_X3Y138_SLICE_X2Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7d287d287d287d28)
  ) CLBLM_R_X3Y138_SLICE_X3Y138_DLUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I1(CLBLL_L_X4Y128_SLICE_X5Y128_BQ),
.I2(CLBLM_R_X3Y153_SLICE_X3Y153_DQ),
.I3(CLBLM_R_X3Y137_SLICE_X3Y137_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y138_SLICE_X3Y138_DO5),
.O6(CLBLM_R_X3Y138_SLICE_X3Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4e1b1b4ee4b1b1e4)
  ) CLBLM_R_X3Y138_SLICE_X3Y138_CLUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I1(BRAM_L_X6Y140_RAMB18_X0Y56_DO7),
.I2(CLBLM_R_X3Y151_SLICE_X2Y151_CQ),
.I3(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO7),
.I4(CLBLL_L_X4Y137_SLICE_X4Y137_DO6),
.I5(CLBLM_R_X5Y125_SLICE_X7Y125_CQ),
.O5(CLBLM_R_X3Y138_SLICE_X3Y138_CO5),
.O6(CLBLM_R_X3Y138_SLICE_X3Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff099990ff06666)
  ) CLBLM_R_X3Y138_SLICE_X3Y138_BLUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y56_DO7),
.I1(CLBLL_L_X4Y138_SLICE_X4Y138_CO6),
.I2(CLBLM_R_X5Y126_SLICE_X6Y126_BQ),
.I3(CLBLM_R_X3Y153_SLICE_X3Y153_AQ),
.I4(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I5(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO7),
.O5(CLBLM_R_X3Y138_SLICE_X3Y138_BO5),
.O6(CLBLM_R_X3Y138_SLICE_X3Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33a5cca5335acc5a)
  ) CLBLM_R_X3Y138_SLICE_X3Y138_ALUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y56_DO7),
.I1(CLBLM_R_X3Y133_SLICE_X3Y133_BQ),
.I2(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO7),
.I3(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I4(CLBLL_L_X2Y157_SLICE_X0Y157_AQ),
.I5(CLBLL_L_X4Y138_SLICE_X5Y138_BO6),
.O5(CLBLM_R_X3Y138_SLICE_X3Y138_AO5),
.O6(CLBLM_R_X3Y138_SLICE_X3Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y139_SLICE_X2Y139_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y139_SLICE_X2Y139_DO5),
.O6(CLBLM_R_X3Y139_SLICE_X2Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y139_SLICE_X2Y139_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y139_SLICE_X2Y139_CO5),
.O6(CLBLM_R_X3Y139_SLICE_X2Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y139_SLICE_X2Y139_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y139_SLICE_X2Y139_BO5),
.O6(CLBLM_R_X3Y139_SLICE_X2Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ccf0f033ccf0f0)
  ) CLBLM_R_X3Y139_SLICE_X2Y139_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y130_SLICE_X2Y130_AQ),
.I2(CLBLM_R_X3Y137_SLICE_X2Y137_AO6),
.I3(CLBLM_R_X3Y157_SLICE_X3Y157_BQ),
.I4(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y139_SLICE_X2Y139_AO5),
.O6(CLBLM_R_X3Y139_SLICE_X2Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y139_SLICE_X3Y139_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y139_SLICE_X3Y139_DO5),
.O6(CLBLM_R_X3Y139_SLICE_X3Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y139_SLICE_X3Y139_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y139_SLICE_X3Y139_CO5),
.O6(CLBLM_R_X3Y139_SLICE_X3Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y139_SLICE_X3Y139_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y139_SLICE_X3Y139_BO5),
.O6(CLBLM_R_X3Y139_SLICE_X3Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y139_SLICE_X3Y139_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y139_SLICE_X3Y139_AO5),
.O6(CLBLM_R_X3Y139_SLICE_X3Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y141_SLICE_X2Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.Q(CLBLM_R_X3Y141_SLICE_X2Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y141_SLICE_X2Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y159_IOB_X0Y160_I),
.Q(CLBLM_R_X3Y141_SLICE_X2Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y141_SLICE_X2Y141_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y157_IOB_X0Y158_I),
.Q(CLBLM_R_X3Y141_SLICE_X2Y141_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y141_SLICE_X2Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y141_SLICE_X2Y141_DO5),
.O6(CLBLM_R_X3Y141_SLICE_X2Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y141_SLICE_X2Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y141_SLICE_X2Y141_CO5),
.O6(CLBLM_R_X3Y141_SLICE_X2Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y141_SLICE_X2Y141_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y141_SLICE_X2Y141_BO5),
.O6(CLBLM_R_X3Y141_SLICE_X2Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y141_SLICE_X2Y141_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y141_SLICE_X2Y141_AO5),
.O6(CLBLM_R_X3Y141_SLICE_X2Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y141_SLICE_X3Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y141_SLICE_X3Y141_DO5),
.O6(CLBLM_R_X3Y141_SLICE_X3Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y141_SLICE_X3Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y141_SLICE_X3Y141_CO5),
.O6(CLBLM_R_X3Y141_SLICE_X3Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y141_SLICE_X3Y141_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y141_SLICE_X3Y141_BO5),
.O6(CLBLM_R_X3Y141_SLICE_X3Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y141_SLICE_X3Y141_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y141_SLICE_X3Y141_AO5),
.O6(CLBLM_R_X3Y141_SLICE_X3Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y161_IOB_X0Y161_I),
.Q(CLBLM_R_X3Y142_SLICE_X2Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y151_IOB_X0Y151_I),
.Q(CLBLM_R_X3Y142_SLICE_X2Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y153_IOB_X0Y153_I),
.Q(CLBLM_R_X3Y142_SLICE_X2Y142_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y159_IOB_X0Y159_I),
.Q(CLBLM_R_X3Y142_SLICE_X2Y142_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y142_SLICE_X2Y142_DO5),
.O6(CLBLM_R_X3Y142_SLICE_X2Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y142_SLICE_X2Y142_CO5),
.O6(CLBLM_R_X3Y142_SLICE_X2Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y142_SLICE_X2Y142_BO5),
.O6(CLBLM_R_X3Y142_SLICE_X2Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y142_SLICE_X2Y142_AO5),
.O6(CLBLM_R_X3Y142_SLICE_X2Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y142_SLICE_X3Y142_DO5),
.O6(CLBLM_R_X3Y142_SLICE_X3Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y142_SLICE_X3Y142_CO5),
.O6(CLBLM_R_X3Y142_SLICE_X3Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y142_SLICE_X3Y142_BO5),
.O6(CLBLM_R_X3Y142_SLICE_X3Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y142_SLICE_X3Y142_AO5),
.O6(CLBLM_R_X3Y142_SLICE_X3Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y153_IOB_X0Y154_I),
.Q(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y155_IOB_X0Y155_I),
.Q(CLBLM_R_X3Y145_SLICE_X2Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y155_IOB_X0Y156_I),
.Q(CLBLM_R_X3Y145_SLICE_X2Y145_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y157_IOB_X0Y157_I),
.Q(CLBLM_R_X3Y145_SLICE_X2Y145_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y145_SLICE_X2Y145_DO5),
.O6(CLBLM_R_X3Y145_SLICE_X2Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y145_SLICE_X2Y145_CO5),
.O6(CLBLM_R_X3Y145_SLICE_X2Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y145_SLICE_X2Y145_BO5),
.O6(CLBLM_R_X3Y145_SLICE_X2Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y145_SLICE_X2Y145_AO5),
.O6(CLBLM_R_X3Y145_SLICE_X2Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y165_IOB_X0Y165_I),
.Q(CLBLM_R_X3Y145_SLICE_X3Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y151_IOB_X0Y152_I),
.Q(CLBLM_R_X3Y145_SLICE_X3Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y145_SLICE_X3Y145_DO5),
.O6(CLBLM_R_X3Y145_SLICE_X3Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y145_SLICE_X3Y145_CO5),
.O6(CLBLM_R_X3Y145_SLICE_X3Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y145_SLICE_X3Y145_BO5),
.O6(CLBLM_R_X3Y145_SLICE_X3Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y145_SLICE_X3Y145_AO5),
.O6(CLBLM_R_X3Y145_SLICE_X3Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y169_IOB_X0Y170_I),
.Q(CLBLM_R_X3Y147_SLICE_X2Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y171_IOB_X0Y171_I),
.Q(CLBLM_R_X3Y147_SLICE_X2Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y171_IOB_X0Y172_I),
.Q(CLBLM_R_X3Y147_SLICE_X2Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y173_IOB_X0Y173_I),
.Q(CLBLM_R_X3Y147_SLICE_X2Y147_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y147_SLICE_X2Y147_DO5),
.O6(CLBLM_R_X3Y147_SLICE_X2Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y147_SLICE_X2Y147_CO5),
.O6(CLBLM_R_X3Y147_SLICE_X2Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y147_SLICE_X2Y147_BO5),
.O6(CLBLM_R_X3Y147_SLICE_X2Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y147_SLICE_X2Y147_AO5),
.O6(CLBLM_R_X3Y147_SLICE_X2Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y161_IOB_X0Y162_I),
.Q(CLBLM_R_X3Y147_SLICE_X3Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y163_IOB_X0Y163_I),
.Q(CLBLM_R_X3Y147_SLICE_X3Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y163_IOB_X0Y164_I),
.Q(CLBLM_R_X3Y147_SLICE_X3Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y167_IOB_X0Y168_I),
.Q(CLBLM_R_X3Y147_SLICE_X3Y147_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y147_SLICE_X3Y147_DO5),
.O6(CLBLM_R_X3Y147_SLICE_X3Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y147_SLICE_X3Y147_CO5),
.O6(CLBLM_R_X3Y147_SLICE_X3Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y147_SLICE_X3Y147_BO5),
.O6(CLBLM_R_X3Y147_SLICE_X3Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y147_SLICE_X3Y147_AO5),
.O6(CLBLM_R_X3Y147_SLICE_X3Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y175_IOB_X0Y175_I),
.Q(CLBLM_R_X3Y149_SLICE_X2Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y175_IOB_X0Y176_I),
.Q(CLBLM_R_X3Y149_SLICE_X2Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y177_IOB_X0Y177_I),
.Q(CLBLM_R_X3Y149_SLICE_X2Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y177_IOB_X0Y178_I),
.Q(CLBLM_R_X3Y149_SLICE_X2Y149_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y149_SLICE_X2Y149_DO5),
.O6(CLBLM_R_X3Y149_SLICE_X2Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y149_SLICE_X2Y149_CO5),
.O6(CLBLM_R_X3Y149_SLICE_X2Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y149_SLICE_X2Y149_BO5),
.O6(CLBLM_R_X3Y149_SLICE_X2Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y149_SLICE_X2Y149_AO5),
.O6(CLBLM_R_X3Y149_SLICE_X2Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y173_IOB_X0Y174_I),
.Q(CLBLM_R_X3Y149_SLICE_X3Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y149_SLICE_X3Y149_DO5),
.O6(CLBLM_R_X3Y149_SLICE_X3Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y149_SLICE_X3Y149_CO5),
.O6(CLBLM_R_X3Y149_SLICE_X3Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y149_SLICE_X3Y149_BO5),
.O6(CLBLM_R_X3Y149_SLICE_X3Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y149_SLICE_X3Y149_AO5),
.O6(CLBLM_R_X3Y149_SLICE_X3Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y151_SLICE_X2Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y181_IOB_X0Y181_I),
.Q(CLBLM_R_X3Y151_SLICE_X2Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y151_SLICE_X2Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y181_IOB_X0Y182_I),
.Q(CLBLM_R_X3Y151_SLICE_X2Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y151_SLICE_X2Y151_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y183_IOB_X0Y183_I),
.Q(CLBLM_R_X3Y151_SLICE_X2Y151_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y151_SLICE_X2Y151_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y183_IOB_X0Y184_I),
.Q(CLBLM_R_X3Y151_SLICE_X2Y151_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y151_SLICE_X2Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y151_SLICE_X2Y151_DO5),
.O6(CLBLM_R_X3Y151_SLICE_X2Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y151_SLICE_X2Y151_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y151_SLICE_X2Y151_CO5),
.O6(CLBLM_R_X3Y151_SLICE_X2Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y151_SLICE_X2Y151_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y151_SLICE_X2Y151_BO5),
.O6(CLBLM_R_X3Y151_SLICE_X2Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y151_SLICE_X2Y151_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y151_SLICE_X2Y151_AO5),
.O6(CLBLM_R_X3Y151_SLICE_X2Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y151_SLICE_X3Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y179_IOB_X0Y179_I),
.Q(CLBLM_R_X3Y151_SLICE_X3Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y151_SLICE_X3Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y179_IOB_X0Y180_I),
.Q(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y151_SLICE_X3Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y151_SLICE_X3Y151_DO5),
.O6(CLBLM_R_X3Y151_SLICE_X3Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y151_SLICE_X3Y151_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y151_SLICE_X3Y151_CO5),
.O6(CLBLM_R_X3Y151_SLICE_X3Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y151_SLICE_X3Y151_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y151_SLICE_X3Y151_BO5),
.O6(CLBLM_R_X3Y151_SLICE_X3Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y151_SLICE_X3Y151_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y151_SLICE_X3Y151_AO5),
.O6(CLBLM_R_X3Y151_SLICE_X3Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y153_SLICE_X2Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y189_IOB_X0Y190_I),
.Q(CLBLM_R_X3Y153_SLICE_X2Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y153_SLICE_X2Y153_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y191_IOB_X0Y191_I),
.Q(CLBLM_R_X3Y153_SLICE_X2Y153_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y153_SLICE_X2Y153_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y191_IOB_X0Y192_I),
.Q(CLBLM_R_X3Y153_SLICE_X2Y153_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y153_SLICE_X2Y153_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y193_IOB_X0Y193_I),
.Q(CLBLM_R_X3Y153_SLICE_X2Y153_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y153_SLICE_X2Y153_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y153_SLICE_X2Y153_DO5),
.O6(CLBLM_R_X3Y153_SLICE_X2Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y153_SLICE_X2Y153_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y153_SLICE_X2Y153_CO5),
.O6(CLBLM_R_X3Y153_SLICE_X2Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y153_SLICE_X2Y153_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y153_SLICE_X2Y153_BO5),
.O6(CLBLM_R_X3Y153_SLICE_X2Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y153_SLICE_X2Y153_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y153_SLICE_X2Y153_AO5),
.O6(CLBLM_R_X3Y153_SLICE_X2Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y153_SLICE_X3Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y185_IOB_X0Y185_I),
.Q(CLBLM_R_X3Y153_SLICE_X3Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y153_SLICE_X3Y153_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y185_IOB_X0Y186_I),
.Q(CLBLM_R_X3Y153_SLICE_X3Y153_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y153_SLICE_X3Y153_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y187_IOB_X0Y188_I),
.Q(CLBLM_R_X3Y153_SLICE_X3Y153_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y153_SLICE_X3Y153_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y189_IOB_X0Y189_I),
.Q(CLBLM_R_X3Y153_SLICE_X3Y153_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y153_SLICE_X3Y153_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y153_SLICE_X3Y153_DO5),
.O6(CLBLM_R_X3Y153_SLICE_X3Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y153_SLICE_X3Y153_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y153_SLICE_X3Y153_CO5),
.O6(CLBLM_R_X3Y153_SLICE_X3Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y153_SLICE_X3Y153_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y153_SLICE_X3Y153_BO5),
.O6(CLBLM_R_X3Y153_SLICE_X3Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y153_SLICE_X3Y153_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y153_SLICE_X3Y153_AO5),
.O6(CLBLM_R_X3Y153_SLICE_X3Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y155_SLICE_X2Y155_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y221_IOB_X0Y222_I),
.Q(CLBLM_R_X3Y155_SLICE_X2Y155_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y155_SLICE_X2Y155_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y225_IOB_X0Y225_I),
.Q(CLBLM_R_X3Y155_SLICE_X2Y155_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y155_SLICE_X2Y155_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y231_IOB_X0Y231_I),
.Q(CLBLM_R_X3Y155_SLICE_X2Y155_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y155_SLICE_X2Y155_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y239_IOB_X0Y240_I),
.Q(CLBLM_R_X3Y155_SLICE_X2Y155_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y155_SLICE_X2Y155_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y155_SLICE_X2Y155_DO5),
.O6(CLBLM_R_X3Y155_SLICE_X2Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y155_SLICE_X2Y155_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y155_SLICE_X2Y155_CO5),
.O6(CLBLM_R_X3Y155_SLICE_X2Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y155_SLICE_X2Y155_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y155_SLICE_X2Y155_BO5),
.O6(CLBLM_R_X3Y155_SLICE_X2Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y155_SLICE_X2Y155_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y155_SLICE_X2Y155_AO5),
.O6(CLBLM_R_X3Y155_SLICE_X2Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y155_SLICE_X3Y155_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y195_IOB_X0Y196_I),
.Q(CLBLM_R_X3Y155_SLICE_X3Y155_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y155_SLICE_X3Y155_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y197_IOB_X0Y198_I),
.Q(CLBLM_R_X3Y155_SLICE_X3Y155_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y155_SLICE_X3Y155_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y201_IOB_X0Y202_I),
.Q(CLBLM_R_X3Y155_SLICE_X3Y155_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y155_SLICE_X3Y155_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y155_SLICE_X3Y155_DO5),
.O6(CLBLM_R_X3Y155_SLICE_X3Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y155_SLICE_X3Y155_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y155_SLICE_X3Y155_CO5),
.O6(CLBLM_R_X3Y155_SLICE_X3Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y155_SLICE_X3Y155_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y155_SLICE_X3Y155_BO5),
.O6(CLBLM_R_X3Y155_SLICE_X3Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y155_SLICE_X3Y155_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y155_SLICE_X3Y155_AO5),
.O6(CLBLM_R_X3Y155_SLICE_X3Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y157_SLICE_X2Y157_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y227_IOB_X0Y227_I),
.Q(CLBLM_R_X3Y157_SLICE_X2Y157_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y157_SLICE_X2Y157_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y243_IOB_X0Y243_I),
.Q(CLBLM_R_X3Y157_SLICE_X2Y157_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y157_SLICE_X2Y157_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y247_IOB_X0Y248_I),
.Q(CLBLM_R_X3Y157_SLICE_X2Y157_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y157_SLICE_X2Y157_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_SING_X0Y249_IOB_X0Y249_I),
.Q(CLBLM_R_X3Y157_SLICE_X2Y157_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y157_SLICE_X2Y157_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y157_SLICE_X2Y157_DO5),
.O6(CLBLM_R_X3Y157_SLICE_X2Y157_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y157_SLICE_X2Y157_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y157_SLICE_X2Y157_CO5),
.O6(CLBLM_R_X3Y157_SLICE_X2Y157_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y157_SLICE_X2Y157_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y157_SLICE_X2Y157_BO5),
.O6(CLBLM_R_X3Y157_SLICE_X2Y157_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y157_SLICE_X2Y157_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y157_SLICE_X2Y157_AO5),
.O6(CLBLM_R_X3Y157_SLICE_X2Y157_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y157_SLICE_X3Y157_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y205_IOB_X0Y205_I),
.Q(CLBLM_R_X3Y157_SLICE_X3Y157_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y157_SLICE_X3Y157_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y205_IOB_X0Y206_I),
.Q(CLBLM_R_X3Y157_SLICE_X3Y157_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y157_SLICE_X3Y157_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y219_IOB_X0Y220_I),
.Q(CLBLM_R_X3Y157_SLICE_X3Y157_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y157_SLICE_X3Y157_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y221_IOB_X0Y221_I),
.Q(CLBLM_R_X3Y157_SLICE_X3Y157_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y157_SLICE_X3Y157_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y157_SLICE_X3Y157_DO5),
.O6(CLBLM_R_X3Y157_SLICE_X3Y157_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y157_SLICE_X3Y157_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y157_SLICE_X3Y157_CO5),
.O6(CLBLM_R_X3Y157_SLICE_X3Y157_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y157_SLICE_X3Y157_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y157_SLICE_X3Y157_BO5),
.O6(CLBLM_R_X3Y157_SLICE_X3Y157_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y157_SLICE_X3Y157_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y157_SLICE_X3Y157_AO5),
.O6(CLBLM_R_X3Y157_SLICE_X3Y157_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y158_SLICE_X2Y158_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y225_IOB_X0Y226_I),
.Q(CLBLM_R_X3Y158_SLICE_X2Y158_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y158_SLICE_X2Y158_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y233_IOB_X0Y234_I),
.Q(CLBLM_R_X3Y158_SLICE_X2Y158_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y158_SLICE_X2Y158_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y235_IOB_X0Y236_I),
.Q(CLBLM_R_X3Y158_SLICE_X2Y158_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y158_SLICE_X2Y158_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y237_IOB_X0Y238_I),
.Q(CLBLM_R_X3Y158_SLICE_X2Y158_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y158_SLICE_X2Y158_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y158_SLICE_X2Y158_DO5),
.O6(CLBLM_R_X3Y158_SLICE_X2Y158_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y158_SLICE_X2Y158_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y158_SLICE_X2Y158_CO5),
.O6(CLBLM_R_X3Y158_SLICE_X2Y158_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y158_SLICE_X2Y158_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y158_SLICE_X2Y158_BO5),
.O6(CLBLM_R_X3Y158_SLICE_X2Y158_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y158_SLICE_X2Y158_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y158_SLICE_X2Y158_AO5),
.O6(CLBLM_R_X3Y158_SLICE_X2Y158_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y158_SLICE_X3Y158_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y213_IOB_X0Y214_I),
.Q(CLBLM_R_X3Y158_SLICE_X3Y158_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y158_SLICE_X3Y158_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y217_IOB_X0Y218_I),
.Q(CLBLM_R_X3Y158_SLICE_X3Y158_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y158_SLICE_X3Y158_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y223_IOB_X0Y223_I),
.Q(CLBLM_R_X3Y158_SLICE_X3Y158_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y158_SLICE_X3Y158_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y223_IOB_X0Y224_I),
.Q(CLBLM_R_X3Y158_SLICE_X3Y158_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y158_SLICE_X3Y158_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y158_SLICE_X3Y158_DO5),
.O6(CLBLM_R_X3Y158_SLICE_X3Y158_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y158_SLICE_X3Y158_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y158_SLICE_X3Y158_CO5),
.O6(CLBLM_R_X3Y158_SLICE_X3Y158_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y158_SLICE_X3Y158_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y158_SLICE_X3Y158_BO5),
.O6(CLBLM_R_X3Y158_SLICE_X3Y158_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y158_SLICE_X3Y158_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y158_SLICE_X3Y158_AO5),
.O6(CLBLM_R_X3Y158_SLICE_X3Y158_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y125_SLICE_X6Y125_AO6),
.Q(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y125_SLICE_X6Y125_DO5),
.O6(CLBLM_R_X5Y125_SLICE_X6Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y125_SLICE_X6Y125_CO5),
.O6(CLBLM_R_X5Y125_SLICE_X6Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y125_SLICE_X6Y125_BO5),
.O6(CLBLM_R_X5Y125_SLICE_X6Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff699600006996)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_ALUT (
.I0(BRAM_L_X6Y125_RAMB18_X0Y50_DO2),
.I1(CLBLM_R_X7Y125_SLICE_X8Y125_C5Q),
.I2(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.I3(CLBLM_R_X5Y125_SLICE_X7Y125_BQ),
.I4(LIOB33_X0Y147_IOB_X0Y148_I),
.I5(LIOB33_X0Y17_IOB_X0Y17_I),
.O5(CLBLM_R_X5Y125_SLICE_X6Y125_AO5),
.O6(CLBLM_R_X5Y125_SLICE_X6Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y125_SLICE_X7Y125_AO6),
.Q(CLBLM_R_X5Y125_SLICE_X7Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y125_SLICE_X7Y125_BO6),
.Q(CLBLM_R_X5Y125_SLICE_X7Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y125_SLICE_X7Y125_CO6),
.Q(CLBLM_R_X5Y125_SLICE_X7Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc5aa5a55a)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_DLUT (
.I0(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.I1(LIOB33_X0Y1_IOB_X0Y2_I),
.I2(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.I3(BRAM_L_X6Y125_RAMB18_X0Y50_DO2),
.I4(CLBLM_R_X5Y125_SLICE_X7Y125_BO5),
.I5(LIOB33_X0Y147_IOB_X0Y148_I),
.O5(CLBLM_R_X5Y125_SLICE_X7Y125_DO5),
.O6(CLBLM_R_X5Y125_SLICE_X7Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000069966996)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_CLUT (
.I0(BRAM_L_X6Y125_RAMB18_X0Y50_DO1),
.I1(CLBLM_R_X5Y125_SLICE_X7Y125_CQ),
.I2(CLBLM_R_X7Y125_SLICE_X8Y125_B5Q),
.I3(CLBLM_R_X5Y125_SLICE_X7Y125_AQ),
.I4(LIOB33_X0Y51_IOB_X0Y51_I),
.I5(LIOB33_X0Y147_IOB_X0Y148_I),
.O5(CLBLM_R_X5Y125_SLICE_X7Y125_CO5),
.O6(CLBLM_R_X5Y125_SLICE_X7Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf099f0663333cccc)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_BLUT (
.I0(BRAM_L_X6Y125_RAMB18_X0Y50_DO2),
.I1(CLBLM_R_X5Y125_SLICE_X7Y125_BQ),
.I2(LIOB33_X0Y65_IOB_X0Y66_I),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(CLBLM_R_X7Y125_SLICE_X8Y125_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y125_SLICE_X7Y125_BO5),
.O6(CLBLM_R_X5Y125_SLICE_X7Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb88b8bb80f0ff0f0)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_ALUT (
.I0(LIOB33_X0Y65_IOB_X0Y65_I),
.I1(LIOB33_X0Y147_IOB_X0Y148_I),
.I2(CLBLM_R_X5Y125_SLICE_X7Y125_AQ),
.I3(BRAM_L_X6Y125_RAMB18_X0Y50_DO1),
.I4(CLBLM_R_X7Y125_SLICE_X8Y125_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y125_SLICE_X7Y125_AO5),
.O6(CLBLM_R_X5Y125_SLICE_X7Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y126_SLICE_X6Y126_AO6),
.Q(CLBLM_R_X5Y126_SLICE_X6Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y126_SLICE_X6Y126_BO6),
.Q(CLBLM_R_X5Y126_SLICE_X6Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y126_SLICE_X6Y126_DO5),
.O6(CLBLM_R_X5Y126_SLICE_X6Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff699600006996)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_CLUT (
.I0(CLBLM_R_X5Y126_SLICE_X6Y126_BQ),
.I1(BRAM_L_X6Y125_RAMB18_X0Y50_DO3),
.I2(CLBLM_R_X5Y126_SLICE_X7Y126_B5Q),
.I3(CLBLM_R_X5Y126_SLICE_X6Y126_AO5),
.I4(LIOB33_X0Y147_IOB_X0Y148_I),
.I5(LIOB33_X0Y3_IOB_X0Y3_I),
.O5(CLBLM_R_X5Y126_SLICE_X6Y126_CO5),
.O6(CLBLM_R_X5Y126_SLICE_X6Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8bb8b88bb88b8bb8)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_BLUT (
.I0(LIOB33_X0Y51_IOB_X0Y52_I),
.I1(LIOB33_X0Y147_IOB_X0Y148_I),
.I2(CLBLM_R_X5Y126_SLICE_X6Y126_AQ),
.I3(CLBLM_R_X7Y126_SLICE_X8Y126_D5Q),
.I4(CLBLM_R_X5Y126_SLICE_X6Y126_BQ),
.I5(BRAM_L_X6Y125_RAMB18_X0Y50_DO3),
.O5(CLBLM_R_X5Y126_SLICE_X6Y126_BO5),
.O6(CLBLM_R_X5Y126_SLICE_X6Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haac3aa3c0f0ff0f0)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_ALUT (
.I0(LIOB33_X0Y67_IOB_X0Y67_I),
.I1(BRAM_L_X6Y125_RAMB18_X0Y50_DO3),
.I2(CLBLM_R_X5Y126_SLICE_X6Y126_AQ),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(CLBLM_R_X7Y126_SLICE_X8Y126_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y126_SLICE_X6Y126_AO5),
.O6(CLBLM_R_X5Y126_SLICE_X6Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y126_SLICE_X6Y126_CO6),
.Q(CLBLM_R_X5Y126_SLICE_X7Y126_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y126_SLICE_X7Y126_AO6),
.Q(CLBLM_R_X5Y126_SLICE_X7Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y126_SLICE_X7Y126_BO6),
.Q(CLBLM_R_X5Y126_SLICE_X7Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y126_SLICE_X7Y126_DO5),
.O6(CLBLM_R_X5Y126_SLICE_X7Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdeed1221edde2112)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_CLUT (
.I0(BRAM_L_X6Y125_RAMB18_X0Y50_DO4),
.I1(LIOB33_X0Y147_IOB_X0Y148_I),
.I2(CLBLM_R_X5Y126_SLICE_X7Y126_BQ),
.I3(CLBLM_R_X5Y126_SLICE_X7Y126_AO5),
.I4(LIOB33_X0Y3_IOB_X0Y4_I),
.I5(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.O5(CLBLM_R_X5Y126_SLICE_X7Y126_CO5),
.O6(CLBLM_R_X5Y126_SLICE_X7Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff69ff9600690096)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_BLUT (
.I0(CLBLM_R_X7Y129_SLICE_X9Y129_A5Q),
.I1(CLBLM_R_X5Y126_SLICE_X7Y126_BQ),
.I2(CLBLM_R_X5Y126_SLICE_X7Y126_AQ),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(BRAM_L_X6Y125_RAMB18_X0Y50_DO4),
.I5(LIOB33_X0Y17_IOB_X0Y18_I),
.O5(CLBLM_R_X5Y126_SLICE_X7Y126_BO5),
.O6(CLBLM_R_X5Y126_SLICE_X7Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haac3aa3c3c3c3c3c)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_ALUT (
.I0(LIOB33_X0Y67_IOB_X0Y68_I),
.I1(CLBLM_R_X7Y129_SLICE_X9Y129_A5Q),
.I2(CLBLM_R_X5Y126_SLICE_X7Y126_AQ),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(BRAM_L_X6Y125_RAMB18_X0Y50_DO4),
.I5(1'b1),
.O5(CLBLM_R_X5Y126_SLICE_X7Y126_AO5),
.O6(CLBLM_R_X5Y126_SLICE_X7Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X6Y127_AO6),
.Q(CLBLM_R_X5Y127_SLICE_X6Y127_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X6Y127_CO5),
.Q(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X6Y127_BO6),
.Q(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X6Y127_DO6),
.Q(CLBLM_R_X5Y127_SLICE_X6Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f066999966)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_DLUT (
.I0(BRAM_L_X6Y125_RAMB18_X0Y50_DO0),
.I1(CLBLM_R_X5Y127_SLICE_X6Y127_CQ),
.I2(LIOB33_SING_X0Y0_IOB_X0Y0_I),
.I3(CLBLM_R_X5Y127_SLICE_X6Y127_CO6),
.I4(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.I5(LIOB33_X0Y147_IOB_X0Y148_I),
.O5(CLBLM_R_X5Y127_SLICE_X6Y127_DO5),
.O6(CLBLM_R_X5Y127_SLICE_X6Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0ff0f0cca5cc5a)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_CLUT (
.I0(BRAM_L_X6Y125_RAMB18_X0Y50_DO0),
.I1(LIOB33_X0Y63_IOB_X0Y64_I),
.I2(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(CLBLM_R_X7Y127_SLICE_X8Y127_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y127_SLICE_X6Y127_CO5),
.O6(CLBLM_R_X5Y127_SLICE_X6Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa3caac3aac3aa3c)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.I2(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(BRAM_L_X6Y125_RAMB18_X0Y50_DO0),
.I5(CLBLM_R_X7Y127_SLICE_X8Y127_A5Q),
.O5(CLBLM_R_X5Y127_SLICE_X6Y127_BO5),
.O6(CLBLM_R_X5Y127_SLICE_X6Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff96009666666666)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_ALUT (
.I0(CLBLM_R_X7Y129_SLICE_X9Y129_B5Q),
.I1(CLBLM_R_X5Y127_SLICE_X6Y127_B5Q),
.I2(BRAM_L_X6Y125_RAMB18_X0Y50_DO6),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(LIOB33_X0Y69_IOB_X0Y70_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y127_SLICE_X6Y127_AO5),
.O6(CLBLM_R_X5Y127_SLICE_X6Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X7Y127_DO6),
.Q(CLBLM_R_X5Y127_SLICE_X7Y127_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X7Y127_AO6),
.Q(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X7Y127_BO6),
.Q(CLBLM_R_X5Y127_SLICE_X7Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X7Y127_CO6),
.Q(CLBLM_R_X5Y127_SLICE_X7Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y127_SLICE_X5Y127_BO6),
.Q(CLBLM_R_X5Y127_SLICE_X7Y127_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f066999966)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_DLUT (
.I0(CLBLM_R_X5Y127_SLICE_X7Y127_BQ),
.I1(BRAM_L_X6Y125_RAMB18_X0Y50_DO5),
.I2(LIOB33_X0Y5_IOB_X0Y5_I),
.I3(CLBLM_R_X5Y127_SLICE_X7Y127_AO5),
.I4(CLBLM_R_X5Y127_SLICE_X7Y127_B5Q),
.I5(LIOB33_X0Y147_IOB_X0Y148_I),
.O5(CLBLM_R_X5Y127_SLICE_X7Y127_DO5),
.O6(CLBLM_R_X5Y127_SLICE_X7Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf066f099f099f066)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_CLUT (
.I0(BRAM_L_X6Y125_RAMB18_X0Y50_DO6),
.I1(CLBLM_R_X5Y127_SLICE_X7Y127_CQ),
.I2(LIOB33_X0Y5_IOB_X0Y6_I),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(CLBLM_R_X5Y127_SLICE_X6Y127_AO5),
.I5(CLBLL_L_X4Y127_SLICE_X5Y127_AQ),
.O5(CLBLM_R_X5Y127_SLICE_X7Y127_CO5),
.O6(CLBLM_R_X5Y127_SLICE_X7Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc5acca5cca5cc5a)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_BLUT (
.I0(CLBLM_R_X7Y128_SLICE_X8Y128_A5Q),
.I1(LIOB33_X0Y19_IOB_X0Y19_I),
.I2(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(CLBLM_R_X5Y127_SLICE_X7Y127_BQ),
.I5(BRAM_L_X6Y125_RAMB18_X0Y50_DO5),
.O5(CLBLM_R_X5Y127_SLICE_X7Y127_BO5),
.O6(CLBLM_R_X5Y127_SLICE_X7Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff9600965a5a5a5a)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_ALUT (
.I0(CLBLM_R_X7Y128_SLICE_X8Y128_A5Q),
.I1(BRAM_L_X6Y125_RAMB18_X0Y50_DO5),
.I2(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(LIOB33_X0Y69_IOB_X0Y69_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y127_SLICE_X7Y127_AO5),
.O6(CLBLM_R_X5Y127_SLICE_X7Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X6Y128_AO6),
.Q(CLBLM_R_X5Y128_SLICE_X6Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X6Y128_BO6),
.Q(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y128_SLICE_X6Y128_DO5),
.O6(CLBLM_R_X5Y128_SLICE_X6Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y128_SLICE_X6Y128_CO5),
.O6(CLBLM_R_X5Y128_SLICE_X6Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff69ff9600690096)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_BLUT (
.I0(CLBLM_L_X8Y130_SLICE_X10Y130_B5Q),
.I1(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.I2(CLBLM_R_X5Y128_SLICE_X6Y128_AQ),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(BRAM_L_X6Y125_RAMB18_X0Y50_DO19),
.I5(LIOB33_X0Y25_IOB_X0Y25_I),
.O5(CLBLM_R_X5Y128_SLICE_X6Y128_BO5),
.O6(CLBLM_R_X5Y128_SLICE_X6Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hed21de125a5a5a5a)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_ALUT (
.I0(CLBLM_L_X8Y130_SLICE_X10Y130_B5Q),
.I1(LIOB33_X0Y147_IOB_X0Y148_I),
.I2(CLBLM_R_X5Y128_SLICE_X6Y128_AQ),
.I3(LIOB33_X0Y75_IOB_X0Y75_I),
.I4(BRAM_L_X6Y125_RAMB18_X0Y50_DO19),
.I5(1'b1),
.O5(CLBLM_R_X5Y128_SLICE_X6Y128_AO5),
.O6(CLBLM_R_X5Y128_SLICE_X6Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y129_SLICE_X7Y129_AO6),
.Q(CLBLM_R_X5Y128_SLICE_X7Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y128_SLICE_X7Y128_DO5),
.O6(CLBLM_R_X5Y128_SLICE_X7Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y128_SLICE_X7Y128_CO5),
.O6(CLBLM_R_X5Y128_SLICE_X7Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y128_SLICE_X7Y128_BO5),
.O6(CLBLM_R_X5Y128_SLICE_X7Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y128_SLICE_X7Y128_AO5),
.O6(CLBLM_R_X5Y128_SLICE_X7Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y129_SLICE_X6Y129_CO6),
.Q(CLBLM_R_X5Y129_SLICE_X6Y129_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y129_SLICE_X6Y129_AO6),
.Q(CLBLM_R_X5Y129_SLICE_X6Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y129_SLICE_X6Y129_BO6),
.Q(CLBLM_R_X5Y129_SLICE_X6Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff699600006996)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_DLUT (
.I0(CLBLM_R_X5Y129_SLICE_X7Y129_AQ),
.I1(CLBLM_R_X5Y129_SLICE_X6Y129_AQ),
.I2(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.I3(CLBLM_R_X5Y130_SLICE_X6Y130_AO5),
.I4(LIOB33_X0Y147_IOB_X0Y148_I),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_R_X5Y129_SLICE_X6Y129_DO5),
.O6(CLBLM_R_X5Y129_SLICE_X6Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f066999966)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_CLUT (
.I0(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.I1(CLBLM_R_X5Y128_SLICE_X6Y128_AO5),
.I2(LIOB33_X0Y9_IOB_X0Y10_I),
.I3(CLBLM_R_X5Y129_SLICE_X6Y129_A5Q),
.I4(BRAM_L_X6Y125_RAMB18_X0Y50_DO19),
.I5(LIOB33_X0Y147_IOB_X0Y148_I),
.O5(CLBLM_R_X5Y129_SLICE_X6Y129_CO5),
.O6(CLBLM_R_X5Y129_SLICE_X6Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff690069ff960096)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_BLUT (
.I0(CLBLM_R_X7Y136_SLICE_X8Y136_A5Q),
.I1(CLBLM_R_X5Y129_SLICE_X6Y129_BQ),
.I2(BRAM_L_X6Y125_RAMB18_X0Y50_DO17),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(LIOB33_X0Y23_IOB_X0Y23_I),
.I5(CLBLL_L_X4Y129_SLICE_X4Y129_AQ),
.O5(CLBLM_R_X5Y129_SLICE_X6Y129_BO5),
.O6(CLBLM_R_X5Y129_SLICE_X6Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hed21ed21de12de12)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_ALUT (
.I0(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.I1(LIOB33_X0Y147_IOB_X0Y148_I),
.I2(CLBLM_R_X5Y129_SLICE_X6Y129_AQ),
.I3(LIOB33_X0Y59_IOB_X0Y59_I),
.I4(1'b1),
.I5(CLBLM_R_X5Y130_SLICE_X6Y130_AO5),
.O5(CLBLM_R_X5Y129_SLICE_X6Y129_AO5),
.O6(CLBLM_R_X5Y129_SLICE_X6Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y129_SLICE_X7Y129_CO6),
.Q(CLBLM_R_X5Y129_SLICE_X7Y129_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y129_SLICE_X6Y129_DO6),
.Q(CLBLM_R_X5Y129_SLICE_X7Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y129_SLICE_X7Y129_BO6),
.Q(CLBLM_R_X5Y129_SLICE_X7Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdeed1221edde2112)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_DLUT (
.I0(BRAM_L_X6Y125_RAMB18_X0Y50_DO16),
.I1(LIOB33_X0Y147_IOB_X0Y148_I),
.I2(CLBLM_R_X5Y129_SLICE_X7Y129_BQ),
.I3(CLBLM_R_X5Y129_SLICE_X7Y129_AO5),
.I4(LIOB33_X0Y7_IOB_X0Y7_I),
.I5(CLBLM_R_X5Y130_SLICE_X7Y130_CQ),
.O5(CLBLM_R_X5Y129_SLICE_X7Y129_DO5),
.O6(CLBLM_R_X5Y129_SLICE_X7Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f066999966)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_CLUT (
.I0(BRAM_L_X6Y125_RAMB18_X0Y50_DO17),
.I1(CLBLM_R_X5Y129_SLICE_X6Y129_BQ),
.I2(LIOB33_X0Y7_IOB_X0Y8_I),
.I3(CLBLL_L_X4Y129_SLICE_X5Y129_BO5),
.I4(CLBLM_R_X5Y129_SLICE_X7Y129_B5Q),
.I5(LIOB33_X0Y147_IOB_X0Y148_I),
.O5(CLBLM_R_X5Y129_SLICE_X7Y129_CO5),
.O6(CLBLM_R_X5Y129_SLICE_X7Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa3caac3aac3aa3c)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_BLUT (
.I0(LIOB33_X0Y21_IOB_X0Y22_I),
.I1(CLBLM_R_X5Y129_SLICE_X7Y129_BQ),
.I2(CLBLM_R_X5Y128_SLICE_X7Y128_AQ),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(BRAM_L_X6Y125_RAMB18_X0Y50_DO16),
.I5(CLBLM_R_X7Y129_SLICE_X8Y129_A5Q),
.O5(CLBLM_R_X5Y129_SLICE_X7Y129_BO5),
.O6(CLBLM_R_X5Y129_SLICE_X7Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he2d1d1e25555aaaa)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_ALUT (
.I0(CLBLM_R_X7Y129_SLICE_X8Y129_A5Q),
.I1(LIOB33_X0Y147_IOB_X0Y148_I),
.I2(LIOB33_X0Y71_IOB_X0Y72_I),
.I3(BRAM_L_X6Y125_RAMB18_X0Y50_DO16),
.I4(CLBLM_R_X5Y128_SLICE_X7Y128_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y129_SLICE_X7Y129_AO5),
.O6(CLBLM_R_X5Y129_SLICE_X7Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y130_SLICE_X5Y130_CO6),
.Q(CLBLM_R_X5Y130_SLICE_X6Y130_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y130_SLICE_X6Y130_AO6),
.Q(CLBLM_R_X5Y130_SLICE_X6Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y130_SLICE_X6Y130_BO6),
.Q(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y130_SLICE_X6Y130_CO6),
.Q(CLBLM_R_X5Y130_SLICE_X6Y130_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y130_SLICE_X4Y130_CO6),
.Q(CLBLM_R_X5Y130_SLICE_X6Y130_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f066999966)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_DLUT (
.I0(BRAM_L_X6Y125_RAMB18_X0Y50_DO20),
.I1(CLBLM_R_X5Y130_SLICE_X7Y130_A5Q),
.I2(LIOB33_X0Y11_IOB_X0Y11_I),
.I3(CLBLL_L_X4Y131_SLICE_X4Y131_AO5),
.I4(CLBLL_L_X4Y131_SLICE_X5Y131_BQ),
.I5(LIOB33_X0Y147_IOB_X0Y148_I),
.O5(CLBLM_R_X5Y130_SLICE_X6Y130_DO5),
.O6(CLBLM_R_X5Y130_SLICE_X6Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa3cc3c33c)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_CLUT (
.I0(LIOB33_X0Y15_IOB_X0Y15_I),
.I1(CLBLM_R_X5Y130_SLICE_X6Y130_CQ),
.I2(CLBLM_R_X5Y131_SLICE_X6Y131_BO5),
.I3(CLBLM_R_X5Y131_SLICE_X6Y131_CQ),
.I4(BRAM_L_X6Y130_RAMB18_X0Y52_DO0),
.I5(LIOB33_X0Y147_IOB_X0Y148_I),
.O5(CLBLM_R_X5Y130_SLICE_X6Y130_CO5),
.O6(CLBLM_R_X5Y130_SLICE_X6Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff690069ff960096)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_BLUT (
.I0(CLBLM_R_X5Y130_SLICE_X6Y130_AQ),
.I1(BRAM_L_X6Y130_RAMB18_X0Y52_DO19),
.I2(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(LIOB33_X0Y91_IOB_X0Y91_I),
.I5(CLBLM_R_X3Y131_SLICE_X2Y131_B5Q),
.O5(CLBLM_R_X5Y130_SLICE_X6Y130_BO5),
.O6(CLBLM_R_X5Y130_SLICE_X6Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haac3aa3cc3c33c3c)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_ALUT (
.I0(LIOB33_X0Y143_IOB_X0Y143_I),
.I1(BRAM_L_X6Y130_RAMB18_X0Y52_DO19),
.I2(CLBLM_R_X5Y130_SLICE_X6Y130_AQ),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(CLBLM_R_X3Y131_SLICE_X2Y131_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y130_SLICE_X6Y130_AO5),
.O6(CLBLM_R_X5Y130_SLICE_X6Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y130_SLICE_X6Y130_DO6),
.Q(CLBLM_R_X5Y130_SLICE_X7Y130_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y130_SLICE_X7Y130_AO6),
.Q(CLBLM_R_X5Y130_SLICE_X7Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y130_SLICE_X3Y130_CO6),
.Q(CLBLM_R_X5Y130_SLICE_X7Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y129_SLICE_X7Y129_DO6),
.Q(CLBLM_R_X5Y130_SLICE_X7Y130_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y130_SLICE_X7Y130_DO5),
.O6(CLBLM_R_X5Y130_SLICE_X7Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y130_SLICE_X7Y130_CO5),
.O6(CLBLM_R_X5Y130_SLICE_X7Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y130_SLICE_X7Y130_BO5),
.O6(CLBLM_R_X5Y130_SLICE_X7Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6666666666666666)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_ALUT (
.I0(CLBLL_L_X4Y131_SLICE_X4Y131_DQ),
.I1(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO2),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y130_SLICE_X7Y130_AO5),
.O6(CLBLM_R_X5Y130_SLICE_X7Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X6Y131_DO6),
.Q(CLBLM_R_X5Y131_SLICE_X6Y131_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X6Y131_AO6),
.Q(CLBLM_R_X5Y131_SLICE_X6Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X6Y131_CO6),
.Q(CLBLM_R_X5Y131_SLICE_X6Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000069966996)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_DLUT (
.I0(BRAM_L_X6Y130_RAMB18_X0Y52_DO4),
.I1(CLBLM_R_X5Y131_SLICE_X6Y131_A5Q),
.I2(CLBLM_R_X5Y131_SLICE_X7Y131_BO5),
.I3(CLBLM_R_X5Y131_SLICE_X7Y131_CQ),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(LIOB33_X0Y147_IOB_X0Y148_I),
.O5(CLBLM_R_X5Y131_SLICE_X6Y131_DO5),
.O6(CLBLM_R_X5Y131_SLICE_X6Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff690069ff960096)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_CLUT (
.I0(BRAM_L_X6Y130_RAMB18_X0Y52_DO0),
.I1(CLBLM_R_X5Y131_SLICE_X6Y131_CQ),
.I2(CLBLM_L_X8Y132_SLICE_X11Y132_A5Q),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(LIOB33_X0Y29_IOB_X0Y30_I),
.I5(CLBLM_R_X5Y131_SLICE_X7Y131_A5Q),
.O5(CLBLM_R_X5Y131_SLICE_X6Y131_CO5),
.O6(CLBLM_R_X5Y131_SLICE_X6Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haac3aa3c3c3c3c3c)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_BLUT (
.I0(LIOB33_X0Y79_IOB_X0Y80_I),
.I1(CLBLM_L_X8Y132_SLICE_X11Y132_A5Q),
.I2(CLBLM_R_X5Y131_SLICE_X7Y131_A5Q),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(BRAM_L_X6Y130_RAMB18_X0Y52_DO0),
.I5(1'b1),
.O5(CLBLM_R_X5Y131_SLICE_X6Y131_BO5),
.O6(CLBLM_R_X5Y131_SLICE_X6Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5a5a5a5a5a)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_ALUT (
.I0(CLBLM_R_X5Y129_SLICE_X6Y129_AQ),
.I1(1'b1),
.I2(BRAM_L_X6Y140_RAMB18_X0Y56_DO3),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y131_SLICE_X6Y131_AO5),
.O6(CLBLM_R_X5Y131_SLICE_X6Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X6Y131_BO6),
.Q(CLBLM_R_X5Y131_SLICE_X7Y131_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X7Y131_AO6),
.Q(CLBLM_R_X5Y131_SLICE_X7Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X7Y131_BO6),
.Q(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X7Y131_CO6),
.Q(CLBLM_R_X5Y131_SLICE_X7Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_DLUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y54_DO23),
.I1(BRAM_R_X17Y135_RAMB18_X1Y54_DO22),
.I2(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO7),
.I3(CLBLL_L_X4Y128_SLICE_X5Y128_AQ),
.I4(BRAM_R_X17Y135_RAMB18_X1Y54_DO23),
.I5(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO6),
.O5(CLBLM_R_X5Y131_SLICE_X7Y131_DO5),
.O6(CLBLM_R_X5Y131_SLICE_X7Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0069699696)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_CLUT (
.I0(BRAM_L_X6Y130_RAMB18_X0Y52_DO4),
.I1(CLBLM_R_X5Y131_SLICE_X7Y131_CQ),
.I2(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.I3(LIOB33_X0Y53_IOB_X0Y54_I),
.I4(CLBLM_L_X8Y136_SLICE_X10Y136_A5Q),
.I5(LIOB33_X0Y147_IOB_X0Y148_I),
.O5(CLBLM_R_X5Y131_SLICE_X7Y131_CO5),
.O6(CLBLM_R_X5Y131_SLICE_X7Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf099f06666666666)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_BLUT (
.I0(CLBLM_L_X8Y136_SLICE_X10Y136_A5Q),
.I1(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.I2(LIOB33_X0Y83_IOB_X0Y84_I),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(BRAM_L_X6Y130_RAMB18_X0Y52_DO4),
.I5(1'b1),
.O5(CLBLM_R_X5Y131_SLICE_X7Y131_BO5),
.O6(CLBLM_R_X5Y131_SLICE_X7Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555555aaaaaaaa)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_ALUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO6),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y127_SLICE_X7Y127_CQ),
.O5(CLBLM_R_X5Y131_SLICE_X7Y131_AO5),
.O6(CLBLM_R_X5Y131_SLICE_X7Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y132_SLICE_X5Y132_DO6),
.Q(CLBLM_R_X5Y132_SLICE_X6Y132_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y132_SLICE_X6Y132_AO6),
.Q(CLBLM_R_X5Y132_SLICE_X6Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y132_SLICE_X6Y132_BO6),
.Q(CLBLM_R_X5Y132_SLICE_X6Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf6f9f9f606090906)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_DLUT (
.I0(CLBLM_R_X5Y132_SLICE_X6Y132_BQ),
.I1(CLBLM_R_X7Y132_SLICE_X8Y132_BQ),
.I2(LIOB33_X0Y147_IOB_X0Y148_I),
.I3(BRAM_L_X6Y130_RAMB18_X0Y52_DO3),
.I4(CLBLM_R_X5Y133_SLICE_X6Y133_AO5),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLM_R_X5Y132_SLICE_X6Y132_DO5),
.O6(CLBLM_R_X5Y132_SLICE_X6Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f06699f0f09966)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_CLUT (
.I0(BRAM_L_X6Y130_RAMB18_X0Y52_DO5),
.I1(CLBLM_R_X7Y132_SLICE_X8Y132_CQ),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(CLBLM_R_X5Y132_SLICE_X6Y132_AO5),
.I4(LIOB33_X0Y147_IOB_X0Y148_I),
.I5(CLBLL_L_X4Y132_SLICE_X5Y132_AQ),
.O5(CLBLM_R_X5Y132_SLICE_X6Y132_CO5),
.O6(CLBLM_R_X5Y132_SLICE_X6Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb1e4e4b1e4b1b1e4)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_BLUT (
.I0(LIOB33_X0Y147_IOB_X0Y148_I),
.I1(CLBLM_R_X5Y132_SLICE_X6Y132_BQ),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(CLBLM_R_X5Y133_SLICE_X6Y133_AQ),
.I4(CLBLM_R_X7Y134_SLICE_X9Y134_B5Q),
.I5(BRAM_L_X6Y130_RAMB18_X0Y52_DO3),
.O5(CLBLM_R_X5Y132_SLICE_X6Y132_BO5),
.O6(CLBLM_R_X5Y132_SLICE_X6Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hebbe41140ff00ff0)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_ALUT (
.I0(LIOB33_X0Y147_IOB_X0Y148_I),
.I1(BRAM_L_X6Y130_RAMB18_X0Y52_DO5),
.I2(CLBLM_R_X5Y132_SLICE_X6Y132_AQ),
.I3(CLBLM_L_X10Y135_SLICE_X12Y135_A5Q),
.I4(LIOB33_X0Y85_IOB_X0Y85_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y132_SLICE_X6Y132_AO5),
.O6(CLBLM_R_X5Y132_SLICE_X6Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y132_SLICE_X4Y132_DO6),
.Q(CLBLM_R_X5Y132_SLICE_X7Y132_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y132_SLICE_X5Y132_CO6),
.Q(CLBLM_R_X5Y132_SLICE_X7Y132_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y132_SLICE_X7Y132_AO6),
.Q(CLBLM_R_X5Y132_SLICE_X7Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y132_SLICE_X7Y132_BO6),
.Q(CLBLM_R_X5Y132_SLICE_X7Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f30cfc03f30cfc0)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y157_SLICE_X3Y157_CQ),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I3(CLBLM_R_X5Y132_SLICE_X7Y132_CO6),
.I4(CLBLM_R_X5Y127_SLICE_X6Y127_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y132_SLICE_X7Y132_DO5),
.O6(CLBLM_R_X5Y132_SLICE_X7Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_CLUT (
.I0(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO5),
.I1(BRAM_R_X17Y135_RAMB18_X1Y54_DO22),
.I2(CLBLM_R_X5Y127_SLICE_X6Y127_B5Q),
.I3(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO6),
.I4(BRAM_L_X6Y135_RAMB18_X0Y54_DO22),
.I5(BRAM_R_X17Y135_RAMB18_X1Y54_DO21),
.O5(CLBLM_R_X5Y132_SLICE_X7Y132_CO5),
.O6(CLBLM_R_X5Y132_SLICE_X7Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ffff00ff00)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X5Y132_SLICE_X6Y132_BQ),
.I4(1'b1),
.I5(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO3),
.O5(CLBLM_R_X5Y132_SLICE_X7Y132_BO5),
.O6(CLBLM_R_X5Y132_SLICE_X7Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cc33cc33cc33cc)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y132_SLICE_X6Y132_B5Q),
.I2(1'b1),
.I3(BRAM_L_X6Y140_RAMB18_X0Y56_DO17),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y132_SLICE_X7Y132_AO5),
.O6(CLBLM_R_X5Y132_SLICE_X7Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X6Y133_AO6),
.Q(CLBLM_R_X5Y133_SLICE_X6Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y133_SLICE_X5Y133_DO6),
.Q(CLBLM_R_X5Y133_SLICE_X6Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f0cf3c03f0cf3c0)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I2(CLBLM_R_X5Y130_SLICE_X6Y130_DQ),
.I3(CLBLM_R_X5Y133_SLICE_X6Y133_CO6),
.I4(CLBLM_R_X3Y147_SLICE_X3Y147_DQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y133_SLICE_X6Y133_DO5),
.O6(CLBLM_R_X5Y133_SLICE_X6Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_CLUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO1),
.I1(BRAM_L_X6Y140_RAMB18_X0Y56_DO18),
.I2(CLBLM_R_X5Y130_SLICE_X6Y130_DQ),
.I3(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO1),
.I4(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO2),
.I5(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO2),
.O5(CLBLM_R_X5Y133_SLICE_X6Y133_CO5),
.O6(CLBLM_R_X5Y133_SLICE_X6Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0ff0f099669966)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_BLUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO7),
.I1(CLBLM_R_X5Y133_SLICE_X7Y133_DO6),
.I2(CLBLM_R_X7Y130_SLICE_X8Y130_B5Q),
.I3(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO7),
.I4(CLBLL_L_X4Y145_SLICE_X4Y145_BQ),
.I5(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.O5(CLBLM_R_X5Y133_SLICE_X6Y133_BO5),
.O6(CLBLM_R_X5Y133_SLICE_X6Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaac33c0ff00ff0)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_ALUT (
.I0(LIOB33_X0Y83_IOB_X0Y83_I),
.I1(BRAM_L_X6Y130_RAMB18_X0Y52_DO3),
.I2(CLBLM_R_X5Y133_SLICE_X6Y133_AQ),
.I3(CLBLM_R_X7Y134_SLICE_X9Y134_B5Q),
.I4(LIOB33_X0Y147_IOB_X0Y148_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y133_SLICE_X6Y133_AO5),
.O6(CLBLM_R_X5Y133_SLICE_X6Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X7Y133_AO6),
.Q(CLBLM_R_X5Y133_SLICE_X7Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X7Y133_BO6),
.Q(CLBLM_R_X5Y133_SLICE_X7Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X7Y133_CO6),
.Q(CLBLM_R_X5Y133_SLICE_X7Y133_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_DLUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO1),
.I1(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO1),
.I2(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO0),
.I3(BRAM_L_X6Y140_RAMB18_X0Y56_DO17),
.I4(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO0),
.I5(CLBLM_R_X7Y130_SLICE_X8Y130_B5Q),
.O5(CLBLM_R_X5Y133_SLICE_X7Y133_DO5),
.O6(CLBLM_R_X5Y133_SLICE_X7Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5a5a5a5a5a)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_CLUT (
.I0(CLBLM_R_X3Y130_SLICE_X2Y130_AQ),
.I1(1'b1),
.I2(BRAM_L_X6Y140_RAMB18_X0Y56_DO0),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y133_SLICE_X7Y133_CO5),
.O6(CLBLM_R_X5Y133_SLICE_X7Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3c3c3c3c3c)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_BLUT (
.I0(1'b1),
.I1(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO2),
.I2(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y133_SLICE_X7Y133_BO5),
.O6(CLBLM_R_X5Y133_SLICE_X7Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffff0000ffff00)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(BRAM_L_X6Y140_RAMB18_X0Y56_DO19),
.I4(CLBLM_R_X5Y129_SLICE_X7Y129_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y133_SLICE_X7Y133_AO5),
.O6(CLBLM_R_X5Y133_SLICE_X7Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f303f30cfc0cfc0)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y155_SLICE_X0Y155_CQ),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I3(CLBLM_R_X5Y135_SLICE_X6Y135_AO6),
.I4(1'b1),
.I5(CLBLL_L_X4Y132_SLICE_X5Y132_AQ),
.O5(CLBLM_R_X5Y134_SLICE_X6Y134_DO5),
.O6(CLBLM_R_X5Y134_SLICE_X6Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_CLUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO7),
.I1(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO7),
.I2(BRAM_L_X6Y140_RAMB18_X0Y56_DO23),
.I3(CLBLL_L_X4Y132_SLICE_X5Y132_A5Q),
.I4(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO6),
.I5(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO6),
.O5(CLBLM_R_X5Y134_SLICE_X6Y134_CO5),
.O6(CLBLM_R_X5Y134_SLICE_X6Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffff000ff00ff0)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X5Y127_SLICE_X7Y127_DQ),
.I3(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO7),
.I4(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO7),
.I5(1'b1),
.O5(CLBLM_R_X5Y134_SLICE_X6Y134_BO5),
.O6(CLBLM_R_X5Y134_SLICE_X6Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333cccc00ffff00)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_ALUT (
.I0(1'b1),
.I1(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO7),
.I2(1'b1),
.I3(CLBLL_L_X4Y134_SLICE_X4Y134_AQ),
.I4(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO7),
.I5(1'b1),
.O5(CLBLM_R_X5Y134_SLICE_X6Y134_AO5),
.O6(CLBLM_R_X5Y134_SLICE_X6Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X7Y134_AO5),
.Q(CLBLM_R_X5Y134_SLICE_X7Y134_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X7Y134_AO6),
.Q(CLBLM_R_X5Y134_SLICE_X7Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X7Y134_BO6),
.Q(CLBLM_R_X5Y134_SLICE_X7Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X7Y134_CO6),
.Q(CLBLM_R_X5Y134_SLICE_X7Y134_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3fcf30c03fcf30c0)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y132_SLICE_X8Y132_CQ),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I3(CLBLM_R_X3Y147_SLICE_X2Y147_BQ),
.I4(CLBLM_R_X7Y134_SLICE_X8Y134_AO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y134_SLICE_X7Y134_DO5),
.O6(CLBLM_R_X5Y134_SLICE_X7Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555555aaaaaaaa)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_CLUT (
.I0(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO4),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y131_SLICE_X7Y131_CQ),
.O5(CLBLM_R_X5Y134_SLICE_X7Y134_CO5),
.O6(CLBLM_R_X5Y134_SLICE_X7Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5a5a5a5a5a)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_BLUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y56_DO23),
.I1(1'b1),
.I2(CLBLL_L_X4Y132_SLICE_X5Y132_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y134_SLICE_X7Y134_BO5),
.O6(CLBLM_R_X5Y134_SLICE_X7Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ccccaa3caa3c)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_ALUT (
.I0(LIOB33_X0Y131_IOB_X0Y131_I),
.I1(CLBLM_R_X5Y134_SLICE_X7Y134_A5Q),
.I2(BRAM_L_X6Y125_RAMB18_X0Y50_DO23),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(BRAM_L_X6Y135_RAMB18_X0Y54_DO7),
.I5(1'b1),
.O5(CLBLM_R_X5Y134_SLICE_X7Y134_AO5),
.O6(CLBLM_R_X5Y134_SLICE_X7Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_DLUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO5),
.I1(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO6),
.I2(BRAM_L_X6Y140_RAMB18_X0Y56_DO22),
.I3(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO6),
.I4(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO5),
.I5(CLBLM_R_X5Y130_SLICE_X6Y130_B5Q),
.O5(CLBLM_R_X5Y135_SLICE_X6Y135_DO5),
.O6(CLBLM_R_X5Y135_SLICE_X6Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_CLUT (
.I0(CLBLM_R_X3Y134_SLICE_X2Y134_AQ),
.I1(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO7),
.I2(BRAM_R_X17Y135_RAMB18_X1Y54_DO23),
.I3(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO7),
.I4(BRAM_L_X6Y135_RAMB18_X0Y54_DO22),
.I5(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO6),
.O5(CLBLM_R_X5Y135_SLICE_X6Y135_CO5),
.O6(CLBLM_R_X5Y135_SLICE_X6Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_BLUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO6),
.I1(BRAM_L_X6Y140_RAMB18_X0Y56_DO22),
.I2(CLBLM_R_X5Y132_SLICE_X7Y132_A5Q),
.I3(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO5),
.I4(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO5),
.I5(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO6),
.O5(CLBLM_R_X5Y135_SLICE_X6Y135_BO5),
.O6(CLBLM_R_X5Y135_SLICE_X6Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_ALUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y56_DO5),
.I1(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO5),
.I2(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO4),
.I3(CLBLL_L_X4Y132_SLICE_X5Y132_AQ),
.I4(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO4),
.I5(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO5),
.O5(CLBLM_R_X5Y135_SLICE_X6Y135_AO5),
.O6(CLBLM_R_X5Y135_SLICE_X6Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y135_SLICE_X7Y135_AO6),
.Q(CLBLM_R_X5Y135_SLICE_X7Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_DLUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y56_DO19),
.I1(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO3),
.I2(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO3),
.I3(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO2),
.I4(CLBLM_R_X5Y129_SLICE_X6Y129_A5Q),
.I5(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO2),
.O5(CLBLM_R_X5Y135_SLICE_X7Y135_DO5),
.O6(CLBLM_R_X5Y135_SLICE_X7Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f990f66f099f066)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_CLUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO7),
.I1(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO7),
.I2(CLBLM_R_X5Y129_SLICE_X6Y129_A5Q),
.I3(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I4(CLBLM_R_X5Y135_SLICE_X7Y135_DO6),
.I5(CLBLM_R_X3Y142_SLICE_X2Y142_AQ),
.O5(CLBLM_R_X5Y135_SLICE_X7Y135_CO5),
.O6(CLBLM_R_X5Y135_SLICE_X7Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_BLUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y54_DO21),
.I1(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO6),
.I2(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO5),
.I3(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO6),
.I4(BRAM_R_X17Y135_RAMB18_X1Y54_DO22),
.I5(CLBLL_L_X4Y131_SLICE_X5Y131_B5Q),
.O5(CLBLM_R_X5Y135_SLICE_X7Y135_BO5),
.O6(CLBLM_R_X5Y135_SLICE_X7Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa55aa55aa55aa)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_ALUT (
.I0(CLBLM_R_X5Y126_SLICE_X7Y126_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO4),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y135_SLICE_X7Y135_AO5),
.O6(CLBLM_R_X5Y135_SLICE_X7Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f99f0990f66f066)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_DLUT (
.I0(CLBLM_R_X5Y137_SLICE_X7Y137_BO6),
.I1(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO7),
.I2(CLBLM_R_X3Y153_SLICE_X2Y153_BQ),
.I3(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I4(CLBLM_R_X5Y129_SLICE_X6Y129_BQ),
.I5(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO7),
.O5(CLBLM_R_X5Y136_SLICE_X6Y136_DO5),
.O6(CLBLM_R_X5Y136_SLICE_X6Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_CLUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO1),
.I1(BRAM_L_X6Y140_RAMB18_X0Y56_DO18),
.I2(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO2),
.I3(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.I4(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO1),
.I5(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO2),
.O5(CLBLM_R_X5Y136_SLICE_X6Y136_CO5),
.O6(CLBLM_R_X5Y136_SLICE_X6Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h74474774b88b8bb8)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_BLUT (
.I0(CLBLL_L_X4Y155_SLICE_X4Y155_BQ),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I2(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO7),
.I3(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO7),
.I4(CLBLM_R_X5Y136_SLICE_X6Y136_AO6),
.I5(CLBLM_R_X5Y132_SLICE_X6Y132_BQ),
.O5(CLBLM_R_X5Y136_SLICE_X6Y136_BO5),
.O6(CLBLM_R_X5Y136_SLICE_X6Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_ALUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y56_DO3),
.I1(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO2),
.I2(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO2),
.I3(CLBLM_R_X5Y132_SLICE_X6Y132_BQ),
.I4(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO3),
.I5(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO3),
.O5(CLBLM_R_X5Y136_SLICE_X6Y136_AO5),
.O6(CLBLM_R_X5Y136_SLICE_X6Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6666ffff66660000)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_DLUT (
.I0(CLBLM_R_X3Y155_SLICE_X3Y155_AQ),
.I1(CLBLL_L_X4Y131_SLICE_X5Y131_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I5(CLBLM_R_X5Y136_SLICE_X7Y136_BO6),
.O5(CLBLM_R_X5Y136_SLICE_X7Y136_DO5),
.O6(CLBLM_R_X5Y136_SLICE_X7Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_CLUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO1),
.I1(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO0),
.I2(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO0),
.I3(BRAM_L_X6Y140_RAMB18_X0Y56_DO17),
.I4(CLBLM_R_X5Y129_SLICE_X7Y129_B5Q),
.I5(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO1),
.O5(CLBLM_R_X5Y136_SLICE_X7Y136_CO5),
.O6(CLBLM_R_X5Y136_SLICE_X7Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_BLUT (
.I0(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO6),
.I1(CLBLL_L_X4Y131_SLICE_X5Y131_CQ),
.I2(BRAM_L_X6Y140_RAMB18_X0Y56_DO6),
.I3(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO5),
.I4(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO5),
.I5(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO6),
.O5(CLBLM_R_X5Y136_SLICE_X7Y136_BO5),
.O6(CLBLM_R_X5Y136_SLICE_X7Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h66f0660f660f66f0)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_ALUT (
.I0(CLBLM_R_X3Y142_SLICE_X2Y142_DQ),
.I1(CLBLM_R_X5Y129_SLICE_X7Y129_B5Q),
.I2(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO7),
.I3(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I4(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO7),
.I5(CLBLM_R_X5Y136_SLICE_X7Y136_CO6),
.O5(CLBLM_R_X5Y136_SLICE_X7Y136_AO5),
.O6(CLBLM_R_X5Y136_SLICE_X7Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h77bb77bb44884488)
  ) CLBLM_R_X5Y137_SLICE_X6Y137_DLUT (
.I0(CLBLL_L_X4Y134_SLICE_X4Y134_AQ),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I2(1'b1),
.I3(CLBLM_R_X3Y145_SLICE_X3Y145_AQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y137_SLICE_X6Y137_BO6),
.O5(CLBLM_R_X5Y137_SLICE_X6Y137_DO5),
.O6(CLBLM_R_X5Y137_SLICE_X6Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h77447744bb88bb88)
  ) CLBLM_R_X5Y137_SLICE_X6Y137_CLUT (
.I0(CLBLM_R_X3Y130_SLICE_X3Y130_BQ),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y137_SLICE_X6Y137_AO6),
.I4(1'b1),
.I5(CLBLL_L_X2Y155_SLICE_X1Y155_AQ),
.O5(CLBLM_R_X5Y137_SLICE_X6Y137_CO5),
.O6(CLBLM_R_X5Y137_SLICE_X6Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X5Y137_SLICE_X6Y137_BLUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO6),
.I1(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO7),
.I2(CLBLL_L_X4Y134_SLICE_X4Y134_AQ),
.I3(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO6),
.I4(BRAM_L_X6Y140_RAMB18_X0Y56_DO23),
.I5(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO7),
.O5(CLBLM_R_X5Y137_SLICE_X6Y137_BO5),
.O6(CLBLM_R_X5Y137_SLICE_X6Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X5Y137_SLICE_X6Y137_ALUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO4),
.I1(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO5),
.I2(CLBLM_R_X3Y130_SLICE_X3Y130_BQ),
.I3(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO4),
.I4(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO5),
.I5(BRAM_L_X6Y140_RAMB18_X0Y56_DO5),
.O5(CLBLM_R_X5Y137_SLICE_X6Y137_AO5),
.O6(CLBLM_R_X5Y137_SLICE_X6Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y137_SLICE_X7Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y137_SLICE_X7Y137_AO6),
.Q(CLBLM_R_X5Y137_SLICE_X7Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2112eddeedde2112)
  ) CLBLM_R_X5Y137_SLICE_X7Y137_DLUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y56_DO7),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I2(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO7),
.I3(CLBLM_R_X5Y137_SLICE_X7Y137_CO6),
.I4(CLBLM_R_X5Y126_SLICE_X7Y126_BQ),
.I5(CLBLM_R_X3Y153_SLICE_X3Y153_BQ),
.O5(CLBLM_R_X5Y137_SLICE_X7Y137_DO5),
.O6(CLBLM_R_X5Y137_SLICE_X7Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X5Y137_SLICE_X7Y137_CLUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO4),
.I1(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO3),
.I2(CLBLM_R_X5Y126_SLICE_X7Y126_BQ),
.I3(BRAM_L_X6Y140_RAMB18_X0Y56_DO4),
.I4(BRAM_L_X6Y140_RAMB18_X0Y56_DO3),
.I5(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO4),
.O5(CLBLM_R_X5Y137_SLICE_X7Y137_CO5),
.O6(CLBLM_R_X5Y137_SLICE_X7Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X5Y137_SLICE_X7Y137_BLUT (
.I0(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO1),
.I1(BRAM_L_X6Y140_RAMB18_X0Y56_DO1),
.I2(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO0),
.I3(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO1),
.I4(CLBLM_R_X5Y129_SLICE_X6Y129_BQ),
.I5(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO0),
.O5(CLBLM_R_X5Y137_SLICE_X7Y137_BO5),
.O6(CLBLM_R_X5Y137_SLICE_X7Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff00ff00ff00ff0)
  ) CLBLM_R_X5Y137_SLICE_X7Y137_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO5),
.I3(CLBLM_R_X5Y127_SLICE_X7Y127_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y137_SLICE_X7Y137_AO5),
.O6(CLBLM_R_X5Y137_SLICE_X7Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y138_SLICE_X6Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y138_SLICE_X6Y138_AO6),
.Q(CLBLM_R_X5Y138_SLICE_X6Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y138_SLICE_X6Y138_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.Q(CLBLM_R_X5Y138_SLICE_X6Y138_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7b487b487b487b48)
  ) CLBLM_R_X5Y138_SLICE_X6Y138_DLUT (
.I0(CLBLL_L_X4Y127_SLICE_X5Y127_AQ),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I2(CLBLM_R_X3Y153_SLICE_X3Y153_CQ),
.I3(CLBLM_R_X5Y138_SLICE_X6Y138_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y138_SLICE_X6Y138_DO5),
.O6(CLBLM_R_X5Y138_SLICE_X6Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X5Y138_SLICE_X6Y138_CLUT (
.I0(CLBLL_L_X4Y127_SLICE_X5Y127_AQ),
.I1(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO6),
.I2(BRAM_L_X6Y140_RAMB18_X0Y56_DO5),
.I3(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO5),
.I4(BRAM_L_X6Y140_RAMB18_X0Y56_DO6),
.I5(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO6),
.O5(CLBLM_R_X5Y138_SLICE_X6Y138_CO5),
.O6(CLBLM_R_X5Y138_SLICE_X6Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff00ff00ff00ff0)
  ) CLBLM_R_X5Y138_SLICE_X6Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X3Y130_SLICE_X3Y130_BQ),
.I3(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO5),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y138_SLICE_X6Y138_BO5),
.O6(CLBLM_R_X5Y138_SLICE_X6Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa55aa55aa55aa)
  ) CLBLM_R_X5Y138_SLICE_X6Y138_ALUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO4),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_L_X4Y131_SLICE_X5Y131_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y138_SLICE_X6Y138_AO5),
.O6(CLBLM_R_X5Y138_SLICE_X6Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y138_SLICE_X7Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y138_SLICE_X7Y138_AO6),
.Q(CLBLM_R_X5Y138_SLICE_X7Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X5Y138_SLICE_X7Y138_DLUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y56_DO18),
.I1(CLBLM_R_X5Y126_SLICE_X7Y126_B5Q),
.I2(BRAM_L_X6Y140_RAMB18_X0Y56_DO19),
.I3(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO3),
.I4(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO3),
.I5(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO2),
.O5(CLBLM_R_X5Y138_SLICE_X7Y138_DO5),
.O6(CLBLM_R_X5Y138_SLICE_X7Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cc33cca5a55a5a)
  ) CLBLM_R_X5Y138_SLICE_X7Y138_CLUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y56_DO23),
.I1(CLBLM_R_X5Y126_SLICE_X7Y126_B5Q),
.I2(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO7),
.I3(CLBLM_R_X3Y142_SLICE_X2Y142_CQ),
.I4(CLBLM_R_X5Y138_SLICE_X7Y138_DO6),
.I5(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.O5(CLBLM_R_X5Y138_SLICE_X7Y138_CO5),
.O6(CLBLM_R_X5Y138_SLICE_X7Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X5Y138_SLICE_X7Y138_BLUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO3),
.I1(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO3),
.I2(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO2),
.I3(BRAM_L_X6Y140_RAMB18_X0Y56_DO18),
.I4(CLBLM_R_X5Y129_SLICE_X7Y129_AQ),
.I5(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO3),
.O5(CLBLM_R_X5Y138_SLICE_X7Y138_BO5),
.O6(CLBLM_R_X5Y138_SLICE_X7Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6666666666666666)
  ) CLBLM_R_X5Y138_SLICE_X7Y138_ALUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO6),
.I1(CLBLL_L_X4Y131_SLICE_X5Y131_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y138_SLICE_X7Y138_AO5),
.O6(CLBLM_R_X5Y138_SLICE_X7Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X5Y139_SLICE_X6Y139_DLUT (
.I0(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO7),
.I1(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO6),
.I2(BRAM_L_X6Y140_RAMB18_X0Y56_DO22),
.I3(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO7),
.I4(CLBLM_R_X5Y127_SLICE_X7Y127_DQ),
.I5(BRAM_L_X6Y140_RAMB18_X0Y56_DO23),
.O5(CLBLM_R_X5Y139_SLICE_X6Y139_DO5),
.O6(CLBLM_R_X5Y139_SLICE_X6Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X5Y139_SLICE_X6Y139_CLUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO1),
.I1(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO1),
.I2(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO0),
.I3(CLBLM_R_X5Y132_SLICE_X6Y132_B5Q),
.I4(BRAM_L_X6Y140_RAMB18_X0Y56_DO16),
.I5(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO1),
.O5(CLBLM_R_X5Y139_SLICE_X6Y139_CO5),
.O6(CLBLM_R_X5Y139_SLICE_X6Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X5Y139_SLICE_X6Y139_BLUT (
.I0(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I1(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO2),
.I2(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO2),
.I3(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO1),
.I4(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO2),
.I5(BRAM_L_X6Y140_RAMB18_X0Y56_DO17),
.O5(CLBLM_R_X5Y139_SLICE_X6Y139_BO5),
.O6(CLBLM_R_X5Y139_SLICE_X6Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X5Y139_SLICE_X6Y139_ALUT (
.I0(CLBLL_L_X4Y132_SLICE_X5Y132_BQ),
.I1(BRAM_L_X6Y140_RAMB18_X0Y56_DO22),
.I2(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO7),
.I3(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO7),
.I4(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO7),
.I5(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO6),
.O5(CLBLM_R_X5Y139_SLICE_X6Y139_AO5),
.O6(CLBLM_R_X5Y139_SLICE_X6Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3300ffccffcc3300)
  ) CLBLM_R_X5Y139_SLICE_X7Y139_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y139_SLICE_X7Y139_CO6),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_CQ),
.I5(CLBLM_R_X5Y127_SLICE_X7Y127_CQ),
.O5(CLBLM_R_X5Y139_SLICE_X7Y139_DO5),
.O6(CLBLM_R_X5Y139_SLICE_X7Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X5Y139_SLICE_X7Y139_CLUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y56_DO21),
.I1(CLBLM_R_X5Y127_SLICE_X7Y127_CQ),
.I2(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO6),
.I3(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO5),
.I4(BRAM_L_X6Y140_RAMB18_X0Y56_DO22),
.I5(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO6),
.O5(CLBLM_R_X5Y139_SLICE_X7Y139_CO5),
.O6(CLBLM_R_X5Y139_SLICE_X7Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X5Y139_SLICE_X7Y139_BLUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y56_DO6),
.I1(CLBLM_R_X3Y132_SLICE_X3Y132_CQ),
.I2(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO7),
.I3(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO7),
.I4(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO7),
.I5(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO6),
.O5(CLBLM_R_X5Y139_SLICE_X7Y139_BO5),
.O6(CLBLM_R_X5Y139_SLICE_X7Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555aaaac33cc33c)
  ) CLBLM_R_X5Y139_SLICE_X7Y139_ALUT (
.I0(CLBLM_R_X3Y149_SLICE_X2Y149_CQ),
.I1(CLBLM_R_X5Y138_SLICE_X7Y138_BO6),
.I2(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO7),
.I3(BRAM_L_X6Y140_RAMB18_X0Y56_DO23),
.I4(CLBLM_R_X5Y129_SLICE_X7Y129_AQ),
.I5(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.O5(CLBLM_R_X5Y139_SLICE_X7Y139_AO5),
.O6(CLBLM_R_X5Y139_SLICE_X7Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f50afa05f50afa0)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_DLUT (
.I0(CLBLM_R_X5Y127_SLICE_X7Y127_DQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I3(CLBLM_R_X5Y139_SLICE_X6Y139_DO6),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_DQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y140_SLICE_X6Y140_DO5),
.O6(CLBLM_R_X5Y140_SLICE_X6Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3a3a3a3acacacaca)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_CLUT (
.I0(CLBLM_R_X5Y139_SLICE_X6Y139_AO6),
.I1(CLBLL_L_X4Y132_SLICE_X5Y132_BQ),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X3Y151_SLICE_X2Y151_AQ),
.O5(CLBLM_R_X5Y140_SLICE_X6Y140_CO5),
.O6(CLBLM_R_X5Y140_SLICE_X6Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h22ee22eeee22ee22)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_BLUT (
.I0(CLBLM_R_X5Y139_SLICE_X6Y139_BO6),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y149_SLICE_X2Y149_BQ),
.O5(CLBLM_R_X5Y140_SLICE_X6Y140_BO5),
.O6(CLBLM_R_X5Y140_SLICE_X6Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5c53535caca3a3ac)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_ALUT (
.I0(CLBLM_R_X5Y132_SLICE_X6Y132_B5Q),
.I1(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO7),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I3(CLBLM_R_X5Y139_SLICE_X6Y139_CO6),
.I4(BRAM_L_X6Y140_RAMB18_X0Y56_DO23),
.I5(CLBLM_R_X3Y149_SLICE_X2Y149_AQ),
.O5(CLBLM_R_X5Y140_SLICE_X6Y140_AO5),
.O6(CLBLM_R_X5Y140_SLICE_X6Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y140_SLICE_X7Y140_DO5),
.O6(CLBLM_R_X5Y140_SLICE_X7Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y140_SLICE_X7Y140_CO5),
.O6(CLBLM_R_X5Y140_SLICE_X7Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y140_SLICE_X7Y140_BO5),
.O6(CLBLM_R_X5Y140_SLICE_X7Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff0cccc0ff0cccc)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y139_SLICE_X7Y139_BO6),
.I2(CLBLM_R_X3Y132_SLICE_X3Y132_CQ),
.I3(CLBLL_L_X2Y155_SLICE_X0Y155_DQ),
.I4(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y140_SLICE_X7Y140_AO5),
.O6(CLBLM_R_X5Y140_SLICE_X7Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y158_SLICE_X6Y158_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y229_IOB_X0Y230_I),
.Q(CLBLM_R_X5Y158_SLICE_X6Y158_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y158_SLICE_X6Y158_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y233_IOB_X0Y233_I),
.Q(CLBLM_R_X5Y158_SLICE_X6Y158_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y158_SLICE_X6Y158_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y239_IOB_X0Y239_I),
.Q(CLBLM_R_X5Y158_SLICE_X6Y158_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y158_SLICE_X6Y158_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(LIOB33_X0Y241_IOB_X0Y241_I),
.Q(CLBLM_R_X5Y158_SLICE_X6Y158_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y158_SLICE_X6Y158_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y158_SLICE_X6Y158_DO5),
.O6(CLBLM_R_X5Y158_SLICE_X6Y158_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y158_SLICE_X6Y158_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y158_SLICE_X6Y158_CO5),
.O6(CLBLM_R_X5Y158_SLICE_X6Y158_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y158_SLICE_X6Y158_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y158_SLICE_X6Y158_BO5),
.O6(CLBLM_R_X5Y158_SLICE_X6Y158_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y158_SLICE_X6Y158_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y158_SLICE_X6Y158_AO5),
.O6(CLBLM_R_X5Y158_SLICE_X6Y158_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y158_SLICE_X7Y158_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y158_SLICE_X7Y158_DO5),
.O6(CLBLM_R_X5Y158_SLICE_X7Y158_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y158_SLICE_X7Y158_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y158_SLICE_X7Y158_CO5),
.O6(CLBLM_R_X5Y158_SLICE_X7Y158_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y158_SLICE_X7Y158_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y158_SLICE_X7Y158_BO5),
.O6(CLBLM_R_X5Y158_SLICE_X7Y158_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y158_SLICE_X7Y158_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y158_SLICE_X7Y158_AO5),
.O6(CLBLM_R_X5Y158_SLICE_X7Y158_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X8Y125_BO5),
.Q(CLBLM_R_X7Y125_SLICE_X8Y125_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X8Y125_CO5),
.Q(CLBLM_R_X7Y125_SLICE_X8Y125_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X8Y125_AO6),
.Q(CLBLM_R_X7Y125_SLICE_X8Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X8Y125_BO6),
.Q(CLBLM_R_X7Y125_SLICE_X8Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X8Y125_CO6),
.Q(CLBLM_R_X7Y125_SLICE_X8Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff699600006996)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_DLUT (
.I0(BRAM_L_X6Y125_RAMB18_X0Y50_DO1),
.I1(CLBLM_R_X5Y125_SLICE_X7Y125_CQ),
.I2(CLBLM_R_X7Y125_SLICE_X9Y125_AQ),
.I3(CLBLM_R_X5Y125_SLICE_X7Y125_AO5),
.I4(LIOB33_X0Y147_IOB_X0Y148_I),
.I5(LIOB33_X0Y1_IOB_X0Y1_I),
.O5(CLBLM_R_X7Y125_SLICE_X8Y125_DO5),
.O6(CLBLM_R_X7Y125_SLICE_X8Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa55aad1d1e2e2)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_CLUT (
.I0(CLBLM_R_X7Y125_SLICE_X8Y125_C5Q),
.I1(LIOB33_X0Y147_IOB_X0Y148_I),
.I2(LIOB33_X0Y97_IOB_X0Y98_I),
.I3(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO2),
.I4(BRAM_L_X6Y125_RAMB18_X0Y50_DO2),
.I5(1'b1),
.O5(CLBLM_R_X7Y125_SLICE_X8Y125_CO5),
.O6(CLBLM_R_X7Y125_SLICE_X8Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa55aadede1212)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_BLUT (
.I0(CLBLM_R_X7Y125_SLICE_X8Y125_B5Q),
.I1(LIOB33_X0Y147_IOB_X0Y148_I),
.I2(BRAM_L_X6Y125_RAMB18_X0Y50_DO1),
.I3(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO1),
.I4(LIOB33_X0Y97_IOB_X0Y97_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y125_SLICE_X8Y125_BO5),
.O6(CLBLM_R_X7Y125_SLICE_X8Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cc33cc33cc33cc)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y125_SLICE_X7Y125_BQ),
.I2(1'b1),
.I3(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO2),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y125_SLICE_X8Y125_AO5),
.O6(CLBLM_R_X7Y125_SLICE_X8Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X8Y125_DO6),
.Q(CLBLM_R_X7Y125_SLICE_X9Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y125_SLICE_X7Y125_DO6),
.Q(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y125_SLICE_X9Y125_DO5),
.O6(CLBLM_R_X7Y125_SLICE_X9Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y125_SLICE_X9Y125_CO5),
.O6(CLBLM_R_X7Y125_SLICE_X9Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y125_SLICE_X9Y125_BO5),
.O6(CLBLM_R_X7Y125_SLICE_X9Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y125_SLICE_X9Y125_AO5),
.O6(CLBLM_R_X7Y125_SLICE_X9Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X8Y126_DO5),
.Q(CLBLM_R_X7Y126_SLICE_X8Y126_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X8Y126_AO6),
.Q(CLBLM_R_X7Y126_SLICE_X8Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X8Y126_BO6),
.Q(CLBLM_R_X7Y126_SLICE_X8Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X8Y126_CO6),
.Q(CLBLM_R_X7Y126_SLICE_X8Y126_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X8Y126_DO6),
.Q(CLBLM_R_X7Y126_SLICE_X8Y126_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffff008b8bb8b8)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_DLUT (
.I0(LIOB33_SING_X0Y99_IOB_X0Y99_I),
.I1(LIOB33_X0Y147_IOB_X0Y148_I),
.I2(BRAM_L_X6Y125_RAMB18_X0Y50_DO3),
.I3(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO3),
.I4(CLBLM_R_X7Y126_SLICE_X8Y126_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y126_SLICE_X8Y126_DO5),
.O6(CLBLM_R_X7Y126_SLICE_X8Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0ff0f0f0f0)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X5Y126_SLICE_X7Y126_B5Q),
.I3(1'b1),
.I4(1'b1),
.I5(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO3),
.O5(CLBLM_R_X7Y126_SLICE_X8Y126_CO5),
.O6(CLBLM_R_X7Y126_SLICE_X8Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333cccc3333cccc)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_BLUT (
.I0(1'b1),
.I1(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO2),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y126_SLICE_X8Y126_BO5),
.O6(CLBLM_R_X7Y126_SLICE_X8Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffff0000ffff00)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO1),
.I4(CLBLM_R_X7Y125_SLICE_X9Y125_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y126_SLICE_X8Y126_AO5),
.O6(CLBLM_R_X7Y126_SLICE_X8Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y126_SLICE_X7Y126_CO6),
.Q(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y126_SLICE_X9Y126_DO5),
.O6(CLBLM_R_X7Y126_SLICE_X9Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y126_SLICE_X9Y126_CO5),
.O6(CLBLM_R_X7Y126_SLICE_X9Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y126_SLICE_X9Y126_BO5),
.O6(CLBLM_R_X7Y126_SLICE_X9Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y126_SLICE_X9Y126_AO5),
.O6(CLBLM_R_X7Y126_SLICE_X9Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y127_SLICE_X8Y127_AO5),
.Q(CLBLM_R_X7Y127_SLICE_X8Y127_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y127_SLICE_X8Y127_AO6),
.Q(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y127_SLICE_X8Y127_DO5),
.O6(CLBLM_R_X7Y127_SLICE_X8Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y127_SLICE_X8Y127_CO5),
.O6(CLBLM_R_X7Y127_SLICE_X8Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y127_SLICE_X8Y127_BO5),
.O6(CLBLM_R_X7Y127_SLICE_X8Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h66666666ff3c003c)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_ALUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO0),
.I1(CLBLM_R_X7Y127_SLICE_X8Y127_A5Q),
.I2(BRAM_L_X6Y125_RAMB18_X0Y50_DO0),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(LIOB33_X0Y95_IOB_X0Y96_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y127_SLICE_X8Y127_AO5),
.O6(CLBLM_R_X7Y127_SLICE_X8Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y127_SLICE_X9Y127_DO5),
.O6(CLBLM_R_X7Y127_SLICE_X9Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y127_SLICE_X9Y127_CO5),
.O6(CLBLM_R_X7Y127_SLICE_X9Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y127_SLICE_X9Y127_BO5),
.O6(CLBLM_R_X7Y127_SLICE_X9Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y127_SLICE_X9Y127_AO5),
.O6(CLBLM_R_X7Y127_SLICE_X9Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X8Y128_AO5),
.Q(CLBLM_R_X7Y128_SLICE_X8Y128_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X8Y128_AO6),
.Q(CLBLM_R_X7Y128_SLICE_X8Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X8Y128_BO6),
.Q(CLBLM_R_X7Y128_SLICE_X8Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y128_SLICE_X8Y128_DO5),
.O6(CLBLM_R_X7Y128_SLICE_X8Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y128_SLICE_X8Y128_CO5),
.O6(CLBLM_R_X7Y128_SLICE_X8Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0ff0f00f0ff0f0)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO4),
.I3(1'b1),
.I4(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y128_SLICE_X8Y128_BO5),
.O6(CLBLM_R_X7Y128_SLICE_X8Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0ff0f088bbbb88)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_ALUT (
.I0(LIOB33_X0Y119_IOB_X0Y120_I),
.I1(LIOB33_X0Y147_IOB_X0Y148_I),
.I2(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO5),
.I3(BRAM_L_X6Y125_RAMB18_X0Y50_DO5),
.I4(CLBLM_R_X7Y128_SLICE_X8Y128_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y128_SLICE_X8Y128_AO5),
.O6(CLBLM_R_X7Y128_SLICE_X8Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X9Y128_AO6),
.Q(CLBLM_R_X7Y128_SLICE_X9Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y128_SLICE_X9Y128_DO5),
.O6(CLBLM_R_X7Y128_SLICE_X9Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y128_SLICE_X9Y128_CO5),
.O6(CLBLM_R_X7Y128_SLICE_X9Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y128_SLICE_X9Y128_BO5),
.O6(CLBLM_R_X7Y128_SLICE_X9Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff00ff00ff00ff0)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X5Y128_SLICE_X7Y128_AQ),
.I3(BRAM_L_X6Y135_RAMB18_X0Y54_DO16),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y128_SLICE_X9Y128_AO5),
.O6(CLBLM_R_X7Y128_SLICE_X9Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X8Y129_AO5),
.Q(CLBLM_R_X7Y129_SLICE_X8Y129_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X8Y129_BO5),
.Q(CLBLM_R_X7Y129_SLICE_X8Y129_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X8Y129_AO6),
.Q(CLBLM_R_X7Y129_SLICE_X8Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X8Y129_BO6),
.Q(CLBLM_R_X7Y129_SLICE_X8Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X8Y129_CO6),
.Q(CLBLM_R_X7Y129_SLICE_X8Y129_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X8Y129_DO6),
.Q(CLBLM_R_X7Y129_SLICE_X8Y129_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555555aaaaaaaa)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_DLUT (
.I0(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO2),
.O5(CLBLM_R_X7Y129_SLICE_X8Y129_DO5),
.O6(CLBLM_R_X7Y129_SLICE_X8Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555aaaa5555aaaa)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_CLUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X5Y129_SLICE_X7Y129_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X8Y129_CO5),
.O6(CLBLM_R_X7Y129_SLICE_X8Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ccccf066f066)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_BLUT (
.I0(BRAM_L_X6Y125_RAMB18_X0Y50_DO18),
.I1(CLBLM_R_X7Y129_SLICE_X8Y129_B5Q),
.I2(LIOB33_X0Y125_IOB_X0Y125_I),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(BRAM_L_X6Y135_RAMB18_X0Y54_DO2),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X8Y129_BO5),
.O6(CLBLM_R_X7Y129_SLICE_X8Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555aaaaf033f0cc)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_ALUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y54_DO0),
.I1(BRAM_L_X6Y125_RAMB18_X0Y50_DO16),
.I2(LIOB33_X0Y123_IOB_X0Y123_I),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(CLBLM_R_X7Y129_SLICE_X8Y129_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X8Y129_AO5),
.O6(CLBLM_R_X7Y129_SLICE_X8Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X9Y129_AO5),
.Q(CLBLM_R_X7Y129_SLICE_X9Y129_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X9Y129_BO5),
.Q(CLBLM_R_X7Y129_SLICE_X9Y129_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X9Y129_AO6),
.Q(CLBLM_R_X7Y129_SLICE_X9Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X9Y129_BO6),
.Q(CLBLM_R_X7Y129_SLICE_X9Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X9Y129_CO6),
.Q(CLBLM_R_X7Y129_SLICE_X9Y129_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X9Y129_DO5),
.O6(CLBLM_R_X7Y129_SLICE_X9Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0ff0f0f0f0)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X5Y127_SLICE_X7Y127_B5Q),
.I3(1'b1),
.I4(1'b1),
.I5(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO5),
.O5(CLBLM_R_X7Y129_SLICE_X9Y129_CO5),
.O6(CLBLM_R_X7Y129_SLICE_X9Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa55aad1d1e2e2)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_BLUT (
.I0(CLBLM_R_X7Y129_SLICE_X9Y129_B5Q),
.I1(LIOB33_X0Y147_IOB_X0Y148_I),
.I2(LIOB33_X0Y121_IOB_X0Y121_I),
.I3(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO6),
.I4(BRAM_L_X6Y125_RAMB18_X0Y50_DO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X9Y129_BO5),
.O6(CLBLM_R_X7Y129_SLICE_X9Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0ff0f08bb88bb8)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_ALUT (
.I0(LIOB33_X0Y119_IOB_X0Y119_I),
.I1(LIOB33_X0Y147_IOB_X0Y148_I),
.I2(CLBLM_R_X7Y129_SLICE_X9Y129_A5Q),
.I3(BRAM_L_X6Y125_RAMB18_X0Y50_DO4),
.I4(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO4),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X9Y129_AO5),
.O6(CLBLM_R_X7Y129_SLICE_X9Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y130_SLICE_X5Y130_BO6),
.Q(CLBLM_R_X7Y130_SLICE_X8Y130_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y129_SLICE_X5Y129_DO6),
.Q(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X8Y130_BO6),
.Q(CLBLM_R_X7Y130_SLICE_X8Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f50afa05f50afa0)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_DLUT (
.I0(CLBLM_R_X5Y125_SLICE_X7Y125_BQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I3(CLBLM_R_X7Y130_SLICE_X8Y130_CO6),
.I4(CLBLL_L_X4Y156_SLICE_X4Y156_CQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y130_SLICE_X8Y130_DO5),
.O6(CLBLM_R_X7Y130_SLICE_X8Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_CLUT (
.I0(CLBLM_R_X5Y125_SLICE_X7Y125_BQ),
.I1(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO2),
.I2(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO1),
.I3(BRAM_R_X17Y135_RAMB18_X1Y54_DO17),
.I4(BRAM_L_X6Y135_RAMB18_X0Y54_DO18),
.I5(BRAM_R_X17Y135_RAMB18_X1Y54_DO18),
.O5(CLBLM_R_X7Y130_SLICE_X8Y130_CO5),
.O6(CLBLM_R_X7Y130_SLICE_X8Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555555aaaaaaaa)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_BLUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO0),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y130_SLICE_X7Y130_CQ),
.O5(CLBLM_R_X7Y130_SLICE_X8Y130_BO5),
.O6(CLBLM_R_X7Y130_SLICE_X8Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffff000ff00ff0)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X4Y128_SLICE_X5Y128_AQ),
.I3(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO7),
.I4(BRAM_L_X6Y135_RAMB18_X0Y54_DO23),
.I5(1'b1),
.O5(CLBLM_R_X7Y130_SLICE_X8Y130_AO5),
.O6(CLBLM_R_X7Y130_SLICE_X8Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X9Y130_AO6),
.Q(CLBLM_R_X7Y130_SLICE_X9Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X9Y130_BO6),
.Q(CLBLM_R_X7Y130_SLICE_X9Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X9Y130_CO6),
.Q(CLBLM_R_X7Y130_SLICE_X9Y130_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X9Y130_DO6),
.Q(CLBLM_R_X7Y130_SLICE_X9Y130_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5a5a5a5a5a)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_DLUT (
.I0(CLBLL_L_X4Y129_SLICE_X5Y129_AQ),
.I1(1'b1),
.I2(BRAM_L_X6Y135_RAMB18_X0Y54_DO18),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y130_SLICE_X9Y130_DO5),
.O6(CLBLM_R_X7Y130_SLICE_X9Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cc33cc33cc33cc)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_CLUT (
.I0(1'b1),
.I1(BRAM_L_X6Y140_RAMB18_X0Y56_DO18),
.I2(1'b1),
.I3(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y130_SLICE_X9Y130_CO5),
.O6(CLBLM_R_X7Y130_SLICE_X9Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cc33cc33cc33cc)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_BLUT (
.I0(1'b1),
.I1(BRAM_L_X6Y140_RAMB18_X0Y56_DO16),
.I2(1'b1),
.I3(CLBLM_R_X5Y130_SLICE_X7Y130_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y130_SLICE_X9Y130_BO5),
.O6(CLBLM_R_X7Y130_SLICE_X9Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffff0000ffff00)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X5Y129_SLICE_X6Y129_A5Q),
.I4(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO3),
.I5(1'b1),
.O5(CLBLM_R_X7Y130_SLICE_X9Y130_AO5),
.O6(CLBLM_R_X7Y130_SLICE_X9Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5c53aca3535ca3ac)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_DLUT (
.I0(CLBLL_L_X4Y156_SLICE_X4Y156_BQ),
.I1(BRAM_R_X17Y135_RAMB18_X1Y54_DO23),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I3(CLBLM_L_X8Y131_SLICE_X10Y131_DO6),
.I4(CLBLM_R_X5Y125_SLICE_X7Y125_AQ),
.I5(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO7),
.O5(CLBLM_R_X7Y131_SLICE_X8Y131_DO5),
.O6(CLBLM_R_X7Y131_SLICE_X8Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h09f9f90906f6f606)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_CLUT (
.I0(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO7),
.I1(BRAM_R_X17Y135_RAMB18_X1Y54_DO23),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I3(CLBLM_R_X5Y126_SLICE_X6Y126_AQ),
.I4(CLBLL_L_X4Y156_SLICE_X4Y156_DQ),
.I5(CLBLM_L_X8Y131_SLICE_X10Y131_CO6),
.O5(CLBLM_R_X7Y131_SLICE_X8Y131_CO5),
.O6(CLBLM_R_X7Y131_SLICE_X8Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_BLUT (
.I0(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO1),
.I1(CLBLL_L_X4Y129_SLICE_X4Y129_AQ),
.I2(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO1),
.I3(BRAM_L_X6Y135_RAMB18_X0Y54_DO16),
.I4(BRAM_R_X17Y135_RAMB18_X1Y54_DO17),
.I5(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO0),
.O5(CLBLM_R_X7Y131_SLICE_X8Y131_BO5),
.O6(CLBLM_R_X7Y131_SLICE_X8Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h1eb44be14be11eb4)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_ALUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I1(CLBLM_R_X7Y130_SLICE_X8Y130_AO6),
.I2(CLBLM_R_X5Y128_SLICE_X7Y128_AQ),
.I3(CLBLM_R_X3Y155_SLICE_X2Y155_AQ),
.I4(CLBLM_L_X8Y130_SLICE_X11Y130_AO6),
.I5(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO0),
.O5(CLBLM_R_X7Y131_SLICE_X8Y131_AO5),
.O6(CLBLM_R_X7Y131_SLICE_X8Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X9Y131_AO5),
.Q(CLBLM_R_X7Y131_SLICE_X9Y131_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X9Y131_AO6),
.Q(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X9Y131_BO6),
.Q(CLBLM_R_X7Y131_SLICE_X9Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X9Y131_CO6),
.Q(CLBLM_R_X7Y131_SLICE_X9Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X9Y131_DO6),
.Q(CLBLM_R_X7Y131_SLICE_X9Y131_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6666666666666666)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_DLUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO6),
.I1(CLBLM_R_X5Y130_SLICE_X6Y130_B5Q),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y131_SLICE_X9Y131_DO5),
.O6(CLBLM_R_X7Y131_SLICE_X9Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cc33cc33cc33cc)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_CLUT (
.I0(1'b1),
.I1(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO5),
.I2(1'b1),
.I3(CLBLL_L_X4Y130_SLICE_X5Y130_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y131_SLICE_X9Y131_CO5),
.O6(CLBLM_R_X7Y131_SLICE_X9Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333cccc3333cccc)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y130_SLICE_X7Y130_A5Q),
.I2(1'b1),
.I3(1'b1),
.I4(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO4),
.I5(1'b1),
.O5(CLBLM_R_X7Y131_SLICE_X9Y131_BO5),
.O6(CLBLM_R_X7Y131_SLICE_X9Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555aaaaf033f0cc)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_ALUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y54_DO5),
.I1(BRAM_L_X6Y125_RAMB18_X0Y50_DO21),
.I2(LIOB33_X0Y129_IOB_X0Y129_I),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(CLBLM_R_X7Y131_SLICE_X9Y131_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y131_SLICE_X9Y131_AO5),
.O6(CLBLM_R_X7Y131_SLICE_X9Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y132_SLICE_X8Y132_AO5),
.Q(CLBLM_R_X7Y132_SLICE_X8Y132_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y132_SLICE_X8Y132_AO6),
.Q(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y132_SLICE_X6Y132_DO6),
.Q(CLBLM_R_X7Y132_SLICE_X8Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y132_SLICE_X6Y132_CO6),
.Q(CLBLM_R_X7Y132_SLICE_X8Y132_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555f0f0aaaaf0f0)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_DLUT (
.I0(CLBLM_R_X3Y158_SLICE_X3Y158_AQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y132_SLICE_X9Y132_DO6),
.I3(1'b1),
.I4(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I5(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.O5(CLBLM_R_X7Y132_SLICE_X8Y132_DO5),
.O6(CLBLM_R_X7Y132_SLICE_X8Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f9966f0f09966)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_CLUT (
.I0(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO7),
.I1(CLBLM_R_X7Y132_SLICE_X9Y132_CO6),
.I2(CLBLM_R_X5Y126_SLICE_X7Y126_AQ),
.I3(BRAM_R_X17Y135_RAMB18_X1Y54_DO23),
.I4(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I5(CLBLM_R_X3Y158_SLICE_X3Y158_BQ),
.O5(CLBLM_R_X7Y132_SLICE_X8Y132_CO5),
.O6(CLBLM_R_X7Y132_SLICE_X8Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h72d8278d278d72d8)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_BLUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I1(CLBLL_L_X4Y129_SLICE_X4Y129_AQ),
.I2(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO7),
.I3(CLBLM_R_X3Y158_SLICE_X3Y158_CQ),
.I4(CLBLM_R_X7Y131_SLICE_X8Y131_BO6),
.I5(BRAM_L_X6Y135_RAMB18_X0Y54_DO23),
.O5(CLBLM_R_X7Y132_SLICE_X8Y132_BO5),
.O6(CLBLM_R_X7Y132_SLICE_X8Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3cbbee1144)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_ALUT (
.I0(LIOB33_X0Y147_IOB_X0Y148_I),
.I1(CLBLM_R_X7Y132_SLICE_X8Y132_A5Q),
.I2(BRAM_L_X6Y135_RAMB18_X0Y54_DO4),
.I3(BRAM_L_X6Y125_RAMB18_X0Y50_DO20),
.I4(LIOB33_X0Y127_IOB_X0Y127_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y132_SLICE_X8Y132_AO5),
.O6(CLBLM_R_X7Y132_SLICE_X8Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y132_SLICE_X9Y132_AO6),
.Q(CLBLM_R_X7Y132_SLICE_X9Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_DLUT (
.I0(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO7),
.I1(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO0),
.I2(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.I3(BRAM_L_X6Y135_RAMB18_X0Y54_DO16),
.I4(BRAM_R_X17Y135_RAMB18_X1Y54_DO23),
.I5(BRAM_R_X17Y135_RAMB18_X1Y54_DO16),
.O5(CLBLM_R_X7Y132_SLICE_X9Y132_DO5),
.O6(CLBLM_R_X7Y132_SLICE_X9Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_CLUT (
.I0(BRAM_R_X17Y135_RAMB18_X1Y54_DO20),
.I1(BRAM_L_X6Y135_RAMB18_X0Y54_DO20),
.I2(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO3),
.I3(BRAM_R_X17Y135_RAMB18_X1Y54_DO19),
.I4(CLBLM_R_X5Y126_SLICE_X7Y126_AQ),
.I5(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO4),
.O5(CLBLM_R_X7Y132_SLICE_X9Y132_CO5),
.O6(CLBLM_R_X7Y132_SLICE_X9Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_BLUT (
.I0(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO2),
.I1(BRAM_R_X17Y135_RAMB18_X1Y54_DO18),
.I2(CLBLL_L_X4Y129_SLICE_X5Y129_AQ),
.I3(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO2),
.I4(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO1),
.I5(BRAM_L_X6Y135_RAMB18_X0Y54_DO17),
.O5(CLBLM_R_X7Y132_SLICE_X9Y132_BO5),
.O6(CLBLM_R_X7Y132_SLICE_X9Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5a5a5a5a5a)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_ALUT (
.I0(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO6),
.I1(1'b1),
.I2(CLBLL_L_X4Y133_SLICE_X4Y133_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y132_SLICE_X9Y132_AO5),
.O6(CLBLM_R_X7Y132_SLICE_X9Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h74747474b8b8b8b8)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_DLUT (
.I0(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I2(CLBLM_R_X7Y133_SLICE_X9Y133_DO6),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X2Y157_SLICE_X0Y157_DQ),
.O5(CLBLM_R_X7Y133_SLICE_X8Y133_DO5),
.O6(CLBLM_R_X7Y133_SLICE_X8Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f99f0990f66f066)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_CLUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y54_DO23),
.I1(CLBLM_R_X7Y133_SLICE_X9Y133_CO6),
.I2(CLBLM_R_X5Y128_SLICE_X6Y128_AQ),
.I3(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I4(CLBLM_R_X3Y155_SLICE_X2Y155_BQ),
.I5(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO7),
.O5(CLBLM_R_X7Y133_SLICE_X8Y133_CO5),
.O6(CLBLM_R_X7Y133_SLICE_X8Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_BLUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO3),
.I1(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO2),
.I2(BRAM_L_X6Y140_RAMB18_X0Y56_DO19),
.I3(CLBLM_R_X7Y132_SLICE_X8Y132_BQ),
.I4(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO2),
.I5(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO3),
.O5(CLBLM_R_X7Y133_SLICE_X8Y133_BO5),
.O6(CLBLM_R_X7Y133_SLICE_X8Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3caa553c3c55aa)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_ALUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO7),
.I1(CLBLM_R_X7Y132_SLICE_X8Y132_BQ),
.I2(CLBLL_L_X4Y146_SLICE_X4Y146_AQ),
.I3(CLBLM_R_X7Y133_SLICE_X8Y133_BO6),
.I4(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I5(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO7),
.O5(CLBLM_R_X7Y133_SLICE_X8Y133_AO5),
.O6(CLBLM_R_X7Y133_SLICE_X8Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X9Y133_AO6),
.Q(CLBLM_R_X7Y133_SLICE_X9Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X9Y133_BO6),
.Q(CLBLM_R_X7Y133_SLICE_X9Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_DLUT (
.I0(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO4),
.I1(BRAM_R_X17Y135_RAMB18_X1Y54_DO21),
.I2(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO5),
.I3(BRAM_R_X17Y135_RAMB18_X1Y54_DO20),
.I4(BRAM_L_X6Y135_RAMB18_X0Y54_DO21),
.I5(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.O5(CLBLM_R_X7Y133_SLICE_X9Y133_DO5),
.O6(CLBLM_R_X7Y133_SLICE_X9Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_CLUT (
.I0(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO2),
.I1(BRAM_R_X17Y135_RAMB18_X1Y54_DO19),
.I2(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO3),
.I3(BRAM_L_X6Y135_RAMB18_X0Y54_DO18),
.I4(CLBLM_R_X5Y128_SLICE_X6Y128_AQ),
.I5(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO3),
.O5(CLBLM_R_X7Y133_SLICE_X9Y133_CO5),
.O6(CLBLM_R_X7Y133_SLICE_X9Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0ff0f0f0f0)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y125_SLICE_X7Y125_CQ),
.O5(CLBLM_R_X7Y133_SLICE_X9Y133_BO5),
.O6(CLBLM_R_X7Y133_SLICE_X9Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa55aa55aa55aa)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_ALUT (
.I0(CLBLL_L_X4Y133_SLICE_X4Y133_A5Q),
.I1(1'b1),
.I2(1'b1),
.I3(BRAM_L_X6Y140_RAMB18_X0Y56_DO21),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y133_SLICE_X9Y133_AO5),
.O6(CLBLM_R_X7Y133_SLICE_X9Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aacccc55aacccc)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_DLUT (
.I0(CLBLM_R_X7Y125_SLICE_X8Y125_C5Q),
.I1(CLBLM_L_X8Y134_SLICE_X10Y134_DO6),
.I2(1'b1),
.I3(CLBLM_R_X3Y157_SLICE_X2Y157_CQ),
.I4(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y134_SLICE_X8Y134_DO5),
.O6(CLBLM_R_X7Y134_SLICE_X8Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff9696ff009696)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_CLUT (
.I0(BRAM_R_X17Y135_RAMB18_X1Y54_DO7),
.I1(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO7),
.I2(CLBLM_R_X7Y134_SLICE_X9Y134_DO6),
.I3(CLBLM_R_X7Y126_SLICE_X8Y126_D5Q),
.I4(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I5(CLBLM_R_X3Y157_SLICE_X2Y157_DQ),
.O5(CLBLM_R_X7Y134_SLICE_X8Y134_CO5),
.O6(CLBLM_R_X7Y134_SLICE_X8Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_BLUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y54_DO20),
.I1(BRAM_R_X17Y135_RAMB18_X1Y54_DO21),
.I2(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO5),
.I3(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO5),
.I4(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO4),
.I5(CLBLM_R_X3Y130_SLICE_X3Y130_AQ),
.O5(CLBLM_R_X7Y134_SLICE_X8Y134_BO5),
.O6(CLBLM_R_X7Y134_SLICE_X8Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_ALUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y56_DO21),
.I1(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO5),
.I2(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO4),
.I3(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO5),
.I4(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO4),
.I5(CLBLM_R_X7Y132_SLICE_X8Y132_CQ),
.O5(CLBLM_R_X7Y134_SLICE_X8Y134_AO5),
.O6(CLBLM_R_X7Y134_SLICE_X8Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X9Y134_AO5),
.Q(CLBLM_R_X7Y134_SLICE_X9Y134_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X9Y134_BO5),
.Q(CLBLM_R_X7Y134_SLICE_X9Y134_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X9Y134_AO6),
.Q(CLBLM_R_X7Y134_SLICE_X9Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X9Y134_BO6),
.Q(CLBLM_R_X7Y134_SLICE_X9Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_DLUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y54_DO3),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_D5Q),
.I2(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO2),
.I3(BRAM_R_X17Y135_RAMB18_X1Y54_DO2),
.I4(BRAM_R_X17Y135_RAMB18_X1Y54_DO3),
.I5(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO3),
.O5(CLBLM_R_X7Y134_SLICE_X9Y134_DO5),
.O6(CLBLM_R_X7Y134_SLICE_X9Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_CLUT (
.I0(CLBLL_L_X4Y131_SLICE_X5Y131_AQ),
.I1(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO3),
.I2(BRAM_L_X6Y135_RAMB18_X0Y54_DO19),
.I3(BRAM_R_X17Y135_RAMB18_X1Y54_DO20),
.I4(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO4),
.I5(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO4),
.O5(CLBLM_R_X7Y134_SLICE_X9Y134_CO5),
.O6(CLBLM_R_X7Y134_SLICE_X9Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa55aadede1212)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_BLUT (
.I0(CLBLM_R_X7Y134_SLICE_X9Y134_B5Q),
.I1(LIOB33_X0Y147_IOB_X0Y148_I),
.I2(BRAM_L_X6Y130_RAMB18_X0Y52_DO3),
.I3(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO3),
.I4(LIOB33_X0Y135_IOB_X0Y135_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y134_SLICE_X9Y134_BO5),
.O6(CLBLM_R_X7Y134_SLICE_X9Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ccccf055f0aa)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_ALUT (
.I0(BRAM_L_X6Y130_RAMB18_X0Y52_DO2),
.I1(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO2),
.I2(LIOB33_X0Y133_IOB_X0Y134_I),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(CLBLM_R_X7Y134_SLICE_X9Y134_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y134_SLICE_X9Y134_AO5),
.O6(CLBLM_R_X7Y134_SLICE_X9Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7474b8b87474b8b8)
  ) CLBLM_R_X7Y135_SLICE_X8Y135_DLUT (
.I0(CLBLM_R_X3Y158_SLICE_X3Y158_DQ),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I2(CLBLM_R_X7Y132_SLICE_X9Y132_BO6),
.I3(1'b1),
.I4(CLBLL_L_X4Y129_SLICE_X5Y129_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y135_SLICE_X8Y135_DO5),
.O6(CLBLM_R_X7Y135_SLICE_X8Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7b7b7b7b48484848)
  ) CLBLM_R_X7Y135_SLICE_X8Y135_CLUT (
.I0(CLBLM_R_X3Y130_SLICE_X3Y130_AQ),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I2(CLBLM_R_X3Y157_SLICE_X2Y157_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X7Y134_SLICE_X8Y134_BO6),
.O5(CLBLM_R_X7Y135_SLICE_X8Y135_CO5),
.O6(CLBLM_R_X7Y135_SLICE_X8Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4ee41bb11bb14ee4)
  ) CLBLM_R_X7Y135_SLICE_X8Y135_BLUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I1(CLBLM_R_X7Y134_SLICE_X9Y134_CO6),
.I2(CLBLL_L_X4Y131_SLICE_X5Y131_AQ),
.I3(CLBLM_R_X3Y158_SLICE_X2Y158_AQ),
.I4(BRAM_L_X6Y135_RAMB18_X0Y54_DO23),
.I5(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO7),
.O5(CLBLM_R_X7Y135_SLICE_X8Y135_BO5),
.O6(CLBLM_R_X7Y135_SLICE_X8Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4114ebbeebbe4114)
  ) CLBLM_R_X7Y135_SLICE_X8Y135_ALUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I1(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO7),
.I2(CLBLM_R_X7Y135_SLICE_X9Y135_CO6),
.I3(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO7),
.I4(CLBLM_R_X3Y147_SLICE_X2Y147_AQ),
.I5(CLBLM_R_X5Y131_SLICE_X6Y131_A5Q),
.O5(CLBLM_R_X7Y135_SLICE_X8Y135_AO5),
.O6(CLBLM_R_X7Y135_SLICE_X8Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3caa3caa3caa3caa)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_DLUT (
.I0(CLBLM_R_X7Y135_SLICE_X9Y135_AO6),
.I1(CLBLM_R_X3Y132_SLICE_X2Y132_DQ),
.I2(CLBLL_L_X4Y156_SLICE_X5Y156_CQ),
.I3(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y135_SLICE_X9Y135_DO5),
.O6(CLBLM_R_X7Y135_SLICE_X9Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_CLUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO4),
.I1(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO3),
.I2(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO4),
.I3(CLBLM_R_X5Y131_SLICE_X6Y131_A5Q),
.I4(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO3),
.I5(BRAM_L_X6Y140_RAMB18_X0Y56_DO20),
.O5(CLBLM_R_X7Y135_SLICE_X9Y135_CO5),
.O6(CLBLM_R_X7Y135_SLICE_X9Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_BLUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y54_DO22),
.I1(CLBLL_L_X4Y133_SLICE_X5Y133_AQ),
.I2(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO7),
.I3(BRAM_R_X17Y135_RAMB18_X1Y54_DO23),
.I4(BRAM_L_X6Y135_RAMB18_X0Y54_DO23),
.I5(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO6),
.O5(CLBLM_R_X7Y135_SLICE_X9Y135_BO5),
.O6(CLBLM_R_X7Y135_SLICE_X9Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_ALUT (
.I0(BRAM_R_X17Y135_RAMB18_X1Y54_DO22),
.I1(CLBLM_R_X3Y132_SLICE_X2Y132_DQ),
.I2(BRAM_L_X6Y135_RAMB18_X0Y54_DO23),
.I3(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO7),
.I4(BRAM_L_X6Y125_RAMB18_X0Y51_DOADO7),
.I5(BRAM_L_X6Y130_RAMB18_X0Y53_DOADO6),
.O5(CLBLM_R_X7Y135_SLICE_X9Y135_AO5),
.O6(CLBLM_R_X7Y135_SLICE_X9Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y136_SLICE_X8Y136_AO5),
.Q(CLBLM_R_X7Y136_SLICE_X8Y136_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y136_SLICE_X8Y136_AO6),
.Q(CLBLM_R_X7Y136_SLICE_X8Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y136_SLICE_X8Y136_BO6),
.Q(CLBLM_R_X7Y136_SLICE_X8Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5050fafafafa5050)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_DLUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y136_SLICE_X9Y136_BO6),
.I3(1'b1),
.I4(CLBLL_L_X4Y156_SLICE_X5Y156_DQ),
.I5(CLBLM_R_X7Y127_SLICE_X8Y127_A5Q),
.O5(CLBLM_R_X7Y136_SLICE_X8Y136_DO5),
.O6(CLBLM_R_X7Y136_SLICE_X8Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4114ebbeebbe4114)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_CLUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I1(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO7),
.I2(CLBLM_L_X8Y136_SLICE_X10Y136_DO6),
.I3(BRAM_R_X17Y135_RAMB18_X1Y54_DO7),
.I4(CLBLM_R_X7Y125_SLICE_X8Y125_B5Q),
.I5(CLBLL_L_X4Y156_SLICE_X5Y156_A5Q),
.O5(CLBLM_R_X7Y136_SLICE_X8Y136_CO5),
.O6(CLBLM_R_X7Y136_SLICE_X8Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333333cccccccc)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_BLUT (
.I0(1'b1),
.I1(BRAM_L_X6Y140_RAMB18_X0Y56_DO4),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X3Y133_SLICE_X3Y133_BQ),
.O5(CLBLM_R_X7Y136_SLICE_X8Y136_BO5),
.O6(CLBLM_R_X7Y136_SLICE_X8Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffff00d1d1e2e2)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_ALUT (
.I0(BRAM_L_X6Y125_RAMB18_X0Y50_DO17),
.I1(LIOB33_X0Y147_IOB_X0Y148_I),
.I2(LIOB33_X0Y123_IOB_X0Y124_I),
.I3(BRAM_L_X6Y135_RAMB18_X0Y54_DO1),
.I4(CLBLM_R_X7Y136_SLICE_X8Y136_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y136_SLICE_X8Y136_AO5),
.O6(CLBLM_R_X7Y136_SLICE_X8Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f303f30cfc0cfc0)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y129_SLICE_X8Y129_B5Q),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I3(CLBLM_R_X7Y136_SLICE_X9Y136_AO6),
.I4(1'b1),
.I5(CLBLM_R_X25Y151_SLICE_X36Y151_AQ),
.O5(CLBLM_R_X7Y136_SLICE_X9Y136_DO5),
.O6(CLBLM_R_X7Y136_SLICE_X9Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7d7d7d7d28282828)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_CLUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I1(CLBLL_L_X4Y156_SLICE_X5Y156_AQ),
.I2(CLBLL_L_X4Y133_SLICE_X5Y133_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X7Y135_SLICE_X9Y135_BO6),
.O5(CLBLM_R_X7Y136_SLICE_X9Y136_CO5),
.O6(CLBLM_R_X7Y136_SLICE_X9Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_BLUT (
.I0(BRAM_R_X17Y135_RAMB18_X1Y54_DO0),
.I1(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO0),
.I2(BRAM_L_X6Y135_RAMB18_X0Y54_DO0),
.I3(CLBLM_R_X7Y127_SLICE_X8Y127_A5Q),
.I4(BRAM_R_X17Y135_RAMB18_X1Y54_DO7),
.I5(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO7),
.O5(CLBLM_R_X7Y136_SLICE_X9Y136_BO5),
.O6(CLBLM_R_X7Y136_SLICE_X9Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_ALUT (
.I0(BRAM_R_X17Y135_RAMB18_X1Y54_DO2),
.I1(CLBLM_R_X7Y129_SLICE_X8Y129_B5Q),
.I2(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO2),
.I3(BRAM_L_X6Y135_RAMB18_X0Y54_DO1),
.I4(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO1),
.I5(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO2),
.O5(CLBLM_R_X7Y136_SLICE_X9Y136_AO5),
.O6(CLBLM_R_X7Y136_SLICE_X9Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y137_SLICE_X8Y137_AO5),
.Q(CLBLM_R_X7Y137_SLICE_X8Y137_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y137_SLICE_X8Y137_AO6),
.Q(CLBLM_R_X7Y137_SLICE_X8Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y137_SLICE_X8Y137_BO6),
.Q(CLBLM_R_X7Y137_SLICE_X8Y137_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f0a5f0af5a0f5a0)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_DLUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I1(1'b1),
.I2(CLBLM_R_X3Y147_SLICE_X3Y147_BQ),
.I3(CLBLM_R_X7Y137_SLICE_X8Y137_CO6),
.I4(1'b1),
.I5(CLBLL_L_X4Y130_SLICE_X5Y130_A5Q),
.O5(CLBLM_R_X7Y137_SLICE_X8Y137_DO5),
.O6(CLBLM_R_X7Y137_SLICE_X8Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_CLUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO4),
.I1(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO4),
.I2(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO5),
.I3(CLBLL_L_X4Y130_SLICE_X5Y130_A5Q),
.I4(BRAM_L_X6Y140_RAMB18_X0Y56_DO21),
.I5(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO5),
.O5(CLBLM_R_X7Y137_SLICE_X8Y137_CO5),
.O6(CLBLM_R_X7Y137_SLICE_X8Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0ff0f0f0f0)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO6),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X4Y127_SLICE_X5Y127_AQ),
.O5(CLBLM_R_X7Y137_SLICE_X8Y137_BO5),
.O6(CLBLM_R_X7Y137_SLICE_X8Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3caaaa33cc)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_ALUT (
.I0(LIOB33_X0Y129_IOB_X0Y130_I),
.I1(CLBLM_R_X7Y137_SLICE_X8Y137_A5Q),
.I2(BRAM_L_X6Y135_RAMB18_X0Y54_DO6),
.I3(BRAM_L_X6Y125_RAMB18_X0Y50_DO22),
.I4(LIOB33_X0Y147_IOB_X0Y148_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y137_SLICE_X8Y137_AO5),
.O6(CLBLM_R_X7Y137_SLICE_X8Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y137_SLICE_X9Y137_AO6),
.Q(CLBLM_R_X7Y137_SLICE_X9Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y137_SLICE_X9Y137_BO6),
.Q(CLBLM_R_X7Y137_SLICE_X9Y137_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y137_SLICE_X9Y137_CO6),
.Q(CLBLM_R_X7Y137_SLICE_X9Y137_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y137_SLICE_X9Y137_DO6),
.Q(CLBLM_R_X7Y137_SLICE_X9Y137_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6666666666666666)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_DLUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y56_DO7),
.I1(CLBLM_R_X3Y132_SLICE_X3Y132_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y137_SLICE_X9Y137_DO5),
.O6(CLBLM_R_X7Y137_SLICE_X9Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3c3c3c3c3c)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_CLUT (
.I0(1'b1),
.I1(BRAM_L_X6Y140_RAMB18_X0Y56_DO1),
.I2(CLBLL_L_X4Y132_SLICE_X4Y132_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y137_SLICE_X9Y137_CO5),
.O6(CLBLM_R_X7Y137_SLICE_X9Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3c3c3c3c3c)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y131_SLICE_X6Y131_CQ),
.I2(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO0),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y137_SLICE_X9Y137_BO5),
.O6(CLBLM_R_X7Y137_SLICE_X9Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ffff00ff00)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X5Y126_SLICE_X6Y126_BQ),
.I4(1'b1),
.I5(BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO3),
.O5(CLBLM_R_X7Y137_SLICE_X9Y137_AO5),
.O6(CLBLM_R_X7Y137_SLICE_X9Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f0a5f0af5a0f5a0)
  ) CLBLM_R_X7Y138_SLICE_X8Y138_DLUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I1(1'b1),
.I2(CLBLM_R_X3Y145_SLICE_X2Y145_BQ),
.I3(CLBLM_R_X7Y138_SLICE_X8Y138_CO6),
.I4(1'b1),
.I5(CLBLM_R_X5Y127_SLICE_X7Y127_B5Q),
.O5(CLBLM_R_X7Y138_SLICE_X8Y138_DO5),
.O6(CLBLM_R_X7Y138_SLICE_X8Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X7Y138_SLICE_X8Y138_CLUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO4),
.I1(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO5),
.I2(BRAM_L_X6Y140_RAMB18_X0Y56_DO21),
.I3(CLBLM_R_X5Y127_SLICE_X7Y127_B5Q),
.I4(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO5),
.I5(BRAM_L_X6Y140_RAMB18_X0Y56_DO20),
.O5(CLBLM_R_X7Y138_SLICE_X8Y138_CO5),
.O6(CLBLM_R_X7Y138_SLICE_X8Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X7Y138_SLICE_X8Y138_BLUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO3),
.I1(BRAM_L_X6Y140_RAMB18_X0Y56_DO20),
.I2(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO4),
.I3(CLBLM_R_X5Y130_SLICE_X7Y130_A5Q),
.I4(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO4),
.I5(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO3),
.O5(CLBLM_R_X7Y138_SLICE_X8Y138_BO5),
.O6(CLBLM_R_X7Y138_SLICE_X8Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f9966f0f09966)
  ) CLBLM_R_X7Y138_SLICE_X8Y138_ALUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO7),
.I1(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO7),
.I2(CLBLM_R_X3Y147_SLICE_X3Y147_AQ),
.I3(CLBLM_R_X7Y138_SLICE_X8Y138_BO6),
.I4(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I5(CLBLM_R_X5Y130_SLICE_X7Y130_A5Q),
.O5(CLBLM_R_X7Y138_SLICE_X8Y138_AO5),
.O6(CLBLM_R_X7Y138_SLICE_X8Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y138_SLICE_X9Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y138_SLICE_X9Y138_AO6),
.Q(CLBLM_R_X7Y138_SLICE_X9Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y138_SLICE_X9Y138_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y138_SLICE_X9Y138_BO6),
.Q(CLBLM_R_X7Y138_SLICE_X9Y138_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y138_SLICE_X9Y138_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y138_SLICE_X9Y138_CO6),
.Q(CLBLM_R_X7Y138_SLICE_X9Y138_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y138_SLICE_X9Y138_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y138_SLICE_X9Y138_DO6),
.Q(CLBLM_R_X7Y138_SLICE_X9Y138_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6666666666666666)
  ) CLBLM_R_X7Y138_SLICE_X9Y138_DLUT (
.I0(CLBLL_L_X4Y130_SLICE_X4Y130_BQ),
.I1(BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y138_SLICE_X9Y138_DO5),
.O6(CLBLM_R_X7Y138_SLICE_X9Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cc33cc33cc33cc)
  ) CLBLM_R_X7Y138_SLICE_X9Y138_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y129_SLICE_X5Y129_CQ),
.I2(1'b1),
.I3(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO2),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y138_SLICE_X9Y138_CO5),
.O6(CLBLM_R_X7Y138_SLICE_X9Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3c3c3c3c3c)
  ) CLBLM_R_X7Y138_SLICE_X9Y138_BLUT (
.I0(1'b1),
.I1(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO1),
.I2(CLBLM_R_X5Y129_SLICE_X6Y129_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y138_SLICE_X9Y138_BO5),
.O6(CLBLM_R_X7Y138_SLICE_X9Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff00ff00ff00ff0)
  ) CLBLM_R_X7Y138_SLICE_X9Y138_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X5Y129_SLICE_X7Y129_BQ),
.I3(BRAM_L_X6Y135_RAMB18_X0Y55_DOADO0),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y138_SLICE_X9Y138_AO5),
.O6(CLBLM_R_X7Y138_SLICE_X9Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X7Y139_SLICE_X8Y139_DLUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO1),
.I1(BRAM_L_X6Y140_RAMB18_X0Y56_DO16),
.I2(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO0),
.I3(CLBLM_R_X7Y125_SLICE_X9Y125_AQ),
.I4(BRAM_L_X6Y140_RAMB18_X0Y56_DO17),
.I5(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO1),
.O5(CLBLM_R_X7Y139_SLICE_X8Y139_DO5),
.O6(CLBLM_R_X7Y139_SLICE_X8Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X7Y139_SLICE_X8Y139_CLUT (
.I0(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO2),
.I1(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.I2(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO2),
.I3(BRAM_L_X6Y140_RAMB18_X0Y56_DO18),
.I4(BRAM_L_X6Y140_RAMB18_X0Y56_DO17),
.I5(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO1),
.O5(CLBLM_R_X7Y139_SLICE_X8Y139_CO5),
.O6(CLBLM_R_X7Y139_SLICE_X8Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X7Y139_SLICE_X8Y139_BLUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y56_DO19),
.I1(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.I2(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO3),
.I3(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO4),
.I4(BRAM_L_X6Y140_RAMB18_X0Y56_DO20),
.I5(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO4),
.O5(CLBLM_R_X7Y139_SLICE_X8Y139_BO5),
.O6(CLBLM_R_X7Y139_SLICE_X8Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3a35353acac5c5ca)
  ) CLBLM_R_X7Y139_SLICE_X8Y139_ALUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO7),
.I1(CLBLM_R_X7Y125_SLICE_X9Y125_AQ),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I3(CLBLM_R_X7Y139_SLICE_X8Y139_DO6),
.I4(BRAM_L_X6Y140_RAMB18_X0Y56_DO23),
.I5(CLBLM_R_X3Y142_SLICE_X2Y142_BQ),
.O5(CLBLM_R_X7Y139_SLICE_X8Y139_AO5),
.O6(CLBLM_R_X7Y139_SLICE_X8Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33aa33aaccaaccaa)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_DLUT (
.I0(CLBLM_R_X7Y139_SLICE_X9Y139_AO6),
.I1(CLBLM_R_X5Y132_SLICE_X7Y132_B5Q),
.I2(1'b1),
.I3(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.O5(CLBLM_R_X7Y139_SLICE_X9Y139_DO5),
.O6(CLBLM_R_X7Y139_SLICE_X9Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_CLUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO4),
.I1(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO4),
.I2(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO3),
.I3(CLBLM_R_X5Y133_SLICE_X6Y133_BQ),
.I4(BRAM_L_X6Y140_RAMB18_X0Y56_DO19),
.I5(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO4),
.O5(CLBLM_R_X7Y139_SLICE_X9Y139_CO5),
.O6(CLBLM_R_X7Y139_SLICE_X9Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_BLUT (
.I0(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO4),
.I1(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO5),
.I2(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO5),
.I3(CLBLL_L_X4Y133_SLICE_X4Y133_A5Q),
.I4(BRAM_L_X6Y140_RAMB18_X0Y56_DO20),
.I5(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO5),
.O5(CLBLM_R_X7Y139_SLICE_X9Y139_BO5),
.O6(CLBLM_R_X7Y139_SLICE_X9Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_ALUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO6),
.I1(BRAM_L_X6Y140_RAMB18_X0Y56_DO21),
.I2(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO6),
.I3(BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO6),
.I4(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO5),
.I5(CLBLM_R_X5Y132_SLICE_X7Y132_B5Q),
.O5(CLBLM_R_X7Y139_SLICE_X9Y139_AO5),
.O6(CLBLM_R_X7Y139_SLICE_X9Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4ee44ee44ee44ee4)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_DLUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I1(CLBLM_R_X7Y139_SLICE_X8Y139_CO6),
.I2(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.I3(CLBLM_R_X3Y145_SLICE_X3Y145_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y140_SLICE_X8Y140_DO5),
.O6(CLBLM_R_X7Y140_SLICE_X8Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h50fa50fafa50fa50)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_CLUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y139_SLICE_X9Y139_BO6),
.I3(CLBLL_L_X4Y133_SLICE_X4Y133_A5Q),
.I4(1'b1),
.I5(CLBLM_R_X3Y151_SLICE_X3Y151_AQ),
.O5(CLBLM_R_X7Y140_SLICE_X8Y140_CO5),
.O6(CLBLM_R_X7Y140_SLICE_X8Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3a35353acac5c5ca)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_BLUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y56_DO23),
.I1(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I3(BRAM_L_X6Y140_RAMB18_X0Y57_DOADO7),
.I4(CLBLM_R_X7Y139_SLICE_X8Y139_BO6),
.I5(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.O5(CLBLM_R_X7Y140_SLICE_X8Y140_BO5),
.O6(CLBLM_R_X7Y140_SLICE_X8Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff9696ff009696)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_ALUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y56_DO23),
.I1(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO7),
.I2(CLBLM_R_X7Y139_SLICE_X9Y139_CO6),
.I3(CLBLM_R_X3Y149_SLICE_X2Y149_DQ),
.I4(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I5(CLBLM_R_X5Y133_SLICE_X6Y133_BQ),
.O5(CLBLM_R_X7Y140_SLICE_X8Y140_AO5),
.O6(CLBLM_R_X7Y140_SLICE_X8Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y140_SLICE_X9Y140_DO5),
.O6(CLBLM_R_X7Y140_SLICE_X9Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y140_SLICE_X9Y140_CO5),
.O6(CLBLM_R_X7Y140_SLICE_X9Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y140_SLICE_X9Y140_BO5),
.O6(CLBLM_R_X7Y140_SLICE_X9Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y140_SLICE_X9Y140_AO5),
.O6(CLBLM_R_X7Y140_SLICE_X9Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y130_SLICE_X14Y130_AO6),
.Q(CLBLM_R_X11Y130_SLICE_X14Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y130_SLICE_X14Y130_DO5),
.O6(CLBLM_R_X11Y130_SLICE_X14Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y130_SLICE_X14Y130_CO5),
.O6(CLBLM_R_X11Y130_SLICE_X14Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y130_SLICE_X14Y130_BO5),
.O6(CLBLM_R_X11Y130_SLICE_X14Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff00ff00ff00ff0)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(BRAM_R_X17Y135_RAMB18_X1Y54_DO17),
.I3(CLBLL_L_X4Y131_SLICE_X4Y131_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y130_SLICE_X14Y130_AO5),
.O6(CLBLM_R_X11Y130_SLICE_X14Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y130_SLICE_X15Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y130_SLICE_X15Y130_DO5),
.O6(CLBLM_R_X11Y130_SLICE_X15Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y130_SLICE_X15Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y130_SLICE_X15Y130_CO5),
.O6(CLBLM_R_X11Y130_SLICE_X15Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y130_SLICE_X15Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y130_SLICE_X15Y130_BO5),
.O6(CLBLM_R_X11Y130_SLICE_X15Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y130_SLICE_X15Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y130_SLICE_X15Y130_AO5),
.O6(CLBLM_R_X11Y130_SLICE_X15Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y131_SLICE_X14Y131_AO6),
.Q(CLBLM_R_X11Y131_SLICE_X14Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y131_SLICE_X14Y131_BO6),
.Q(CLBLM_R_X11Y131_SLICE_X14Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y131_SLICE_X14Y131_DO5),
.O6(CLBLM_R_X11Y131_SLICE_X14Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y131_SLICE_X14Y131_CO5),
.O6(CLBLM_R_X11Y131_SLICE_X14Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0ff0f0f0f0)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(BRAM_R_X17Y135_RAMB18_X1Y54_DO23),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X3Y132_SLICE_X2Y132_DQ),
.O5(CLBLM_R_X11Y131_SLICE_X14Y131_BO5),
.O6(CLBLM_R_X11Y131_SLICE_X14Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5a5a5a5a5a)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_ALUT (
.I0(CLBLM_R_X3Y131_SLICE_X3Y131_DQ),
.I1(1'b1),
.I2(BRAM_R_X17Y135_RAMB18_X1Y54_DO20),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y131_SLICE_X14Y131_AO5),
.O6(CLBLM_R_X11Y131_SLICE_X14Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y131_SLICE_X15Y131_DO5),
.O6(CLBLM_R_X11Y131_SLICE_X15Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y131_SLICE_X15Y131_CO5),
.O6(CLBLM_R_X11Y131_SLICE_X15Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y131_SLICE_X15Y131_BO5),
.O6(CLBLM_R_X11Y131_SLICE_X15Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y131_SLICE_X15Y131_AO5),
.O6(CLBLM_R_X11Y131_SLICE_X15Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y133_SLICE_X14Y133_AO6),
.Q(CLBLM_R_X11Y133_SLICE_X14Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y133_SLICE_X14Y133_BO6),
.Q(CLBLM_R_X11Y133_SLICE_X14Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y133_SLICE_X14Y133_DO5),
.O6(CLBLM_R_X11Y133_SLICE_X14Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y133_SLICE_X14Y133_CO5),
.O6(CLBLM_R_X11Y133_SLICE_X14Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ffff00ff00)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO5),
.I4(1'b1),
.I5(CLBLM_R_X7Y132_SLICE_X8Y132_CQ),
.O5(CLBLM_R_X11Y133_SLICE_X14Y133_BO5),
.O6(CLBLM_R_X11Y133_SLICE_X14Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa55aa55aa55aa)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_ALUT (
.I0(BRAM_R_X17Y135_RAMB18_X1Y55_DOADO3),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X7Y132_SLICE_X8Y132_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y133_SLICE_X14Y133_AO5),
.O6(CLBLM_R_X11Y133_SLICE_X14Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y133_SLICE_X15Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y133_SLICE_X15Y133_DO5),
.O6(CLBLM_R_X11Y133_SLICE_X15Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y133_SLICE_X15Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y133_SLICE_X15Y133_CO5),
.O6(CLBLM_R_X11Y133_SLICE_X15Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y133_SLICE_X15Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y133_SLICE_X15Y133_BO5),
.O6(CLBLM_R_X11Y133_SLICE_X15Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y133_SLICE_X15Y133_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y133_SLICE_X15Y133_AO5),
.O6(CLBLM_R_X11Y133_SLICE_X15Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y135_SLICE_X14Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y135_SLICE_X14Y135_DO5),
.O6(CLBLM_R_X11Y135_SLICE_X14Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7744bb887744bb88)
  ) CLBLM_R_X11Y135_SLICE_X14Y135_CLUT (
.I0(CLBLM_R_X25Y153_SLICE_X36Y153_AQ),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y135_SLICE_X12Y135_DO6),
.I4(CLBLM_L_X10Y135_SLICE_X12Y135_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y135_SLICE_X14Y135_CO5),
.O6(CLBLM_R_X11Y135_SLICE_X14Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333cccca55aa55a)
  ) CLBLM_R_X11Y135_SLICE_X14Y135_BLUT (
.I0(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO7),
.I1(CLBLM_L_X8Y135_SLICE_X10Y135_A5Q),
.I2(CLBLM_L_X10Y135_SLICE_X13Y135_DO6),
.I3(BRAM_L_X6Y135_RAMB18_X0Y54_DO7),
.I4(CLBLM_L_X16Y151_SLICE_X22Y151_DQ),
.I5(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.O5(CLBLM_R_X11Y135_SLICE_X14Y135_BO5),
.O6(CLBLM_R_X11Y135_SLICE_X14Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X11Y135_SLICE_X14Y135_ALUT (
.I0(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO7),
.I1(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO0),
.I2(CLBLM_R_X3Y131_SLICE_X3Y131_AQ),
.I3(BRAM_R_X17Y135_RAMB18_X1Y54_DO7),
.I4(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO0),
.I5(BRAM_L_X6Y135_RAMB18_X0Y54_DO0),
.O5(CLBLM_R_X11Y135_SLICE_X14Y135_AO5),
.O6(CLBLM_R_X11Y135_SLICE_X14Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y135_SLICE_X15Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y135_SLICE_X15Y135_DO5),
.O6(CLBLM_R_X11Y135_SLICE_X15Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y135_SLICE_X15Y135_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y135_SLICE_X15Y135_CO5),
.O6(CLBLM_R_X11Y135_SLICE_X15Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y135_SLICE_X15Y135_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y135_SLICE_X15Y135_BO5),
.O6(CLBLM_R_X11Y135_SLICE_X15Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y135_SLICE_X15Y135_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y135_SLICE_X15Y135_AO5),
.O6(CLBLM_R_X11Y135_SLICE_X15Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h77bb77bb44884488)
  ) CLBLM_R_X11Y136_SLICE_X14Y136_DLUT (
.I0(CLBLM_L_X8Y137_SLICE_X10Y137_A5Q),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I2(1'b1),
.I3(CLBLM_R_X25Y153_SLICE_X36Y153_BQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y136_SLICE_X12Y136_AO6),
.O5(CLBLM_R_X11Y136_SLICE_X14Y136_DO5),
.O6(CLBLM_R_X11Y136_SLICE_X14Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X11Y136_SLICE_X14Y136_CLUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO7),
.I1(BRAM_L_X6Y135_RAMB18_X0Y54_DO7),
.I2(BRAM_R_X17Y135_RAMB18_X1Y54_DO7),
.I3(BRAM_L_X6Y135_RAMB18_X0Y54_DO6),
.I4(CLBLM_L_X8Y137_SLICE_X10Y137_B5Q),
.I5(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO6),
.O5(CLBLM_R_X11Y136_SLICE_X14Y136_CO5),
.O6(CLBLM_R_X11Y136_SLICE_X14Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X11Y136_SLICE_X14Y136_BLUT (
.I0(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO6),
.I1(BRAM_R_X17Y135_RAMB18_X1Y54_DO5),
.I2(CLBLM_R_X3Y132_SLICE_X2Y132_AQ),
.I3(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO6),
.I4(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO5),
.I5(BRAM_L_X6Y135_RAMB18_X0Y54_DO6),
.O5(CLBLM_R_X11Y136_SLICE_X14Y136_BO5),
.O6(CLBLM_R_X11Y136_SLICE_X14Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X11Y136_SLICE_X14Y136_ALUT (
.I0(BRAM_R_X17Y135_RAMB18_X1Y54_DO6),
.I1(CLBLM_R_X3Y132_SLICE_X2Y132_BQ),
.I2(BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO7),
.I3(BRAM_L_X6Y135_RAMB18_X0Y54_DO7),
.I4(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO7),
.I5(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO6),
.O5(CLBLM_R_X11Y136_SLICE_X14Y136_AO5),
.O6(CLBLM_R_X11Y136_SLICE_X14Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y136_SLICE_X15Y136_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y136_SLICE_X15Y136_DO5),
.O6(CLBLM_R_X11Y136_SLICE_X15Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y136_SLICE_X15Y136_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y136_SLICE_X15Y136_CO5),
.O6(CLBLM_R_X11Y136_SLICE_X15Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y136_SLICE_X15Y136_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y136_SLICE_X15Y136_BO5),
.O6(CLBLM_R_X11Y136_SLICE_X15Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y136_SLICE_X15Y136_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y136_SLICE_X15Y136_AO5),
.O6(CLBLM_R_X11Y136_SLICE_X15Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y135_SLICE_X18Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y135_SLICE_X18Y135_DO5),
.O6(CLBLM_R_X13Y135_SLICE_X18Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y135_SLICE_X18Y135_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y135_SLICE_X18Y135_CO5),
.O6(CLBLM_R_X13Y135_SLICE_X18Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y135_SLICE_X18Y135_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y135_SLICE_X18Y135_BO5),
.O6(CLBLM_R_X13Y135_SLICE_X18Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cc33ccffff0000)
  ) CLBLM_R_X13Y135_SLICE_X18Y135_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X25Y157_SLICE_X37Y157_AQ),
.I2(1'b1),
.I3(CLBLM_R_X3Y133_SLICE_X3Y133_AQ),
.I4(CLBLM_L_X10Y135_SLICE_X12Y135_BO6),
.I5(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.O5(CLBLM_R_X13Y135_SLICE_X18Y135_AO5),
.O6(CLBLM_R_X13Y135_SLICE_X18Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y135_SLICE_X19Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y135_SLICE_X19Y135_DO5),
.O6(CLBLM_R_X13Y135_SLICE_X19Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y135_SLICE_X19Y135_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y135_SLICE_X19Y135_CO5),
.O6(CLBLM_R_X13Y135_SLICE_X19Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y135_SLICE_X19Y135_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y135_SLICE_X19Y135_BO5),
.O6(CLBLM_R_X13Y135_SLICE_X19Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y135_SLICE_X19Y135_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y135_SLICE_X19Y135_AO5),
.O6(CLBLM_R_X13Y135_SLICE_X19Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y136_SLICE_X18Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y136_SLICE_X18Y136_AO6),
.Q(CLBLM_R_X13Y136_SLICE_X18Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y136_SLICE_X18Y136_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y136_SLICE_X18Y136_DO5),
.O6(CLBLM_R_X13Y136_SLICE_X18Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y136_SLICE_X18Y136_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y136_SLICE_X18Y136_CO5),
.O6(CLBLM_R_X13Y136_SLICE_X18Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7b7b7b7b48484848)
  ) CLBLM_R_X13Y136_SLICE_X18Y136_BLUT (
.I0(CLBLM_L_X8Y137_SLICE_X10Y137_B5Q),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I2(CLBLM_L_X16Y154_SLICE_X22Y154_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X11Y136_SLICE_X14Y136_CO6),
.O5(CLBLM_R_X13Y136_SLICE_X18Y136_BO5),
.O6(CLBLM_R_X13Y136_SLICE_X18Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff00ff00ff00ff0)
  ) CLBLM_R_X13Y136_SLICE_X18Y136_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(BRAM_R_X17Y135_RAMB18_X1Y54_DO5),
.I3(CLBLM_R_X3Y133_SLICE_X3Y133_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y136_SLICE_X18Y136_AO5),
.O6(CLBLM_R_X13Y136_SLICE_X18Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y136_SLICE_X19Y136_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y136_SLICE_X19Y136_DO5),
.O6(CLBLM_R_X13Y136_SLICE_X19Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y136_SLICE_X19Y136_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y136_SLICE_X19Y136_CO5),
.O6(CLBLM_R_X13Y136_SLICE_X19Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y136_SLICE_X19Y136_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y136_SLICE_X19Y136_BO5),
.O6(CLBLM_R_X13Y136_SLICE_X19Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y136_SLICE_X19Y136_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y136_SLICE_X19Y136_AO5),
.O6(CLBLM_R_X13Y136_SLICE_X19Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y135_SLICE_X20Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y135_SLICE_X20Y135_DO5),
.O6(CLBLM_R_X15Y135_SLICE_X20Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y135_SLICE_X20Y135_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y135_SLICE_X20Y135_CO5),
.O6(CLBLM_R_X15Y135_SLICE_X20Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y135_SLICE_X20Y135_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y135_SLICE_X20Y135_BO5),
.O6(CLBLM_R_X15Y135_SLICE_X20Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y135_SLICE_X20Y135_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y135_SLICE_X20Y135_AO5),
.O6(CLBLM_R_X15Y135_SLICE_X20Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y135_SLICE_X21Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X15Y135_SLICE_X21Y135_AO6),
.Q(CLBLM_R_X15Y135_SLICE_X21Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y135_SLICE_X21Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y135_SLICE_X21Y135_DO5),
.O6(CLBLM_R_X15Y135_SLICE_X21Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y135_SLICE_X21Y135_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y135_SLICE_X21Y135_CO5),
.O6(CLBLM_R_X15Y135_SLICE_X21Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555aaaac33cc33c)
  ) CLBLM_R_X15Y135_SLICE_X21Y135_BLUT (
.I0(CLBLL_L_X4Y132_SLICE_X4Y132_AQ),
.I1(BRAM_R_X17Y135_RAMB18_X1Y54_DO7),
.I2(CLBLM_L_X10Y135_SLICE_X13Y135_BO6),
.I3(BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO7),
.I4(CLBLM_R_X25Y157_SLICE_X36Y157_AQ),
.I5(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.O5(CLBLM_R_X15Y135_SLICE_X21Y135_BO5),
.O6(CLBLM_R_X15Y135_SLICE_X21Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6666666666666666)
  ) CLBLM_R_X15Y135_SLICE_X21Y135_ALUT (
.I0(CLBLL_L_X4Y132_SLICE_X4Y132_AQ),
.I1(BRAM_R_X17Y135_RAMB18_X1Y54_DO1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y135_SLICE_X21Y135_AO5),
.O6(CLBLM_R_X15Y135_SLICE_X21Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X25Y149_SLICE_X36Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(RIOB33_X105Y179_IOB_X1Y179_I),
.Q(CLBLM_R_X25Y149_SLICE_X36Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X25Y149_SLICE_X36Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(RIOB33_X105Y179_IOB_X1Y180_I),
.Q(CLBLM_R_X25Y149_SLICE_X36Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y149_SLICE_X36Y149_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y149_SLICE_X36Y149_DO5),
.O6(CLBLM_R_X25Y149_SLICE_X36Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y149_SLICE_X36Y149_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y149_SLICE_X36Y149_CO5),
.O6(CLBLM_R_X25Y149_SLICE_X36Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y149_SLICE_X36Y149_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y149_SLICE_X36Y149_BO5),
.O6(CLBLM_R_X25Y149_SLICE_X36Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y149_SLICE_X36Y149_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y149_SLICE_X36Y149_AO5),
.O6(CLBLM_R_X25Y149_SLICE_X36Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X25Y149_SLICE_X37Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(RIOB33_X105Y181_IOB_X1Y182_I),
.Q(CLBLM_R_X25Y149_SLICE_X37Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y149_SLICE_X37Y149_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y149_SLICE_X37Y149_DO5),
.O6(CLBLM_R_X25Y149_SLICE_X37Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y149_SLICE_X37Y149_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y149_SLICE_X37Y149_CO5),
.O6(CLBLM_R_X25Y149_SLICE_X37Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y149_SLICE_X37Y149_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y149_SLICE_X37Y149_BO5),
.O6(CLBLM_R_X25Y149_SLICE_X37Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y149_SLICE_X37Y149_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y149_SLICE_X37Y149_AO5),
.O6(CLBLM_R_X25Y149_SLICE_X37Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X25Y151_SLICE_X36Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(RIOB33_X105Y183_IOB_X1Y184_I),
.Q(CLBLM_R_X25Y151_SLICE_X36Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X25Y151_SLICE_X36Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(RIOB33_X105Y187_IOB_X1Y188_I),
.Q(CLBLM_R_X25Y151_SLICE_X36Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X25Y151_SLICE_X36Y151_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(RIOB33_X105Y189_IOB_X1Y189_I),
.Q(CLBLM_R_X25Y151_SLICE_X36Y151_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y151_SLICE_X36Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y151_SLICE_X36Y151_DO5),
.O6(CLBLM_R_X25Y151_SLICE_X36Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y151_SLICE_X36Y151_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y151_SLICE_X36Y151_CO5),
.O6(CLBLM_R_X25Y151_SLICE_X36Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y151_SLICE_X36Y151_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y151_SLICE_X36Y151_BO5),
.O6(CLBLM_R_X25Y151_SLICE_X36Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y151_SLICE_X36Y151_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y151_SLICE_X36Y151_AO5),
.O6(CLBLM_R_X25Y151_SLICE_X36Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y151_SLICE_X37Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y151_SLICE_X37Y151_DO5),
.O6(CLBLM_R_X25Y151_SLICE_X37Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y151_SLICE_X37Y151_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y151_SLICE_X37Y151_CO5),
.O6(CLBLM_R_X25Y151_SLICE_X37Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y151_SLICE_X37Y151_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y151_SLICE_X37Y151_BO5),
.O6(CLBLM_R_X25Y151_SLICE_X37Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y151_SLICE_X37Y151_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y151_SLICE_X37Y151_AO5),
.O6(CLBLM_R_X25Y151_SLICE_X37Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X25Y153_SLICE_X36Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(RIOB33_X105Y195_IOB_X1Y195_I),
.Q(CLBLM_R_X25Y153_SLICE_X36Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X25Y153_SLICE_X36Y153_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(RIOB33_X105Y195_IOB_X1Y196_I),
.Q(CLBLM_R_X25Y153_SLICE_X36Y153_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y153_SLICE_X36Y153_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y153_SLICE_X36Y153_DO5),
.O6(CLBLM_R_X25Y153_SLICE_X36Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y153_SLICE_X36Y153_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y153_SLICE_X36Y153_CO5),
.O6(CLBLM_R_X25Y153_SLICE_X36Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y153_SLICE_X36Y153_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y153_SLICE_X36Y153_BO5),
.O6(CLBLM_R_X25Y153_SLICE_X36Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y153_SLICE_X36Y153_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y153_SLICE_X36Y153_AO5),
.O6(CLBLM_R_X25Y153_SLICE_X36Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y153_SLICE_X37Y153_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y153_SLICE_X37Y153_DO5),
.O6(CLBLM_R_X25Y153_SLICE_X37Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y153_SLICE_X37Y153_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y153_SLICE_X37Y153_CO5),
.O6(CLBLM_R_X25Y153_SLICE_X37Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y153_SLICE_X37Y153_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y153_SLICE_X37Y153_BO5),
.O6(CLBLM_R_X25Y153_SLICE_X37Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y153_SLICE_X37Y153_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y153_SLICE_X37Y153_AO5),
.O6(CLBLM_R_X25Y153_SLICE_X37Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X25Y154_SLICE_X36Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(RIOB33_SING_X105Y200_IOB_X1Y200_I),
.Q(CLBLM_R_X25Y154_SLICE_X36Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X25Y154_SLICE_X36Y154_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(RIOB33_X105Y197_IOB_X1Y198_I),
.Q(CLBLM_R_X25Y154_SLICE_X36Y154_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X25Y154_SLICE_X36Y154_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(RIOB33_SING_X105Y199_IOB_X1Y199_I),
.Q(CLBLM_R_X25Y154_SLICE_X36Y154_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y154_SLICE_X36Y154_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y154_SLICE_X36Y154_DO5),
.O6(CLBLM_R_X25Y154_SLICE_X36Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y154_SLICE_X36Y154_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y154_SLICE_X36Y154_CO5),
.O6(CLBLM_R_X25Y154_SLICE_X36Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y154_SLICE_X36Y154_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y154_SLICE_X36Y154_BO5),
.O6(CLBLM_R_X25Y154_SLICE_X36Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y154_SLICE_X36Y154_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y154_SLICE_X36Y154_AO5),
.O6(CLBLM_R_X25Y154_SLICE_X36Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y154_SLICE_X37Y154_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y154_SLICE_X37Y154_DO5),
.O6(CLBLM_R_X25Y154_SLICE_X37Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y154_SLICE_X37Y154_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y154_SLICE_X37Y154_CO5),
.O6(CLBLM_R_X25Y154_SLICE_X37Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y154_SLICE_X37Y154_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y154_SLICE_X37Y154_BO5),
.O6(CLBLM_R_X25Y154_SLICE_X37Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y154_SLICE_X37Y154_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y154_SLICE_X37Y154_AO5),
.O6(CLBLM_R_X25Y154_SLICE_X37Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X25Y157_SLICE_X36Y157_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(RIOB33_X105Y201_IOB_X1Y201_I),
.Q(CLBLM_R_X25Y157_SLICE_X36Y157_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X25Y157_SLICE_X36Y157_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(RIOB33_X105Y203_IOB_X1Y204_I),
.Q(CLBLM_R_X25Y157_SLICE_X36Y157_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y157_SLICE_X36Y157_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y157_SLICE_X36Y157_DO5),
.O6(CLBLM_R_X25Y157_SLICE_X36Y157_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y157_SLICE_X36Y157_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y157_SLICE_X36Y157_CO5),
.O6(CLBLM_R_X25Y157_SLICE_X36Y157_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y157_SLICE_X36Y157_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y157_SLICE_X36Y157_BO5),
.O6(CLBLM_R_X25Y157_SLICE_X36Y157_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y157_SLICE_X36Y157_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y157_SLICE_X36Y157_AO5),
.O6(CLBLM_R_X25Y157_SLICE_X36Y157_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X25Y157_SLICE_X37Y157_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y147_IOB_X0Y148_I),
.D(RIOB33_X105Y205_IOB_X1Y205_I),
.Q(CLBLM_R_X25Y157_SLICE_X37Y157_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y157_SLICE_X37Y157_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y157_SLICE_X37Y157_DO5),
.O6(CLBLM_R_X25Y157_SLICE_X37Y157_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y157_SLICE_X37Y157_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y157_SLICE_X37Y157_CO5),
.O6(CLBLM_R_X25Y157_SLICE_X37Y157_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y157_SLICE_X37Y157_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y157_SLICE_X37Y157_BO5),
.O6(CLBLM_R_X25Y157_SLICE_X37Y157_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y157_SLICE_X37Y157_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y157_SLICE_X37Y157_AO5),
.O6(CLBLM_R_X25Y157_SLICE_X37Y157_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(LIOB33_X0Y127_IOB_X0Y128_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X139Y78_BUFHCE_X0Y20_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X139Y78_BUFHCE_X0Y20_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_TOP_R_X139Y182_BUFHCE_X1Y44_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_TOP_R_X139Y182_BUFHCE_X1Y44_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y1_IOB_X0Y1_IBUF (
.I(LIOB33_X0Y1_IOB_X0Y1_IPAD),
.O(LIOB33_X0Y1_IOB_X0Y1_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y1_IOB_X0Y2_IBUF (
.I(LIOB33_X0Y1_IOB_X0Y2_IPAD),
.O(LIOB33_X0Y1_IOB_X0Y2_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y3_IOB_X0Y3_IBUF (
.I(LIOB33_X0Y3_IOB_X0Y3_IPAD),
.O(LIOB33_X0Y3_IOB_X0Y3_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y3_IOB_X0Y4_IBUF (
.I(LIOB33_X0Y3_IOB_X0Y4_IPAD),
.O(LIOB33_X0Y3_IOB_X0Y4_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y5_IOB_X0Y5_IBUF (
.I(LIOB33_X0Y5_IOB_X0Y5_IPAD),
.O(LIOB33_X0Y5_IOB_X0Y5_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y5_IOB_X0Y6_IBUF (
.I(LIOB33_X0Y5_IOB_X0Y6_IPAD),
.O(LIOB33_X0Y5_IOB_X0Y6_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y7_IOB_X0Y7_IBUF (
.I(LIOB33_X0Y7_IOB_X0Y7_IPAD),
.O(LIOB33_X0Y7_IOB_X0Y7_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y7_IOB_X0Y8_IBUF (
.I(LIOB33_X0Y7_IOB_X0Y8_IPAD),
.O(LIOB33_X0Y7_IOB_X0Y8_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y9_IOB_X0Y9_IBUF (
.I(LIOB33_X0Y9_IOB_X0Y9_IPAD),
.O(LIOB33_X0Y9_IOB_X0Y9_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y9_IOB_X0Y10_IBUF (
.I(LIOB33_X0Y9_IOB_X0Y10_IPAD),
.O(LIOB33_X0Y9_IOB_X0Y10_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y11_IOB_X0Y11_IBUF (
.I(LIOB33_X0Y11_IOB_X0Y11_IPAD),
.O(LIOB33_X0Y11_IOB_X0Y11_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y11_IOB_X0Y12_IBUF (
.I(LIOB33_X0Y11_IOB_X0Y12_IPAD),
.O(LIOB33_X0Y11_IOB_X0Y12_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y13_IOB_X0Y13_IBUF (
.I(LIOB33_X0Y13_IOB_X0Y13_IPAD),
.O(LIOB33_X0Y13_IOB_X0Y13_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y13_IOB_X0Y14_IBUF (
.I(LIOB33_X0Y13_IOB_X0Y14_IPAD),
.O(LIOB33_X0Y13_IOB_X0Y14_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y15_IOB_X0Y15_IBUF (
.I(LIOB33_X0Y15_IOB_X0Y15_IPAD),
.O(LIOB33_X0Y15_IOB_X0Y15_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y15_IOB_X0Y16_IBUF (
.I(LIOB33_X0Y15_IOB_X0Y16_IPAD),
.O(LIOB33_X0Y15_IOB_X0Y16_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y17_IOB_X0Y17_IBUF (
.I(LIOB33_X0Y17_IOB_X0Y17_IPAD),
.O(LIOB33_X0Y17_IOB_X0Y17_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y17_IOB_X0Y18_IBUF (
.I(LIOB33_X0Y17_IOB_X0Y18_IPAD),
.O(LIOB33_X0Y17_IOB_X0Y18_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y19_IOB_X0Y19_IBUF (
.I(LIOB33_X0Y19_IOB_X0Y19_IPAD),
.O(LIOB33_X0Y19_IOB_X0Y19_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y19_IOB_X0Y20_IBUF (
.I(LIOB33_X0Y19_IOB_X0Y20_IPAD),
.O(LIOB33_X0Y19_IOB_X0Y20_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y21_IOB_X0Y21_IBUF (
.I(LIOB33_X0Y21_IOB_X0Y21_IPAD),
.O(LIOB33_X0Y21_IOB_X0Y21_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y21_IOB_X0Y22_IBUF (
.I(LIOB33_X0Y21_IOB_X0Y22_IPAD),
.O(LIOB33_X0Y21_IOB_X0Y22_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y23_IOB_X0Y23_IBUF (
.I(LIOB33_X0Y23_IOB_X0Y23_IPAD),
.O(LIOB33_X0Y23_IOB_X0Y23_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y23_IOB_X0Y24_IBUF (
.I(LIOB33_X0Y23_IOB_X0Y24_IPAD),
.O(LIOB33_X0Y23_IOB_X0Y24_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y25_IOB_X0Y25_IBUF (
.I(LIOB33_X0Y25_IOB_X0Y25_IPAD),
.O(LIOB33_X0Y25_IOB_X0Y25_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y25_IOB_X0Y26_IBUF (
.I(LIOB33_X0Y25_IOB_X0Y26_IPAD),
.O(LIOB33_X0Y25_IOB_X0Y26_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y27_IOB_X0Y27_IBUF (
.I(LIOB33_X0Y27_IOB_X0Y27_IPAD),
.O(LIOB33_X0Y27_IOB_X0Y27_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y27_IOB_X0Y28_IBUF (
.I(LIOB33_X0Y27_IOB_X0Y28_IPAD),
.O(LIOB33_X0Y27_IOB_X0Y28_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y29_IOB_X0Y29_IBUF (
.I(LIOB33_X0Y29_IOB_X0Y29_IPAD),
.O(LIOB33_X0Y29_IOB_X0Y29_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y29_IOB_X0Y30_IBUF (
.I(LIOB33_X0Y29_IOB_X0Y30_IPAD),
.O(LIOB33_X0Y29_IOB_X0Y30_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y31_IOB_X0Y31_IBUF (
.I(LIOB33_X0Y31_IOB_X0Y31_IPAD),
.O(LIOB33_X0Y31_IOB_X0Y31_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y51_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y51_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y51_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y52_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y52_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y52_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y53_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y53_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y53_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y54_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y54_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y54_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y55_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y55_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y55_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y56_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y56_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y56_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y57_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y57_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y57_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y58_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y58_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y58_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y59_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y59_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y59_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y60_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y60_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y60_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y61_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y61_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y61_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y62_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y62_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y62_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y63_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y63_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y63_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y64_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y64_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y64_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y65_IOB_X0Y65_IBUF (
.I(LIOB33_X0Y65_IOB_X0Y65_IPAD),
.O(LIOB33_X0Y65_IOB_X0Y65_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y65_IOB_X0Y66_IBUF (
.I(LIOB33_X0Y65_IOB_X0Y66_IPAD),
.O(LIOB33_X0Y65_IOB_X0Y66_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y67_IOB_X0Y67_IBUF (
.I(LIOB33_X0Y67_IOB_X0Y67_IPAD),
.O(LIOB33_X0Y67_IOB_X0Y67_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y67_IOB_X0Y68_IBUF (
.I(LIOB33_X0Y67_IOB_X0Y68_IPAD),
.O(LIOB33_X0Y67_IOB_X0Y68_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y69_IOB_X0Y69_IBUF (
.I(LIOB33_X0Y69_IOB_X0Y69_IPAD),
.O(LIOB33_X0Y69_IOB_X0Y69_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y69_IOB_X0Y70_IBUF (
.I(LIOB33_X0Y69_IOB_X0Y70_IPAD),
.O(LIOB33_X0Y69_IOB_X0Y70_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y71_IOB_X0Y71_IBUF (
.I(LIOB33_X0Y71_IOB_X0Y71_IPAD),
.O(LIOB33_X0Y71_IOB_X0Y71_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y71_IOB_X0Y72_IBUF (
.I(LIOB33_X0Y71_IOB_X0Y72_IPAD),
.O(LIOB33_X0Y71_IOB_X0Y72_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y73_IOB_X0Y73_IBUF (
.I(LIOB33_X0Y73_IOB_X0Y73_IPAD),
.O(LIOB33_X0Y73_IOB_X0Y73_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y73_IOB_X0Y74_IBUF (
.I(LIOB33_X0Y73_IOB_X0Y74_IPAD),
.O(LIOB33_X0Y73_IOB_X0Y74_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y75_IOB_X0Y75_IBUF (
.I(LIOB33_X0Y75_IOB_X0Y75_IPAD),
.O(LIOB33_X0Y75_IOB_X0Y75_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y75_IOB_X0Y76_IBUF (
.I(LIOB33_X0Y75_IOB_X0Y76_IPAD),
.O(LIOB33_X0Y75_IOB_X0Y76_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y77_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y77_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y77_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y78_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y78_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y78_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y79_IOB_X0Y79_IBUF (
.I(LIOB33_X0Y79_IOB_X0Y79_IPAD),
.O(LIOB33_X0Y79_IOB_X0Y79_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y79_IOB_X0Y80_IBUF (
.I(LIOB33_X0Y79_IOB_X0Y80_IPAD),
.O(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y81_IOB_X0Y81_IBUF (
.I(LIOB33_X0Y81_IOB_X0Y81_IPAD),
.O(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y81_IOB_X0Y82_IBUF (
.I(LIOB33_X0Y81_IOB_X0Y82_IPAD),
.O(LIOB33_X0Y81_IOB_X0Y82_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y83_IOB_X0Y83_IBUF (
.I(LIOB33_X0Y83_IOB_X0Y83_IPAD),
.O(LIOB33_X0Y83_IOB_X0Y83_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y83_IOB_X0Y84_IBUF (
.I(LIOB33_X0Y83_IOB_X0Y84_IPAD),
.O(LIOB33_X0Y83_IOB_X0Y84_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y85_IOB_X0Y85_IBUF (
.I(LIOB33_X0Y85_IOB_X0Y85_IPAD),
.O(LIOB33_X0Y85_IOB_X0Y85_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y85_IOB_X0Y86_IBUF (
.I(LIOB33_X0Y85_IOB_X0Y86_IPAD),
.O(LIOB33_X0Y85_IOB_X0Y86_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y87_IOB_X0Y87_IBUF (
.I(LIOB33_X0Y87_IOB_X0Y87_IPAD),
.O(LIOB33_X0Y87_IOB_X0Y87_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y87_IOB_X0Y88_IBUF (
.I(LIOB33_X0Y87_IOB_X0Y88_IPAD),
.O(LIOB33_X0Y87_IOB_X0Y88_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y89_IOB_X0Y89_IBUF (
.I(LIOB33_X0Y89_IOB_X0Y89_IPAD),
.O(LIOB33_X0Y89_IOB_X0Y89_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y89_IOB_X0Y90_IBUF (
.I(LIOB33_X0Y89_IOB_X0Y90_IPAD),
.O(LIOB33_X0Y89_IOB_X0Y90_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y91_IOB_X0Y91_IBUF (
.I(LIOB33_X0Y91_IOB_X0Y91_IPAD),
.O(LIOB33_X0Y91_IOB_X0Y91_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y91_IOB_X0Y92_IBUF (
.I(LIOB33_X0Y91_IOB_X0Y92_IPAD),
.O(LIOB33_X0Y91_IOB_X0Y92_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y93_IOB_X0Y93_IBUF (
.I(LIOB33_X0Y93_IOB_X0Y93_IPAD),
.O(LIOB33_X0Y93_IOB_X0Y93_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y93_IOB_X0Y94_IBUF (
.I(LIOB33_X0Y93_IOB_X0Y94_IPAD),
.O(LIOB33_X0Y93_IOB_X0Y94_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y95_IOB_X0Y95_IBUF (
.I(LIOB33_X0Y95_IOB_X0Y95_IPAD),
.O(LIOB33_X0Y95_IOB_X0Y95_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y95_IOB_X0Y96_IBUF (
.I(LIOB33_X0Y95_IOB_X0Y96_IPAD),
.O(LIOB33_X0Y95_IOB_X0Y96_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y97_IOB_X0Y97_IBUF (
.I(LIOB33_X0Y97_IOB_X0Y97_IPAD),
.O(LIOB33_X0Y97_IOB_X0Y97_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y97_IOB_X0Y98_IBUF (
.I(LIOB33_X0Y97_IOB_X0Y98_IPAD),
.O(LIOB33_X0Y97_IOB_X0Y98_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y101_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y101_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y102_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y102_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y103_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y103_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y104_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y104_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y105_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y105_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y106_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y106_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y107_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y107_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y108_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y108_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y109_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y109_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y110_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y110_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y111_IOB_X0Y111_IBUF (
.I(LIOB33_X0Y111_IOB_X0Y111_IPAD),
.O(LIOB33_X0Y111_IOB_X0Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y111_IOB_X0Y112_IBUF (
.I(LIOB33_X0Y111_IOB_X0Y112_IPAD),
.O(LIOB33_X0Y111_IOB_X0Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y113_IOB_X0Y113_IBUF (
.I(LIOB33_X0Y113_IOB_X0Y113_IPAD),
.O(LIOB33_X0Y113_IOB_X0Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y113_IOB_X0Y114_IBUF (
.I(LIOB33_X0Y113_IOB_X0Y114_IPAD),
.O(LIOB33_X0Y113_IOB_X0Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y115_IOB_X0Y115_IBUF (
.I(LIOB33_X0Y115_IOB_X0Y115_IPAD),
.O(LIOB33_X0Y115_IOB_X0Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y115_IOB_X0Y116_IBUF (
.I(LIOB33_X0Y115_IOB_X0Y116_IPAD),
.O(LIOB33_X0Y115_IOB_X0Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y117_IOB_X0Y117_IBUF (
.I(LIOB33_X0Y117_IOB_X0Y117_IPAD),
.O(LIOB33_X0Y117_IOB_X0Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y117_IOB_X0Y118_IBUF (
.I(LIOB33_X0Y117_IOB_X0Y118_IPAD),
.O(LIOB33_X0Y117_IOB_X0Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y119_IOB_X0Y119_IBUF (
.I(LIOB33_X0Y119_IOB_X0Y119_IPAD),
.O(LIOB33_X0Y119_IOB_X0Y119_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y119_IOB_X0Y120_IBUF (
.I(LIOB33_X0Y119_IOB_X0Y120_IPAD),
.O(LIOB33_X0Y119_IOB_X0Y120_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y121_IOB_X0Y121_IBUF (
.I(LIOB33_X0Y121_IOB_X0Y121_IPAD),
.O(LIOB33_X0Y121_IOB_X0Y121_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y121_IOB_X0Y122_IBUF (
.I(LIOB33_X0Y121_IOB_X0Y122_IPAD),
.O(LIOB33_X0Y121_IOB_X0Y122_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y123_IOB_X0Y123_IBUF (
.I(LIOB33_X0Y123_IOB_X0Y123_IPAD),
.O(LIOB33_X0Y123_IOB_X0Y123_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y123_IOB_X0Y124_IBUF (
.I(LIOB33_X0Y123_IOB_X0Y124_IPAD),
.O(LIOB33_X0Y123_IOB_X0Y124_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y125_IOB_X0Y125_IBUF (
.I(LIOB33_X0Y125_IOB_X0Y125_IPAD),
.O(LIOB33_X0Y125_IOB_X0Y125_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y125_IOB_X0Y126_IBUF (
.I(LIOB33_X0Y125_IOB_X0Y126_IPAD),
.O(LIOB33_X0Y125_IOB_X0Y126_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y127_IOB_X0Y127_IBUF (
.I(LIOB33_X0Y127_IOB_X0Y127_IPAD),
.O(LIOB33_X0Y127_IOB_X0Y127_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y127_IOB_X0Y128_IBUF (
.I(LIOB33_X0Y127_IOB_X0Y128_IPAD),
.O(LIOB33_X0Y127_IOB_X0Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y129_IOB_X0Y129_IBUF (
.I(LIOB33_X0Y129_IOB_X0Y129_IPAD),
.O(LIOB33_X0Y129_IOB_X0Y129_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y129_IOB_X0Y130_IBUF (
.I(LIOB33_X0Y129_IOB_X0Y130_IPAD),
.O(LIOB33_X0Y129_IOB_X0Y130_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y131_IOB_X0Y131_IBUF (
.I(LIOB33_X0Y131_IOB_X0Y131_IPAD),
.O(LIOB33_X0Y131_IOB_X0Y131_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y131_IOB_X0Y132_IBUF (
.I(LIOB33_X0Y131_IOB_X0Y132_IPAD),
.O(LIOB33_X0Y131_IOB_X0Y132_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y133_IOB_X0Y133_IBUF (
.I(LIOB33_X0Y133_IOB_X0Y133_IPAD),
.O(LIOB33_X0Y133_IOB_X0Y133_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y133_IOB_X0Y134_IBUF (
.I(LIOB33_X0Y133_IOB_X0Y134_IPAD),
.O(LIOB33_X0Y133_IOB_X0Y134_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y135_IOB_X0Y135_IBUF (
.I(LIOB33_X0Y135_IOB_X0Y135_IPAD),
.O(LIOB33_X0Y135_IOB_X0Y135_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y135_IOB_X0Y136_IBUF (
.I(LIOB33_X0Y135_IOB_X0Y136_IPAD),
.O(LIOB33_X0Y135_IOB_X0Y136_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y137_IOB_X0Y137_IBUF (
.I(LIOB33_X0Y137_IOB_X0Y137_IPAD),
.O(LIOB33_X0Y137_IOB_X0Y137_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y137_IOB_X0Y138_IBUF (
.I(LIOB33_X0Y137_IOB_X0Y138_IPAD),
.O(LIOB33_X0Y137_IOB_X0Y138_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y139_IOB_X0Y139_IBUF (
.I(LIOB33_X0Y139_IOB_X0Y139_IPAD),
.O(LIOB33_X0Y139_IOB_X0Y139_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y139_IOB_X0Y140_IBUF (
.I(LIOB33_X0Y139_IOB_X0Y140_IPAD),
.O(LIOB33_X0Y139_IOB_X0Y140_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y141_IOB_X0Y141_IBUF (
.I(LIOB33_X0Y141_IOB_X0Y141_IPAD),
.O(LIOB33_X0Y141_IOB_X0Y141_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y141_IOB_X0Y142_IBUF (
.I(LIOB33_X0Y141_IOB_X0Y142_IPAD),
.O(LIOB33_X0Y141_IOB_X0Y142_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y143_IOB_X0Y143_IBUF (
.I(LIOB33_X0Y143_IOB_X0Y143_IPAD),
.O(LIOB33_X0Y143_IOB_X0Y143_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y145_IOB_X0Y145_IBUF (
.I(LIOB33_X0Y145_IOB_X0Y145_IPAD),
.O(LIOB33_X0Y145_IOB_X0Y145_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y145_IOB_X0Y146_IBUF (
.I(LIOB33_X0Y145_IOB_X0Y146_IPAD),
.O(LIOB33_X0Y145_IOB_X0Y146_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y147_IOB_X0Y147_IBUF (
.I(LIOB33_X0Y147_IOB_X0Y147_IPAD),
.O(LIOB33_X0Y147_IOB_X0Y147_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y147_IOB_X0Y148_IBUF (
.I(LIOB33_X0Y147_IOB_X0Y148_IPAD),
.O(LIOB33_X0Y147_IOB_X0Y148_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y151_IOB_X0Y151_IBUF (
.I(LIOB33_X0Y151_IOB_X0Y151_IPAD),
.O(LIOB33_X0Y151_IOB_X0Y151_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y151_IOB_X0Y152_IBUF (
.I(LIOB33_X0Y151_IOB_X0Y152_IPAD),
.O(LIOB33_X0Y151_IOB_X0Y152_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y153_IOB_X0Y153_IBUF (
.I(LIOB33_X0Y153_IOB_X0Y153_IPAD),
.O(LIOB33_X0Y153_IOB_X0Y153_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y153_IOB_X0Y154_IBUF (
.I(LIOB33_X0Y153_IOB_X0Y154_IPAD),
.O(LIOB33_X0Y153_IOB_X0Y154_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y155_IOB_X0Y155_IBUF (
.I(LIOB33_X0Y155_IOB_X0Y155_IPAD),
.O(LIOB33_X0Y155_IOB_X0Y155_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y155_IOB_X0Y156_IBUF (
.I(LIOB33_X0Y155_IOB_X0Y156_IPAD),
.O(LIOB33_X0Y155_IOB_X0Y156_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y157_IOB_X0Y157_IBUF (
.I(LIOB33_X0Y157_IOB_X0Y157_IPAD),
.O(LIOB33_X0Y157_IOB_X0Y157_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y157_IOB_X0Y158_IBUF (
.I(LIOB33_X0Y157_IOB_X0Y158_IPAD),
.O(LIOB33_X0Y157_IOB_X0Y158_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y159_IOB_X0Y159_IBUF (
.I(LIOB33_X0Y159_IOB_X0Y159_IPAD),
.O(LIOB33_X0Y159_IOB_X0Y159_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y159_IOB_X0Y160_IBUF (
.I(LIOB33_X0Y159_IOB_X0Y160_IPAD),
.O(LIOB33_X0Y159_IOB_X0Y160_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y161_IOB_X0Y161_IBUF (
.I(LIOB33_X0Y161_IOB_X0Y161_IPAD),
.O(LIOB33_X0Y161_IOB_X0Y161_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y161_IOB_X0Y162_IBUF (
.I(LIOB33_X0Y161_IOB_X0Y162_IPAD),
.O(LIOB33_X0Y161_IOB_X0Y162_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y163_IOB_X0Y163_IBUF (
.I(LIOB33_X0Y163_IOB_X0Y163_IPAD),
.O(LIOB33_X0Y163_IOB_X0Y163_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y163_IOB_X0Y164_IBUF (
.I(LIOB33_X0Y163_IOB_X0Y164_IPAD),
.O(LIOB33_X0Y163_IOB_X0Y164_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y165_IOB_X0Y165_IBUF (
.I(LIOB33_X0Y165_IOB_X0Y165_IPAD),
.O(LIOB33_X0Y165_IOB_X0Y165_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y165_IOB_X0Y166_IBUF (
.I(LIOB33_X0Y165_IOB_X0Y166_IPAD),
.O(LIOB33_X0Y165_IOB_X0Y166_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y167_IOB_X0Y167_IBUF (
.I(LIOB33_X0Y167_IOB_X0Y167_IPAD),
.O(LIOB33_X0Y167_IOB_X0Y167_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y167_IOB_X0Y168_IBUF (
.I(LIOB33_X0Y167_IOB_X0Y168_IPAD),
.O(LIOB33_X0Y167_IOB_X0Y168_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y169_IOB_X0Y169_IBUF (
.I(LIOB33_X0Y169_IOB_X0Y169_IPAD),
.O(LIOB33_X0Y169_IOB_X0Y169_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y169_IOB_X0Y170_IBUF (
.I(LIOB33_X0Y169_IOB_X0Y170_IPAD),
.O(LIOB33_X0Y169_IOB_X0Y170_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y171_IOB_X0Y171_IBUF (
.I(LIOB33_X0Y171_IOB_X0Y171_IPAD),
.O(LIOB33_X0Y171_IOB_X0Y171_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y171_IOB_X0Y172_IBUF (
.I(LIOB33_X0Y171_IOB_X0Y172_IPAD),
.O(LIOB33_X0Y171_IOB_X0Y172_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y173_IOB_X0Y173_IBUF (
.I(LIOB33_X0Y173_IOB_X0Y173_IPAD),
.O(LIOB33_X0Y173_IOB_X0Y173_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y173_IOB_X0Y174_IBUF (
.I(LIOB33_X0Y173_IOB_X0Y174_IPAD),
.O(LIOB33_X0Y173_IOB_X0Y174_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y175_IOB_X0Y175_IBUF (
.I(LIOB33_X0Y175_IOB_X0Y175_IPAD),
.O(LIOB33_X0Y175_IOB_X0Y175_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y175_IOB_X0Y176_IBUF (
.I(LIOB33_X0Y175_IOB_X0Y176_IPAD),
.O(LIOB33_X0Y175_IOB_X0Y176_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y177_IOB_X0Y177_IBUF (
.I(LIOB33_X0Y177_IOB_X0Y177_IPAD),
.O(LIOB33_X0Y177_IOB_X0Y177_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y177_IOB_X0Y178_IBUF (
.I(LIOB33_X0Y177_IOB_X0Y178_IPAD),
.O(LIOB33_X0Y177_IOB_X0Y178_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y179_IOB_X0Y179_IBUF (
.I(LIOB33_X0Y179_IOB_X0Y179_IPAD),
.O(LIOB33_X0Y179_IOB_X0Y179_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y179_IOB_X0Y180_IBUF (
.I(LIOB33_X0Y179_IOB_X0Y180_IPAD),
.O(LIOB33_X0Y179_IOB_X0Y180_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y181_IOB_X0Y181_IBUF (
.I(LIOB33_X0Y181_IOB_X0Y181_IPAD),
.O(LIOB33_X0Y181_IOB_X0Y181_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y181_IOB_X0Y182_IBUF (
.I(LIOB33_X0Y181_IOB_X0Y182_IPAD),
.O(LIOB33_X0Y181_IOB_X0Y182_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y183_IOB_X0Y183_IBUF (
.I(LIOB33_X0Y183_IOB_X0Y183_IPAD),
.O(LIOB33_X0Y183_IOB_X0Y183_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y183_IOB_X0Y184_IBUF (
.I(LIOB33_X0Y183_IOB_X0Y184_IPAD),
.O(LIOB33_X0Y183_IOB_X0Y184_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y185_IOB_X0Y185_IBUF (
.I(LIOB33_X0Y185_IOB_X0Y185_IPAD),
.O(LIOB33_X0Y185_IOB_X0Y185_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y185_IOB_X0Y186_IBUF (
.I(LIOB33_X0Y185_IOB_X0Y186_IPAD),
.O(LIOB33_X0Y185_IOB_X0Y186_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y187_IOB_X0Y187_IBUF (
.I(LIOB33_X0Y187_IOB_X0Y187_IPAD),
.O(LIOB33_X0Y187_IOB_X0Y187_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y187_IOB_X0Y188_IBUF (
.I(LIOB33_X0Y187_IOB_X0Y188_IPAD),
.O(LIOB33_X0Y187_IOB_X0Y188_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y189_IOB_X0Y189_IBUF (
.I(LIOB33_X0Y189_IOB_X0Y189_IPAD),
.O(LIOB33_X0Y189_IOB_X0Y189_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y189_IOB_X0Y190_IBUF (
.I(LIOB33_X0Y189_IOB_X0Y190_IPAD),
.O(LIOB33_X0Y189_IOB_X0Y190_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y191_IOB_X0Y191_IBUF (
.I(LIOB33_X0Y191_IOB_X0Y191_IPAD),
.O(LIOB33_X0Y191_IOB_X0Y191_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y191_IOB_X0Y192_IBUF (
.I(LIOB33_X0Y191_IOB_X0Y192_IPAD),
.O(LIOB33_X0Y191_IOB_X0Y192_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y193_IOB_X0Y193_IBUF (
.I(LIOB33_X0Y193_IOB_X0Y193_IPAD),
.O(LIOB33_X0Y193_IOB_X0Y193_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y193_IOB_X0Y194_IBUF (
.I(LIOB33_X0Y193_IOB_X0Y194_IPAD),
.O(LIOB33_X0Y193_IOB_X0Y194_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y195_IOB_X0Y195_IBUF (
.I(LIOB33_X0Y195_IOB_X0Y195_IPAD),
.O(LIOB33_X0Y195_IOB_X0Y195_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y195_IOB_X0Y196_IBUF (
.I(LIOB33_X0Y195_IOB_X0Y196_IPAD),
.O(LIOB33_X0Y195_IOB_X0Y196_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y197_IOB_X0Y197_IBUF (
.I(LIOB33_X0Y197_IOB_X0Y197_IPAD),
.O(LIOB33_X0Y197_IOB_X0Y197_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y197_IOB_X0Y198_IBUF (
.I(LIOB33_X0Y197_IOB_X0Y198_IPAD),
.O(LIOB33_X0Y197_IOB_X0Y198_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y201_IOB_X0Y201_IBUF (
.I(LIOB33_X0Y201_IOB_X0Y201_IPAD),
.O(LIOB33_X0Y201_IOB_X0Y201_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y201_IOB_X0Y202_IBUF (
.I(LIOB33_X0Y201_IOB_X0Y202_IPAD),
.O(LIOB33_X0Y201_IOB_X0Y202_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y203_IOB_X0Y203_IBUF (
.I(LIOB33_X0Y203_IOB_X0Y203_IPAD),
.O(LIOB33_X0Y203_IOB_X0Y203_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y203_IOB_X0Y204_IBUF (
.I(LIOB33_X0Y203_IOB_X0Y204_IPAD),
.O(LIOB33_X0Y203_IOB_X0Y204_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y205_IOB_X0Y205_IBUF (
.I(LIOB33_X0Y205_IOB_X0Y205_IPAD),
.O(LIOB33_X0Y205_IOB_X0Y205_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y205_IOB_X0Y206_IBUF (
.I(LIOB33_X0Y205_IOB_X0Y206_IPAD),
.O(LIOB33_X0Y205_IOB_X0Y206_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y207_IOB_X0Y207_IBUF (
.I(LIOB33_X0Y207_IOB_X0Y207_IPAD),
.O(LIOB33_X0Y207_IOB_X0Y207_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y207_IOB_X0Y208_IBUF (
.I(LIOB33_X0Y207_IOB_X0Y208_IPAD),
.O(LIOB33_X0Y207_IOB_X0Y208_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y209_IOB_X0Y209_IBUF (
.I(LIOB33_X0Y209_IOB_X0Y209_IPAD),
.O(LIOB33_X0Y209_IOB_X0Y209_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y209_IOB_X0Y210_IBUF (
.I(LIOB33_X0Y209_IOB_X0Y210_IPAD),
.O(LIOB33_X0Y209_IOB_X0Y210_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y211_IOB_X0Y211_IBUF (
.I(LIOB33_X0Y211_IOB_X0Y211_IPAD),
.O(LIOB33_X0Y211_IOB_X0Y211_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y211_IOB_X0Y212_IBUF (
.I(LIOB33_X0Y211_IOB_X0Y212_IPAD),
.O(LIOB33_X0Y211_IOB_X0Y212_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y213_IOB_X0Y213_IBUF (
.I(LIOB33_X0Y213_IOB_X0Y213_IPAD),
.O(LIOB33_X0Y213_IOB_X0Y213_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y213_IOB_X0Y214_IBUF (
.I(LIOB33_X0Y213_IOB_X0Y214_IPAD),
.O(LIOB33_X0Y213_IOB_X0Y214_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y215_IOB_X0Y215_IBUF (
.I(LIOB33_X0Y215_IOB_X0Y215_IPAD),
.O(LIOB33_X0Y215_IOB_X0Y215_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y215_IOB_X0Y216_IBUF (
.I(LIOB33_X0Y215_IOB_X0Y216_IPAD),
.O(LIOB33_X0Y215_IOB_X0Y216_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y217_IOB_X0Y217_IBUF (
.I(LIOB33_X0Y217_IOB_X0Y217_IPAD),
.O(LIOB33_X0Y217_IOB_X0Y217_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y217_IOB_X0Y218_IBUF (
.I(LIOB33_X0Y217_IOB_X0Y218_IPAD),
.O(LIOB33_X0Y217_IOB_X0Y218_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y219_IOB_X0Y219_IBUF (
.I(LIOB33_X0Y219_IOB_X0Y219_IPAD),
.O(LIOB33_X0Y219_IOB_X0Y219_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y219_IOB_X0Y220_IBUF (
.I(LIOB33_X0Y219_IOB_X0Y220_IPAD),
.O(LIOB33_X0Y219_IOB_X0Y220_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y221_IOB_X0Y221_IBUF (
.I(LIOB33_X0Y221_IOB_X0Y221_IPAD),
.O(LIOB33_X0Y221_IOB_X0Y221_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y221_IOB_X0Y222_IBUF (
.I(LIOB33_X0Y221_IOB_X0Y222_IPAD),
.O(LIOB33_X0Y221_IOB_X0Y222_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y223_IOB_X0Y223_IBUF (
.I(LIOB33_X0Y223_IOB_X0Y223_IPAD),
.O(LIOB33_X0Y223_IOB_X0Y223_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y223_IOB_X0Y224_IBUF (
.I(LIOB33_X0Y223_IOB_X0Y224_IPAD),
.O(LIOB33_X0Y223_IOB_X0Y224_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y225_IOB_X0Y225_IBUF (
.I(LIOB33_X0Y225_IOB_X0Y225_IPAD),
.O(LIOB33_X0Y225_IOB_X0Y225_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y225_IOB_X0Y226_IBUF (
.I(LIOB33_X0Y225_IOB_X0Y226_IPAD),
.O(LIOB33_X0Y225_IOB_X0Y226_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y227_IOB_X0Y227_IBUF (
.I(LIOB33_X0Y227_IOB_X0Y227_IPAD),
.O(LIOB33_X0Y227_IOB_X0Y227_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y227_IOB_X0Y228_IBUF (
.I(LIOB33_X0Y227_IOB_X0Y228_IPAD),
.O(LIOB33_X0Y227_IOB_X0Y228_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y229_IOB_X0Y229_IBUF (
.I(LIOB33_X0Y229_IOB_X0Y229_IPAD),
.O(LIOB33_X0Y229_IOB_X0Y229_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y229_IOB_X0Y230_IBUF (
.I(LIOB33_X0Y229_IOB_X0Y230_IPAD),
.O(LIOB33_X0Y229_IOB_X0Y230_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y231_IOB_X0Y231_IBUF (
.I(LIOB33_X0Y231_IOB_X0Y231_IPAD),
.O(LIOB33_X0Y231_IOB_X0Y231_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y231_IOB_X0Y232_IBUF (
.I(LIOB33_X0Y231_IOB_X0Y232_IPAD),
.O(LIOB33_X0Y231_IOB_X0Y232_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y233_IOB_X0Y233_IBUF (
.I(LIOB33_X0Y233_IOB_X0Y233_IPAD),
.O(LIOB33_X0Y233_IOB_X0Y233_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y233_IOB_X0Y234_IBUF (
.I(LIOB33_X0Y233_IOB_X0Y234_IPAD),
.O(LIOB33_X0Y233_IOB_X0Y234_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y235_IOB_X0Y235_IBUF (
.I(LIOB33_X0Y235_IOB_X0Y235_IPAD),
.O(LIOB33_X0Y235_IOB_X0Y235_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y235_IOB_X0Y236_IBUF (
.I(LIOB33_X0Y235_IOB_X0Y236_IPAD),
.O(LIOB33_X0Y235_IOB_X0Y236_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y237_IOB_X0Y237_IBUF (
.I(LIOB33_X0Y237_IOB_X0Y237_IPAD),
.O(LIOB33_X0Y237_IOB_X0Y237_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y237_IOB_X0Y238_IBUF (
.I(LIOB33_X0Y237_IOB_X0Y238_IPAD),
.O(LIOB33_X0Y237_IOB_X0Y238_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y239_IOB_X0Y239_IBUF (
.I(LIOB33_X0Y239_IOB_X0Y239_IPAD),
.O(LIOB33_X0Y239_IOB_X0Y239_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y239_IOB_X0Y240_IBUF (
.I(LIOB33_X0Y239_IOB_X0Y240_IPAD),
.O(LIOB33_X0Y239_IOB_X0Y240_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y241_IOB_X0Y241_IBUF (
.I(LIOB33_X0Y241_IOB_X0Y241_IPAD),
.O(LIOB33_X0Y241_IOB_X0Y241_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y241_IOB_X0Y242_IBUF (
.I(LIOB33_X0Y241_IOB_X0Y242_IPAD),
.O(LIOB33_X0Y241_IOB_X0Y242_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y243_IOB_X0Y243_IBUF (
.I(LIOB33_X0Y243_IOB_X0Y243_IPAD),
.O(LIOB33_X0Y243_IOB_X0Y243_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y243_IOB_X0Y244_IBUF (
.I(LIOB33_X0Y243_IOB_X0Y244_IPAD),
.O(LIOB33_X0Y243_IOB_X0Y244_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y245_IOB_X0Y245_IBUF (
.I(LIOB33_X0Y245_IOB_X0Y245_IPAD),
.O(LIOB33_X0Y245_IOB_X0Y245_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y245_IOB_X0Y246_IBUF (
.I(LIOB33_X0Y245_IOB_X0Y246_IPAD),
.O(LIOB33_X0Y245_IOB_X0Y246_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y247_IOB_X0Y247_IBUF (
.I(LIOB33_X0Y247_IOB_X0Y247_IPAD),
.O(LIOB33_X0Y247_IOB_X0Y247_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y247_IOB_X0Y248_IBUF (
.I(LIOB33_X0Y247_IOB_X0Y248_IPAD),
.O(LIOB33_X0Y247_IOB_X0Y248_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y0_IOB_X0Y0_IBUF (
.I(LIOB33_SING_X0Y0_IOB_X0Y0_IPAD),
.O(LIOB33_SING_X0Y0_IOB_X0Y0_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y50_IOB_X0Y50_IBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_IPAD),
.O(LIOB33_SING_X0Y50_IOB_X0Y50_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y99_IOB_X0Y99_IBUF (
.I(LIOB33_SING_X0Y99_IOB_X0Y99_IPAD),
.O(LIOB33_SING_X0Y99_IOB_X0Y99_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y100_IOB_X0Y100_OBUF (
.I(CLBLL_L_X2Y141_SLICE_X0Y141_AQ),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y149_IOB_X0Y149_IBUF (
.I(LIOB33_SING_X0Y149_IOB_X0Y149_IPAD),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y150_IOB_X0Y150_IBUF (
.I(LIOB33_SING_X0Y150_IOB_X0Y150_IPAD),
.O(LIOB33_SING_X0Y150_IOB_X0Y150_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y199_IOB_X0Y199_IBUF (
.I(LIOB33_SING_X0Y199_IOB_X0Y199_IPAD),
.O(LIOB33_SING_X0Y199_IOB_X0Y199_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y200_IOB_X0Y200_IBUF (
.I(LIOB33_SING_X0Y200_IOB_X0Y200_IPAD),
.O(LIOB33_SING_X0Y200_IOB_X0Y200_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y249_IOB_X0Y249_IBUF (
.I(LIOB33_SING_X0Y249_IOB_X0Y249_IPAD),
.O(LIOB33_SING_X0Y249_IOB_X0Y249_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y51_IOB_X1Y51_OBUF (
.I(CLBLM_R_X5Y132_SLICE_X7Y132_BQ),
.O(RIOB33_X105Y51_IOB_X1Y51_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y51_IOB_X1Y52_OBUF (
.I(CLBLM_R_X5Y134_SLICE_X7Y134_CQ),
.O(RIOB33_X105Y51_IOB_X1Y52_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y53_IOB_X1Y53_OBUF (
.I(CLBLM_L_X8Y131_SLICE_X10Y131_AQ),
.O(RIOB33_X105Y53_IOB_X1Y53_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y53_IOB_X1Y54_OBUF (
.I(CLBLM_R_X7Y132_SLICE_X9Y132_AQ),
.O(RIOB33_X105Y53_IOB_X1Y54_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y55_IOB_X1Y55_OBUF (
.I(CLBLL_L_X4Y134_SLICE_X5Y134_AQ),
.O(RIOB33_X105Y55_IOB_X1Y55_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y55_IOB_X1Y56_OBUF (
.I(CLBLM_R_X5Y133_SLICE_X7Y133_CQ),
.O(RIOB33_X105Y55_IOB_X1Y56_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y57_IOB_X1Y57_OBUF (
.I(CLBLM_R_X7Y137_SLICE_X9Y137_CQ),
.O(RIOB33_X105Y57_IOB_X1Y57_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y57_IOB_X1Y58_OBUF (
.I(CLBLM_L_X8Y130_SLICE_X10Y130_CQ),
.O(RIOB33_X105Y57_IOB_X1Y58_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y59_IOB_X1Y59_OBUF (
.I(CLBLM_R_X5Y131_SLICE_X6Y131_AQ),
.O(RIOB33_X105Y59_IOB_X1Y59_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y59_IOB_X1Y60_OBUF (
.I(CLBLM_R_X7Y136_SLICE_X8Y136_BQ),
.O(RIOB33_X105Y59_IOB_X1Y60_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y61_IOB_X1Y61_OBUF (
.I(CLBLL_L_X4Y135_SLICE_X5Y135_BQ),
.O(RIOB33_X105Y61_IOB_X1Y61_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y61_IOB_X1Y62_OBUF (
.I(CLBLL_L_X4Y134_SLICE_X5Y134_BQ),
.O(RIOB33_X105Y61_IOB_X1Y62_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y63_IOB_X1Y63_OBUF (
.I(CLBLM_R_X7Y137_SLICE_X9Y137_DQ),
.O(RIOB33_X105Y63_IOB_X1Y63_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y63_IOB_X1Y64_OBUF (
.I(CLBLL_L_X54Y96_SLICE_X82Y96_AQ),
.O(RIOB33_X105Y63_IOB_X1Y64_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y65_IOB_X1Y65_OBUF (
.I(CLBLM_L_X8Y127_SLICE_X10Y127_AQ),
.O(RIOB33_X105Y65_IOB_X1Y65_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y65_IOB_X1Y66_OBUF (
.I(CLBLM_R_X7Y125_SLICE_X8Y125_AQ),
.O(RIOB33_X105Y65_IOB_X1Y66_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y67_IOB_X1Y67_OBUF (
.I(CLBLM_L_X8Y127_SLICE_X10Y127_BQ),
.O(RIOB33_X105Y67_IOB_X1Y67_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y67_IOB_X1Y68_OBUF (
.I(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.O(RIOB33_X105Y67_IOB_X1Y68_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y69_IOB_X1Y69_OBUF (
.I(CLBLM_L_X8Y129_SLICE_X10Y129_BQ),
.O(RIOB33_X105Y69_IOB_X1Y69_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y69_IOB_X1Y70_OBUF (
.I(CLBLM_L_X8Y129_SLICE_X10Y129_CQ),
.O(RIOB33_X105Y69_IOB_X1Y70_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y71_IOB_X1Y71_OBUF (
.I(CLBLL_L_X54Y101_SLICE_X82Y101_AQ),
.O(RIOB33_X105Y71_IOB_X1Y71_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y71_IOB_X1Y72_OBUF (
.I(CLBLM_R_X7Y128_SLICE_X9Y128_AQ),
.O(RIOB33_X105Y71_IOB_X1Y72_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y73_IOB_X1Y73_OBUF (
.I(CLBLM_L_X8Y130_SLICE_X11Y130_BQ),
.O(RIOB33_X105Y73_IOB_X1Y73_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y73_IOB_X1Y74_OBUF (
.I(CLBLM_R_X7Y130_SLICE_X9Y130_DQ),
.O(RIOB33_X105Y73_IOB_X1Y74_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y75_IOB_X1Y75_OBUF (
.I(CLBLM_L_X8Y130_SLICE_X10Y130_DQ),
.O(RIOB33_X105Y75_IOB_X1Y75_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y75_IOB_X1Y76_OBUF (
.I(CLBLM_L_X10Y132_SLICE_X12Y132_AQ),
.O(RIOB33_X105Y75_IOB_X1Y76_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y77_IOB_X1Y77_OBUF (
.I(CLBLM_L_X8Y130_SLICE_X11Y130_CQ),
.O(RIOB33_X105Y77_IOB_X1Y77_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y77_IOB_X1Y78_OBUF (
.I(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.O(RIOB33_X105Y77_IOB_X1Y78_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y79_IOB_X1Y79_OBUF (
.I(CLBLL_L_X54Y105_SLICE_X82Y105_AQ),
.O(RIOB33_X105Y79_IOB_X1Y79_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y79_IOB_X1Y80_OBUF (
.I(CLBLM_L_X8Y131_SLICE_X11Y131_BQ),
.O(RIOB33_X105Y79_IOB_X1Y80_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y81_IOB_X1Y81_OBUF (
.I(CLBLM_L_X8Y131_SLICE_X11Y131_CQ),
.O(RIOB33_X105Y81_IOB_X1Y81_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y81_IOB_X1Y82_OBUF (
.I(CLBLM_L_X8Y130_SLICE_X11Y130_DQ),
.O(RIOB33_X105Y81_IOB_X1Y82_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y83_IOB_X1Y83_OBUF (
.I(CLBLM_L_X8Y131_SLICE_X10Y131_BQ),
.O(RIOB33_X105Y83_IOB_X1Y83_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y83_IOB_X1Y84_OBUF (
.I(CLBLM_L_X10Y132_SLICE_X12Y132_BQ),
.O(RIOB33_X105Y83_IOB_X1Y84_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y85_IOB_X1Y85_OBUF (
.I(CLBLM_L_X10Y132_SLICE_X12Y132_CQ),
.O(RIOB33_X105Y85_IOB_X1Y85_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y85_IOB_X1Y86_OBUF (
.I(CLBLM_L_X8Y132_SLICE_X11Y132_CQ),
.O(RIOB33_X105Y85_IOB_X1Y86_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y87_IOB_X1Y87_OBUF (
.I(CLBLM_L_X10Y132_SLICE_X12Y132_DQ),
.O(RIOB33_X105Y87_IOB_X1Y87_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y87_IOB_X1Y88_OBUF (
.I(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.O(RIOB33_X105Y87_IOB_X1Y88_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y89_IOB_X1Y89_OBUF (
.I(CLBLM_R_X11Y130_SLICE_X14Y130_AQ),
.O(RIOB33_X105Y89_IOB_X1Y89_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y89_IOB_X1Y90_OBUF (
.I(CLBLM_L_X10Y130_SLICE_X12Y130_BQ),
.O(RIOB33_X105Y89_IOB_X1Y90_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y91_IOB_X1Y91_OBUF (
.I(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.O(RIOB33_X105Y91_IOB_X1Y91_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y91_IOB_X1Y92_OBUF (
.I(CLBLM_R_X11Y131_SLICE_X14Y131_AQ),
.O(RIOB33_X105Y91_IOB_X1Y92_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y93_IOB_X1Y93_OBUF (
.I(CLBLM_L_X12Y132_SLICE_X16Y132_CQ),
.O(RIOB33_X105Y93_IOB_X1Y93_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y93_IOB_X1Y94_OBUF (
.I(CLBLM_L_X10Y131_SLICE_X13Y131_AQ),
.O(RIOB33_X105Y93_IOB_X1Y94_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y95_IOB_X1Y95_OBUF (
.I(CLBLM_R_X11Y131_SLICE_X14Y131_BQ),
.O(RIOB33_X105Y95_IOB_X1Y95_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y95_IOB_X1Y96_OBUF (
.I(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.O(RIOB33_X105Y95_IOB_X1Y96_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y97_IOB_X1Y97_OBUF (
.I(CLBLM_R_X7Y125_SLICE_X8Y125_BQ),
.O(RIOB33_X105Y97_IOB_X1Y97_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y97_IOB_X1Y98_OBUF (
.I(CLBLM_R_X7Y125_SLICE_X8Y125_CQ),
.O(RIOB33_X105Y97_IOB_X1Y98_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y101_IOB_X1Y101_OBUF (
.I(CLBLM_R_X7Y126_SLICE_X8Y126_AQ),
.O(RIOB33_X105Y101_IOB_X1Y101_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y101_IOB_X1Y102_OBUF (
.I(CLBLM_R_X7Y126_SLICE_X8Y126_BQ),
.O(RIOB33_X105Y101_IOB_X1Y102_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y103_IOB_X1Y103_OBUF (
.I(CLBLM_R_X7Y126_SLICE_X8Y126_CQ),
.O(RIOB33_X105Y103_IOB_X1Y103_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y103_IOB_X1Y104_OBUF (
.I(CLBLM_R_X7Y128_SLICE_X8Y128_BQ),
.O(RIOB33_X105Y103_IOB_X1Y104_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y105_IOB_X1Y105_OBUF (
.I(CLBLM_R_X7Y129_SLICE_X9Y129_CQ),
.O(RIOB33_X105Y105_IOB_X1Y105_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y105_IOB_X1Y106_OBUF (
.I(CLBLM_R_X5Y131_SLICE_X7Y131_AQ),
.O(RIOB33_X105Y105_IOB_X1Y106_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y107_IOB_X1Y107_OBUF (
.I(CLBLL_L_X54Y119_SLICE_X82Y119_AQ),
.O(RIOB33_X105Y107_IOB_X1Y107_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y107_IOB_X1Y108_OBUF (
.I(CLBLM_R_X7Y130_SLICE_X8Y130_BQ),
.O(RIOB33_X105Y107_IOB_X1Y108_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y109_IOB_X1Y109_OBUF (
.I(CLBLM_R_X7Y129_SLICE_X8Y129_CQ),
.O(RIOB33_X105Y109_IOB_X1Y109_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y109_IOB_X1Y110_OBUF (
.I(CLBLM_R_X7Y129_SLICE_X8Y129_DQ),
.O(RIOB33_X105Y109_IOB_X1Y110_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y111_IOB_X1Y111_OBUF (
.I(CLBLM_R_X7Y130_SLICE_X9Y130_AQ),
.O(RIOB33_X105Y111_IOB_X1Y111_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y111_IOB_X1Y112_OBUF (
.I(CLBLM_R_X7Y131_SLICE_X9Y131_BQ),
.O(RIOB33_X105Y111_IOB_X1Y112_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y113_IOB_X1Y113_OBUF (
.I(CLBLM_R_X7Y131_SLICE_X9Y131_CQ),
.O(RIOB33_X105Y113_IOB_X1Y113_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y113_IOB_X1Y114_OBUF (
.I(CLBLM_R_X7Y131_SLICE_X9Y131_DQ),
.O(RIOB33_X105Y113_IOB_X1Y114_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y115_IOB_X1Y115_OBUF (
.I(CLBLL_L_X54Y123_SLICE_X82Y123_AQ),
.O(RIOB33_X105Y115_IOB_X1Y115_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y115_IOB_X1Y116_OBUF (
.I(CLBLM_L_X10Y133_SLICE_X13Y133_AQ),
.O(RIOB33_X105Y115_IOB_X1Y116_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y117_IOB_X1Y117_OBUF (
.I(CLBLM_L_X12Y132_SLICE_X16Y132_AQ),
.O(RIOB33_X105Y117_IOB_X1Y117_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y117_IOB_X1Y118_OBUF (
.I(CLBLM_L_X10Y131_SLICE_X12Y131_AQ),
.O(RIOB33_X105Y117_IOB_X1Y118_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y119_IOB_X1Y119_OBUF (
.I(CLBLM_R_X11Y133_SLICE_X14Y133_AQ),
.O(RIOB33_X105Y119_IOB_X1Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y119_IOB_X1Y120_OBUF (
.I(CLBLM_L_X10Y133_SLICE_X13Y133_BQ),
.O(RIOB33_X105Y119_IOB_X1Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y121_IOB_X1Y121_OBUF (
.I(CLBLM_R_X11Y133_SLICE_X14Y133_BQ),
.O(RIOB33_X105Y121_IOB_X1Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y121_IOB_X1Y122_OBUF (
.I(CLBLM_L_X10Y133_SLICE_X13Y133_CQ),
.O(RIOB33_X105Y121_IOB_X1Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y123_IOB_X1Y123_OBUF (
.I(CLBLM_L_X12Y132_SLICE_X16Y132_BQ),
.O(RIOB33_X105Y123_IOB_X1Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y123_IOB_X1Y124_OBUF (
.I(CLBLM_R_X7Y130_SLICE_X9Y130_BQ),
.O(RIOB33_X105Y123_IOB_X1Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y125_IOB_X1Y125_OBUF (
.I(CLBLM_R_X5Y132_SLICE_X7Y132_AQ),
.O(RIOB33_X105Y125_IOB_X1Y125_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y125_IOB_X1Y126_OBUF (
.I(CLBLM_R_X7Y130_SLICE_X9Y130_CQ),
.O(RIOB33_X105Y125_IOB_X1Y126_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y127_IOB_X1Y127_OBUF (
.I(CLBLM_R_X5Y133_SLICE_X7Y133_AQ),
.O(RIOB33_X105Y127_IOB_X1Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y127_IOB_X1Y128_OBUF (
.I(CLBLM_L_X8Y134_SLICE_X10Y134_AQ),
.O(RIOB33_X105Y127_IOB_X1Y128_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y129_IOB_X1Y129_OBUF (
.I(CLBLM_R_X7Y133_SLICE_X9Y133_AQ),
.O(RIOB33_X105Y129_IOB_X1Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y129_IOB_X1Y130_OBUF (
.I(CLBLM_L_X8Y132_SLICE_X11Y132_BQ),
.O(RIOB33_X105Y129_IOB_X1Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y131_IOB_X1Y131_OBUF (
.I(CLBLM_R_X5Y134_SLICE_X7Y134_BQ),
.O(RIOB33_X105Y131_IOB_X1Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y131_IOB_X1Y132_OBUF (
.I(CLBLL_L_X54Y133_SLICE_X82Y133_AQ),
.O(RIOB33_X105Y131_IOB_X1Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y133_IOB_X1Y133_OBUF (
.I(CLBLM_R_X7Y133_SLICE_X9Y133_BQ),
.O(RIOB33_X105Y133_IOB_X1Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y133_IOB_X1Y134_OBUF (
.I(CLBLM_R_X5Y133_SLICE_X7Y133_BQ),
.O(RIOB33_X105Y133_IOB_X1Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y135_IOB_X1Y135_OBUF (
.I(CLBLM_R_X7Y137_SLICE_X9Y137_AQ),
.O(RIOB33_X105Y135_IOB_X1Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y135_IOB_X1Y136_OBUF (
.I(CLBLM_R_X5Y135_SLICE_X7Y135_AQ),
.O(RIOB33_X105Y135_IOB_X1Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y137_IOB_X1Y137_OBUF (
.I(CLBLM_R_X5Y137_SLICE_X7Y137_AQ),
.O(RIOB33_X105Y137_IOB_X1Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y137_IOB_X1Y138_OBUF (
.I(CLBLM_R_X7Y137_SLICE_X8Y137_BQ),
.O(RIOB33_X105Y137_IOB_X1Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y139_IOB_X1Y139_OBUF (
.I(CLBLL_L_X54Y138_SLICE_X82Y138_AQ),
.O(RIOB33_X105Y139_IOB_X1Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y139_IOB_X1Y140_OBUF (
.I(CLBLM_R_X7Y138_SLICE_X9Y138_AQ),
.O(RIOB33_X105Y139_IOB_X1Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y141_IOB_X1Y141_OBUF (
.I(CLBLM_R_X7Y138_SLICE_X9Y138_BQ),
.O(RIOB33_X105Y141_IOB_X1Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y141_IOB_X1Y142_OBUF (
.I(CLBLM_R_X7Y138_SLICE_X9Y138_CQ),
.O(RIOB33_X105Y141_IOB_X1Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y143_IOB_X1Y143_OBUF (
.I(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.O(RIOB33_X105Y143_IOB_X1Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y143_IOB_X1Y144_OBUF (
.I(CLBLM_R_X5Y138_SLICE_X6Y138_AQ),
.O(RIOB33_X105Y143_IOB_X1Y144_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y145_IOB_X1Y145_OBUF (
.I(CLBLM_R_X5Y138_SLICE_X6Y138_BQ),
.O(RIOB33_X105Y145_IOB_X1Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y145_IOB_X1Y146_OBUF (
.I(CLBLM_R_X5Y138_SLICE_X7Y138_AQ),
.O(RIOB33_X105Y145_IOB_X1Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y147_IOB_X1Y147_OBUF (
.I(CLBLL_L_X54Y141_SLICE_X82Y141_AQ),
.O(RIOB33_X105Y147_IOB_X1Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y147_IOB_X1Y148_OBUF (
.I(CLBLM_R_X7Y137_SLICE_X9Y137_BQ),
.O(RIOB33_X105Y147_IOB_X1Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y151_OBUF (
.I(CLBLM_R_X7Y128_SLICE_X8Y128_AQ),
.O(RIOB33_X105Y151_IOB_X1Y151_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y152_OBUF (
.I(CLBLM_R_X7Y129_SLICE_X9Y129_BQ),
.O(RIOB33_X105Y151_IOB_X1Y152_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y153_OBUF (
.I(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.O(RIOB33_X105Y153_IOB_X1Y153_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y154_OBUF (
.I(CLBLM_R_X7Y129_SLICE_X8Y129_AQ),
.O(RIOB33_X105Y153_IOB_X1Y154_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y155_OBUF (
.I(CLBLM_R_X7Y136_SLICE_X8Y136_AQ),
.O(RIOB33_X105Y155_IOB_X1Y155_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y156_OBUF (
.I(CLBLM_R_X7Y129_SLICE_X8Y129_BQ),
.O(RIOB33_X105Y155_IOB_X1Y156_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y157_OBUF (
.I(CLBLM_L_X8Y130_SLICE_X10Y130_BQ),
.O(RIOB33_X105Y157_IOB_X1Y157_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y158_OBUF (
.I(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.O(RIOB33_X105Y157_IOB_X1Y158_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y159_OBUF (
.I(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.O(RIOB33_X105Y159_IOB_X1Y159_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y160_OBUF (
.I(CLBLM_R_X7Y137_SLICE_X8Y137_AQ),
.O(RIOB33_X105Y159_IOB_X1Y160_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y161_OBUF (
.I(CLBLM_R_X5Y134_SLICE_X7Y134_AQ),
.O(RIOB33_X105Y161_IOB_X1Y161_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y162_OBUF (
.I(CLBLM_L_X8Y132_SLICE_X11Y132_AQ),
.O(RIOB33_X105Y161_IOB_X1Y162_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y163_OBUF (
.I(CLBLM_L_X8Y135_SLICE_X10Y135_AQ),
.O(RIOB33_X105Y163_IOB_X1Y163_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y164_OBUF (
.I(CLBLM_R_X7Y134_SLICE_X9Y134_AQ),
.O(RIOB33_X105Y163_IOB_X1Y164_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y165_OBUF (
.I(CLBLM_R_X7Y134_SLICE_X9Y134_BQ),
.O(RIOB33_X105Y165_IOB_X1Y165_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y166_OBUF (
.I(CLBLM_L_X8Y136_SLICE_X10Y136_AQ),
.O(RIOB33_X105Y165_IOB_X1Y166_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y167_OBUF (
.I(CLBLM_L_X10Y135_SLICE_X12Y135_AQ),
.O(RIOB33_X105Y167_IOB_X1Y167_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y168_OBUF (
.I(CLBLM_L_X8Y137_SLICE_X10Y137_AQ),
.O(RIOB33_X105Y167_IOB_X1Y168_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y169_OBUF (
.I(CLBLM_L_X8Y137_SLICE_X10Y137_BQ),
.O(RIOB33_X105Y169_IOB_X1Y169_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y170_OBUF (
.I(CLBLM_L_X56Y151_SLICE_X84Y151_AQ),
.O(RIOB33_X105Y169_IOB_X1Y170_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y171_OBUF (
.I(CLBLM_R_X15Y135_SLICE_X21Y135_AQ),
.O(RIOB33_X105Y171_IOB_X1Y171_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y172_OBUF (
.I(CLBLM_L_X16Y136_SLICE_X22Y136_AQ),
.O(RIOB33_X105Y171_IOB_X1Y172_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y173_OBUF (
.I(CLBLM_L_X16Y135_SLICE_X22Y135_AQ),
.O(RIOB33_X105Y173_IOB_X1Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y174_OBUF (
.I(CLBLM_L_X16Y135_SLICE_X22Y135_BQ),
.O(RIOB33_X105Y173_IOB_X1Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y175_OBUF (
.I(CLBLM_R_X13Y136_SLICE_X18Y136_AQ),
.O(RIOB33_X105Y175_IOB_X1Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y176_OBUF (
.I(CLBLM_L_X16Y137_SLICE_X22Y137_AQ),
.O(RIOB33_X105Y175_IOB_X1Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y177_OBUF (
.I(CLBLM_L_X16Y137_SLICE_X22Y137_BQ),
.O(RIOB33_X105Y177_IOB_X1Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y177_IOB_X1Y178_IBUF (
.I(RIOB33_X105Y177_IOB_X1Y178_IPAD),
.O(RIOB33_X105Y177_IOB_X1Y178_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y179_IOB_X1Y179_IBUF (
.I(RIOB33_X105Y179_IOB_X1Y179_IPAD),
.O(RIOB33_X105Y179_IOB_X1Y179_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y179_IOB_X1Y180_IBUF (
.I(RIOB33_X105Y179_IOB_X1Y180_IPAD),
.O(RIOB33_X105Y179_IOB_X1Y180_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y181_IOB_X1Y181_IBUF (
.I(RIOB33_X105Y181_IOB_X1Y181_IPAD),
.O(RIOB33_X105Y181_IOB_X1Y181_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y181_IOB_X1Y182_IBUF (
.I(RIOB33_X105Y181_IOB_X1Y182_IPAD),
.O(RIOB33_X105Y181_IOB_X1Y182_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y183_IOB_X1Y183_IBUF (
.I(RIOB33_X105Y183_IOB_X1Y183_IPAD),
.O(RIOB33_X105Y183_IOB_X1Y183_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y183_IOB_X1Y184_IBUF (
.I(RIOB33_X105Y183_IOB_X1Y184_IPAD),
.O(RIOB33_X105Y183_IOB_X1Y184_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y185_IOB_X1Y185_IBUF (
.I(RIOB33_X105Y185_IOB_X1Y185_IPAD),
.O(RIOB33_X105Y185_IOB_X1Y185_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y185_IOB_X1Y186_IBUF (
.I(RIOB33_X105Y185_IOB_X1Y186_IPAD),
.O(RIOB33_X105Y185_IOB_X1Y186_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y187_IOB_X1Y187_IBUF (
.I(RIOB33_X105Y187_IOB_X1Y187_IPAD),
.O(RIOB33_X105Y187_IOB_X1Y187_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y187_IOB_X1Y188_IBUF (
.I(RIOB33_X105Y187_IOB_X1Y188_IPAD),
.O(RIOB33_X105Y187_IOB_X1Y188_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y189_IOB_X1Y189_IBUF (
.I(RIOB33_X105Y189_IOB_X1Y189_IPAD),
.O(RIOB33_X105Y189_IOB_X1Y189_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y189_IOB_X1Y190_IBUF (
.I(RIOB33_X105Y189_IOB_X1Y190_IPAD),
.O(RIOB33_X105Y189_IOB_X1Y190_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y191_IOB_X1Y191_IBUF (
.I(RIOB33_X105Y191_IOB_X1Y191_IPAD),
.O(RIOB33_X105Y191_IOB_X1Y191_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y191_IOB_X1Y192_IBUF (
.I(RIOB33_X105Y191_IOB_X1Y192_IPAD),
.O(RIOB33_X105Y191_IOB_X1Y192_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y193_IOB_X1Y193_IBUF (
.I(RIOB33_X105Y193_IOB_X1Y193_IPAD),
.O(RIOB33_X105Y193_IOB_X1Y193_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y193_IOB_X1Y194_IBUF (
.I(RIOB33_X105Y193_IOB_X1Y194_IPAD),
.O(RIOB33_X105Y193_IOB_X1Y194_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y195_IOB_X1Y195_IBUF (
.I(RIOB33_X105Y195_IOB_X1Y195_IPAD),
.O(RIOB33_X105Y195_IOB_X1Y195_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y195_IOB_X1Y196_IBUF (
.I(RIOB33_X105Y195_IOB_X1Y196_IPAD),
.O(RIOB33_X105Y195_IOB_X1Y196_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y197_IOB_X1Y197_IBUF (
.I(RIOB33_X105Y197_IOB_X1Y197_IPAD),
.O(RIOB33_X105Y197_IOB_X1Y197_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y197_IOB_X1Y198_IBUF (
.I(RIOB33_X105Y197_IOB_X1Y198_IPAD),
.O(RIOB33_X105Y197_IOB_X1Y198_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y201_IOB_X1Y201_IBUF (
.I(RIOB33_X105Y201_IOB_X1Y201_IPAD),
.O(RIOB33_X105Y201_IOB_X1Y201_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y201_IOB_X1Y202_IBUF (
.I(RIOB33_X105Y201_IOB_X1Y202_IPAD),
.O(RIOB33_X105Y201_IOB_X1Y202_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y203_IOB_X1Y203_IBUF (
.I(RIOB33_X105Y203_IOB_X1Y203_IPAD),
.O(RIOB33_X105Y203_IOB_X1Y203_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y203_IOB_X1Y204_IBUF (
.I(RIOB33_X105Y203_IOB_X1Y204_IPAD),
.O(RIOB33_X105Y203_IOB_X1Y204_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y205_IOB_X1Y205_IBUF (
.I(RIOB33_X105Y205_IOB_X1Y205_IPAD),
.O(RIOB33_X105Y205_IOB_X1Y205_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y50_IOB_X1Y50_OBUF (
.I(CLBLM_R_X5Y130_SLICE_X7Y130_AQ),
.O(RIOB33_SING_X105Y50_IOB_X1Y50_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y99_IOB_X1Y99_OBUF (
.I(CLBLM_R_X7Y126_SLICE_X8Y126_DQ),
.O(RIOB33_SING_X105Y99_IOB_X1Y99_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y100_IOB_X1Y100_OBUF (
.I(CLBLL_L_X54Y116_SLICE_X82Y116_AQ),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y149_IOB_X1Y149_OBUF (
.I(CLBLM_R_X7Y138_SLICE_X9Y138_DQ),
.O(RIOB33_SING_X105Y149_IOB_X1Y149_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y150_IOB_X1Y150_OBUF (
.I(CLBLM_R_X7Y129_SLICE_X9Y129_AQ),
.O(RIOB33_SING_X105Y150_IOB_X1Y150_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y199_IOB_X1Y199_IBUF (
.I(RIOB33_SING_X105Y199_IOB_X1Y199_IPAD),
.O(RIOB33_SING_X105Y199_IOB_X1Y199_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y200_IOB_X1Y200_IBUF (
.I(RIOB33_SING_X105Y200_IOB_X1Y200_IPAD),
.O(RIOB33_SING_X105Y200_IOB_X1Y200_I)
  );
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A = CLBLL_L_X2Y131_SLICE_X0Y131_AO6;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B = CLBLL_L_X2Y131_SLICE_X0Y131_BO6;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C = CLBLL_L_X2Y131_SLICE_X0Y131_CO6;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D = CLBLL_L_X2Y131_SLICE_X0Y131_DO6;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A = CLBLL_L_X2Y131_SLICE_X1Y131_AO6;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B = CLBLL_L_X2Y131_SLICE_X1Y131_BO6;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C = CLBLL_L_X2Y131_SLICE_X1Y131_CO6;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D = CLBLL_L_X2Y131_SLICE_X1Y131_DO6;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_AMUX = CLBLL_L_X2Y131_SLICE_X1Y131_A5Q;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_A = CLBLL_L_X2Y132_SLICE_X0Y132_AO6;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_B = CLBLL_L_X2Y132_SLICE_X0Y132_BO6;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_C = CLBLL_L_X2Y132_SLICE_X0Y132_CO6;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_D = CLBLL_L_X2Y132_SLICE_X0Y132_DO6;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_A = CLBLL_L_X2Y132_SLICE_X1Y132_AO6;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_B = CLBLL_L_X2Y132_SLICE_X1Y132_BO6;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_C = CLBLL_L_X2Y132_SLICE_X1Y132_CO6;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_D = CLBLL_L_X2Y132_SLICE_X1Y132_DO6;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_A = CLBLL_L_X2Y141_SLICE_X0Y141_AO6;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_B = CLBLL_L_X2Y141_SLICE_X0Y141_BO6;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_C = CLBLL_L_X2Y141_SLICE_X0Y141_CO6;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_D = CLBLL_L_X2Y141_SLICE_X0Y141_DO6;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_A = CLBLL_L_X2Y141_SLICE_X1Y141_AO6;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_B = CLBLL_L_X2Y141_SLICE_X1Y141_BO6;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_C = CLBLL_L_X2Y141_SLICE_X1Y141_CO6;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_D = CLBLL_L_X2Y141_SLICE_X1Y141_DO6;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_A = CLBLL_L_X2Y142_SLICE_X0Y142_AO6;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_B = CLBLL_L_X2Y142_SLICE_X0Y142_BO6;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_C = CLBLL_L_X2Y142_SLICE_X0Y142_CO6;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_D = CLBLL_L_X2Y142_SLICE_X0Y142_DO6;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_A = CLBLL_L_X2Y142_SLICE_X1Y142_AO6;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_B = CLBLL_L_X2Y142_SLICE_X1Y142_BO6;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_C = CLBLL_L_X2Y142_SLICE_X1Y142_CO6;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_D = CLBLL_L_X2Y142_SLICE_X1Y142_DO6;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_A = CLBLL_L_X2Y152_SLICE_X0Y152_AO6;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_B = CLBLL_L_X2Y152_SLICE_X0Y152_BO6;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_C = CLBLL_L_X2Y152_SLICE_X0Y152_CO6;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_D = CLBLL_L_X2Y152_SLICE_X0Y152_DO6;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_A = CLBLL_L_X2Y152_SLICE_X1Y152_AO6;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_B = CLBLL_L_X2Y152_SLICE_X1Y152_BO6;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_C = CLBLL_L_X2Y152_SLICE_X1Y152_CO6;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_D = CLBLL_L_X2Y152_SLICE_X1Y152_DO6;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_A = CLBLL_L_X2Y155_SLICE_X0Y155_AO6;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_B = CLBLL_L_X2Y155_SLICE_X0Y155_BO6;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_C = CLBLL_L_X2Y155_SLICE_X0Y155_CO6;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_D = CLBLL_L_X2Y155_SLICE_X0Y155_DO6;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_A = CLBLL_L_X2Y155_SLICE_X1Y155_AO6;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_B = CLBLL_L_X2Y155_SLICE_X1Y155_BO6;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_C = CLBLL_L_X2Y155_SLICE_X1Y155_CO6;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_D = CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_A = CLBLL_L_X2Y157_SLICE_X0Y157_AO6;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_B = CLBLL_L_X2Y157_SLICE_X0Y157_BO6;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_C = CLBLL_L_X2Y157_SLICE_X0Y157_CO6;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_D = CLBLL_L_X2Y157_SLICE_X0Y157_DO6;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_A = CLBLL_L_X2Y157_SLICE_X1Y157_AO6;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_B = CLBLL_L_X2Y157_SLICE_X1Y157_BO6;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_C = CLBLL_L_X2Y157_SLICE_X1Y157_CO6;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_D = CLBLL_L_X2Y157_SLICE_X1Y157_DO6;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_A = CLBLL_L_X2Y158_SLICE_X0Y158_AO6;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_B = CLBLL_L_X2Y158_SLICE_X0Y158_BO6;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_C = CLBLL_L_X2Y158_SLICE_X0Y158_CO6;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_D = CLBLL_L_X2Y158_SLICE_X0Y158_DO6;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_A = CLBLL_L_X2Y158_SLICE_X1Y158_AO6;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_B = CLBLL_L_X2Y158_SLICE_X1Y158_BO6;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_C = CLBLL_L_X2Y158_SLICE_X1Y158_CO6;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_D = CLBLL_L_X2Y158_SLICE_X1Y158_DO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A = CLBLL_L_X4Y127_SLICE_X4Y127_AO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B = CLBLL_L_X4Y127_SLICE_X4Y127_BO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C = CLBLL_L_X4Y127_SLICE_X4Y127_CO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D = CLBLL_L_X4Y127_SLICE_X4Y127_DO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A = CLBLL_L_X4Y127_SLICE_X5Y127_AO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B = CLBLL_L_X4Y127_SLICE_X5Y127_BO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C = CLBLL_L_X4Y127_SLICE_X5Y127_CO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D = CLBLL_L_X4Y127_SLICE_X5Y127_DO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_A = CLBLL_L_X4Y128_SLICE_X4Y128_AO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_B = CLBLL_L_X4Y128_SLICE_X4Y128_BO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_C = CLBLL_L_X4Y128_SLICE_X4Y128_CO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_D = CLBLL_L_X4Y128_SLICE_X4Y128_DO6;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_A = CLBLL_L_X4Y128_SLICE_X5Y128_AO6;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_B = CLBLL_L_X4Y128_SLICE_X5Y128_BO6;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_C = CLBLL_L_X4Y128_SLICE_X5Y128_CO6;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_D = CLBLL_L_X4Y128_SLICE_X5Y128_DO6;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_AMUX = CLBLL_L_X4Y128_SLICE_X5Y128_AO5;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A = CLBLL_L_X4Y129_SLICE_X4Y129_AO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B = CLBLL_L_X4Y129_SLICE_X4Y129_BO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C = CLBLL_L_X4Y129_SLICE_X4Y129_CO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D = CLBLL_L_X4Y129_SLICE_X4Y129_DO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A = CLBLL_L_X4Y129_SLICE_X5Y129_AO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B = CLBLL_L_X4Y129_SLICE_X5Y129_BO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C = CLBLL_L_X4Y129_SLICE_X5Y129_CO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D = CLBLL_L_X4Y129_SLICE_X5Y129_DO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_AMUX = CLBLL_L_X4Y129_SLICE_X5Y129_AO5;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_BMUX = CLBLL_L_X4Y129_SLICE_X5Y129_BO5;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A = CLBLL_L_X4Y130_SLICE_X4Y130_AO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B = CLBLL_L_X4Y130_SLICE_X4Y130_BO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C = CLBLL_L_X4Y130_SLICE_X4Y130_CO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D = CLBLL_L_X4Y130_SLICE_X4Y130_DO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_AMUX = CLBLL_L_X4Y130_SLICE_X4Y130_AO5;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A = CLBLL_L_X4Y130_SLICE_X5Y130_AO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B = CLBLL_L_X4Y130_SLICE_X5Y130_BO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C = CLBLL_L_X4Y130_SLICE_X5Y130_CO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D = CLBLL_L_X4Y130_SLICE_X5Y130_DO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_AMUX = CLBLL_L_X4Y130_SLICE_X5Y130_A5Q;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_DMUX = CLBLL_L_X4Y130_SLICE_X5Y130_DO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A = CLBLL_L_X4Y131_SLICE_X4Y131_AO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C = CLBLL_L_X4Y131_SLICE_X4Y131_CO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D = CLBLL_L_X4Y131_SLICE_X4Y131_DO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_AMUX = CLBLL_L_X4Y131_SLICE_X4Y131_AO5;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_BMUX = CLBLL_L_X4Y131_SLICE_X4Y131_BO5;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A = CLBLL_L_X4Y131_SLICE_X5Y131_AO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B = CLBLL_L_X4Y131_SLICE_X5Y131_BO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C = CLBLL_L_X4Y131_SLICE_X5Y131_CO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D = CLBLL_L_X4Y131_SLICE_X5Y131_DO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_AMUX = CLBLL_L_X4Y131_SLICE_X5Y131_AO5;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_BMUX = CLBLL_L_X4Y131_SLICE_X5Y131_B5Q;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A = CLBLL_L_X4Y132_SLICE_X4Y132_AO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B = CLBLL_L_X4Y132_SLICE_X4Y132_BO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C = CLBLL_L_X4Y132_SLICE_X4Y132_CO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D = CLBLL_L_X4Y132_SLICE_X4Y132_DO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_AMUX = CLBLL_L_X4Y132_SLICE_X4Y132_AO5;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_BMUX = CLBLL_L_X4Y132_SLICE_X4Y132_BO5;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_DMUX = CLBLL_L_X4Y132_SLICE_X4Y132_DO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A = CLBLL_L_X4Y132_SLICE_X5Y132_AO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B = CLBLL_L_X4Y132_SLICE_X5Y132_BO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C = CLBLL_L_X4Y132_SLICE_X5Y132_CO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D = CLBLL_L_X4Y132_SLICE_X5Y132_DO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_AMUX = CLBLL_L_X4Y132_SLICE_X5Y132_A5Q;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A = CLBLL_L_X4Y133_SLICE_X4Y133_AO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B = CLBLL_L_X4Y133_SLICE_X4Y133_BO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C = CLBLL_L_X4Y133_SLICE_X4Y133_CO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D = CLBLL_L_X4Y133_SLICE_X4Y133_DO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_AMUX = CLBLL_L_X4Y133_SLICE_X4Y133_A5Q;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_CMUX = CLBLL_L_X4Y133_SLICE_X4Y133_CO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A = CLBLL_L_X4Y133_SLICE_X5Y133_AO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B = CLBLL_L_X4Y133_SLICE_X5Y133_BO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C = CLBLL_L_X4Y133_SLICE_X5Y133_CO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D = CLBLL_L_X4Y133_SLICE_X5Y133_DO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_AMUX = CLBLL_L_X4Y133_SLICE_X5Y133_AO5;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A = CLBLL_L_X4Y134_SLICE_X4Y134_AO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B = CLBLL_L_X4Y134_SLICE_X4Y134_BO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C = CLBLL_L_X4Y134_SLICE_X4Y134_CO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D = CLBLL_L_X4Y134_SLICE_X4Y134_DO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A = CLBLL_L_X4Y134_SLICE_X5Y134_AO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B = CLBLL_L_X4Y134_SLICE_X5Y134_BO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C = CLBLL_L_X4Y134_SLICE_X5Y134_CO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D = CLBLL_L_X4Y134_SLICE_X5Y134_DO6;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_A = CLBLL_L_X4Y135_SLICE_X4Y135_AO6;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_B = CLBLL_L_X4Y135_SLICE_X4Y135_BO6;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_C = CLBLL_L_X4Y135_SLICE_X4Y135_CO6;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_D = CLBLL_L_X4Y135_SLICE_X4Y135_DO6;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_AMUX = CLBLL_L_X4Y135_SLICE_X4Y135_AO5;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_A = CLBLL_L_X4Y135_SLICE_X5Y135_AO6;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_B = CLBLL_L_X4Y135_SLICE_X5Y135_BO6;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_C = CLBLL_L_X4Y135_SLICE_X5Y135_CO6;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_D = CLBLL_L_X4Y135_SLICE_X5Y135_DO6;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_AMUX = CLBLL_L_X4Y135_SLICE_X5Y135_AO5;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_A = CLBLL_L_X4Y136_SLICE_X4Y136_AO6;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_B = CLBLL_L_X4Y136_SLICE_X4Y136_BO6;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_C = CLBLL_L_X4Y136_SLICE_X4Y136_CO6;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_D = CLBLL_L_X4Y136_SLICE_X4Y136_DO6;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_A = CLBLL_L_X4Y136_SLICE_X5Y136_AO6;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_B = CLBLL_L_X4Y136_SLICE_X5Y136_BO6;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_C = CLBLL_L_X4Y136_SLICE_X5Y136_CO6;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_D = CLBLL_L_X4Y136_SLICE_X5Y136_DO6;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_CMUX = CLBLL_L_X4Y136_SLICE_X5Y136_CO6;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_A = CLBLL_L_X4Y137_SLICE_X4Y137_AO6;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_B = CLBLL_L_X4Y137_SLICE_X4Y137_BO6;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_C = CLBLL_L_X4Y137_SLICE_X4Y137_CO6;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_D = CLBLL_L_X4Y137_SLICE_X4Y137_DO6;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_BMUX = CLBLL_L_X4Y137_SLICE_X4Y137_BO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_A = CLBLL_L_X4Y137_SLICE_X5Y137_AO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_B = CLBLL_L_X4Y137_SLICE_X5Y137_BO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_C = CLBLL_L_X4Y137_SLICE_X5Y137_CO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_D = CLBLL_L_X4Y137_SLICE_X5Y137_DO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_AMUX = CLBLL_L_X4Y137_SLICE_X5Y137_AO5;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_BMUX = CLBLL_L_X4Y137_SLICE_X5Y137_BO6;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A = CLBLL_L_X4Y138_SLICE_X4Y138_AO6;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B = CLBLL_L_X4Y138_SLICE_X4Y138_BO6;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C = CLBLL_L_X4Y138_SLICE_X4Y138_CO6;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D = CLBLL_L_X4Y138_SLICE_X4Y138_DO6;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_BMUX = CLBLL_L_X4Y138_SLICE_X4Y138_BO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A = CLBLL_L_X4Y138_SLICE_X5Y138_AO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B = CLBLL_L_X4Y138_SLICE_X5Y138_BO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C = CLBLL_L_X4Y138_SLICE_X5Y138_CO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D = CLBLL_L_X4Y138_SLICE_X5Y138_DO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_A = CLBLL_L_X4Y139_SLICE_X4Y139_AO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_B = CLBLL_L_X4Y139_SLICE_X4Y139_BO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_C = CLBLL_L_X4Y139_SLICE_X4Y139_CO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_D = CLBLL_L_X4Y139_SLICE_X4Y139_DO6;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_A = CLBLL_L_X4Y139_SLICE_X5Y139_AO6;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_B = CLBLL_L_X4Y139_SLICE_X5Y139_BO6;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_C = CLBLL_L_X4Y139_SLICE_X5Y139_CO6;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_D = CLBLL_L_X4Y139_SLICE_X5Y139_DO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A = CLBLL_L_X4Y140_SLICE_X4Y140_AO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B = CLBLL_L_X4Y140_SLICE_X4Y140_BO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C = CLBLL_L_X4Y140_SLICE_X4Y140_CO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D = CLBLL_L_X4Y140_SLICE_X4Y140_DO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B = CLBLL_L_X4Y140_SLICE_X5Y140_BO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C = CLBLL_L_X4Y140_SLICE_X5Y140_CO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D = CLBLL_L_X4Y140_SLICE_X5Y140_DO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_AMUX = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A = CLBLL_L_X4Y145_SLICE_X4Y145_AO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B = CLBLL_L_X4Y145_SLICE_X4Y145_BO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C = CLBLL_L_X4Y145_SLICE_X4Y145_CO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D = CLBLL_L_X4Y145_SLICE_X4Y145_DO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A = CLBLL_L_X4Y145_SLICE_X5Y145_AO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B = CLBLL_L_X4Y145_SLICE_X5Y145_BO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C = CLBLL_L_X4Y145_SLICE_X5Y145_CO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D = CLBLL_L_X4Y145_SLICE_X5Y145_DO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A = CLBLL_L_X4Y146_SLICE_X4Y146_AO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B = CLBLL_L_X4Y146_SLICE_X4Y146_BO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C = CLBLL_L_X4Y146_SLICE_X4Y146_CO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D = CLBLL_L_X4Y146_SLICE_X4Y146_DO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A = CLBLL_L_X4Y146_SLICE_X5Y146_AO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B = CLBLL_L_X4Y146_SLICE_X5Y146_BO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C = CLBLL_L_X4Y146_SLICE_X5Y146_CO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D = CLBLL_L_X4Y146_SLICE_X5Y146_DO6;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_A = CLBLL_L_X4Y155_SLICE_X4Y155_AO6;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_B = CLBLL_L_X4Y155_SLICE_X4Y155_BO6;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_C = CLBLL_L_X4Y155_SLICE_X4Y155_CO6;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_D = CLBLL_L_X4Y155_SLICE_X4Y155_DO6;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_A = CLBLL_L_X4Y155_SLICE_X5Y155_AO6;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_B = CLBLL_L_X4Y155_SLICE_X5Y155_BO6;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_C = CLBLL_L_X4Y155_SLICE_X5Y155_CO6;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_D = CLBLL_L_X4Y155_SLICE_X5Y155_DO6;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_A = CLBLL_L_X4Y156_SLICE_X4Y156_AO6;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_B = CLBLL_L_X4Y156_SLICE_X4Y156_BO6;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_C = CLBLL_L_X4Y156_SLICE_X4Y156_CO6;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_D = CLBLL_L_X4Y156_SLICE_X4Y156_DO6;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_A = CLBLL_L_X4Y156_SLICE_X5Y156_AO6;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_B = CLBLL_L_X4Y156_SLICE_X5Y156_BO6;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_C = CLBLL_L_X4Y156_SLICE_X5Y156_CO6;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_D = CLBLL_L_X4Y156_SLICE_X5Y156_DO6;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_AMUX = CLBLL_L_X4Y156_SLICE_X5Y156_A5Q;
  assign CLBLL_L_X54Y96_SLICE_X82Y96_A = CLBLL_L_X54Y96_SLICE_X82Y96_AO6;
  assign CLBLL_L_X54Y96_SLICE_X82Y96_B = CLBLL_L_X54Y96_SLICE_X82Y96_BO6;
  assign CLBLL_L_X54Y96_SLICE_X82Y96_C = CLBLL_L_X54Y96_SLICE_X82Y96_CO6;
  assign CLBLL_L_X54Y96_SLICE_X82Y96_D = CLBLL_L_X54Y96_SLICE_X82Y96_DO6;
  assign CLBLL_L_X54Y96_SLICE_X83Y96_A = CLBLL_L_X54Y96_SLICE_X83Y96_AO6;
  assign CLBLL_L_X54Y96_SLICE_X83Y96_B = CLBLL_L_X54Y96_SLICE_X83Y96_BO6;
  assign CLBLL_L_X54Y96_SLICE_X83Y96_C = CLBLL_L_X54Y96_SLICE_X83Y96_CO6;
  assign CLBLL_L_X54Y96_SLICE_X83Y96_D = CLBLL_L_X54Y96_SLICE_X83Y96_DO6;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_A = CLBLL_L_X54Y101_SLICE_X82Y101_AO6;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_B = CLBLL_L_X54Y101_SLICE_X82Y101_BO6;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_C = CLBLL_L_X54Y101_SLICE_X82Y101_CO6;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_D = CLBLL_L_X54Y101_SLICE_X82Y101_DO6;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_A = CLBLL_L_X54Y101_SLICE_X83Y101_AO6;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_B = CLBLL_L_X54Y101_SLICE_X83Y101_BO6;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_C = CLBLL_L_X54Y101_SLICE_X83Y101_CO6;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_D = CLBLL_L_X54Y101_SLICE_X83Y101_DO6;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_A = CLBLL_L_X54Y105_SLICE_X82Y105_AO6;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_B = CLBLL_L_X54Y105_SLICE_X82Y105_BO6;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_C = CLBLL_L_X54Y105_SLICE_X82Y105_CO6;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_D = CLBLL_L_X54Y105_SLICE_X82Y105_DO6;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_A = CLBLL_L_X54Y105_SLICE_X83Y105_AO6;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_B = CLBLL_L_X54Y105_SLICE_X83Y105_BO6;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_C = CLBLL_L_X54Y105_SLICE_X83Y105_CO6;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_D = CLBLL_L_X54Y105_SLICE_X83Y105_DO6;
  assign CLBLL_L_X54Y116_SLICE_X82Y116_A = CLBLL_L_X54Y116_SLICE_X82Y116_AO6;
  assign CLBLL_L_X54Y116_SLICE_X82Y116_B = CLBLL_L_X54Y116_SLICE_X82Y116_BO6;
  assign CLBLL_L_X54Y116_SLICE_X82Y116_C = CLBLL_L_X54Y116_SLICE_X82Y116_CO6;
  assign CLBLL_L_X54Y116_SLICE_X82Y116_D = CLBLL_L_X54Y116_SLICE_X82Y116_DO6;
  assign CLBLL_L_X54Y116_SLICE_X83Y116_A = CLBLL_L_X54Y116_SLICE_X83Y116_AO6;
  assign CLBLL_L_X54Y116_SLICE_X83Y116_B = CLBLL_L_X54Y116_SLICE_X83Y116_BO6;
  assign CLBLL_L_X54Y116_SLICE_X83Y116_C = CLBLL_L_X54Y116_SLICE_X83Y116_CO6;
  assign CLBLL_L_X54Y116_SLICE_X83Y116_D = CLBLL_L_X54Y116_SLICE_X83Y116_DO6;
  assign CLBLL_L_X54Y119_SLICE_X82Y119_A = CLBLL_L_X54Y119_SLICE_X82Y119_AO6;
  assign CLBLL_L_X54Y119_SLICE_X82Y119_B = CLBLL_L_X54Y119_SLICE_X82Y119_BO6;
  assign CLBLL_L_X54Y119_SLICE_X82Y119_C = CLBLL_L_X54Y119_SLICE_X82Y119_CO6;
  assign CLBLL_L_X54Y119_SLICE_X82Y119_D = CLBLL_L_X54Y119_SLICE_X82Y119_DO6;
  assign CLBLL_L_X54Y119_SLICE_X83Y119_A = CLBLL_L_X54Y119_SLICE_X83Y119_AO6;
  assign CLBLL_L_X54Y119_SLICE_X83Y119_B = CLBLL_L_X54Y119_SLICE_X83Y119_BO6;
  assign CLBLL_L_X54Y119_SLICE_X83Y119_C = CLBLL_L_X54Y119_SLICE_X83Y119_CO6;
  assign CLBLL_L_X54Y119_SLICE_X83Y119_D = CLBLL_L_X54Y119_SLICE_X83Y119_DO6;
  assign CLBLL_L_X54Y123_SLICE_X82Y123_A = CLBLL_L_X54Y123_SLICE_X82Y123_AO6;
  assign CLBLL_L_X54Y123_SLICE_X82Y123_B = CLBLL_L_X54Y123_SLICE_X82Y123_BO6;
  assign CLBLL_L_X54Y123_SLICE_X82Y123_C = CLBLL_L_X54Y123_SLICE_X82Y123_CO6;
  assign CLBLL_L_X54Y123_SLICE_X82Y123_D = CLBLL_L_X54Y123_SLICE_X82Y123_DO6;
  assign CLBLL_L_X54Y123_SLICE_X83Y123_A = CLBLL_L_X54Y123_SLICE_X83Y123_AO6;
  assign CLBLL_L_X54Y123_SLICE_X83Y123_B = CLBLL_L_X54Y123_SLICE_X83Y123_BO6;
  assign CLBLL_L_X54Y123_SLICE_X83Y123_C = CLBLL_L_X54Y123_SLICE_X83Y123_CO6;
  assign CLBLL_L_X54Y123_SLICE_X83Y123_D = CLBLL_L_X54Y123_SLICE_X83Y123_DO6;
  assign CLBLL_L_X54Y133_SLICE_X82Y133_A = CLBLL_L_X54Y133_SLICE_X82Y133_AO6;
  assign CLBLL_L_X54Y133_SLICE_X82Y133_B = CLBLL_L_X54Y133_SLICE_X82Y133_BO6;
  assign CLBLL_L_X54Y133_SLICE_X82Y133_C = CLBLL_L_X54Y133_SLICE_X82Y133_CO6;
  assign CLBLL_L_X54Y133_SLICE_X82Y133_D = CLBLL_L_X54Y133_SLICE_X82Y133_DO6;
  assign CLBLL_L_X54Y133_SLICE_X83Y133_A = CLBLL_L_X54Y133_SLICE_X83Y133_AO6;
  assign CLBLL_L_X54Y133_SLICE_X83Y133_B = CLBLL_L_X54Y133_SLICE_X83Y133_BO6;
  assign CLBLL_L_X54Y133_SLICE_X83Y133_C = CLBLL_L_X54Y133_SLICE_X83Y133_CO6;
  assign CLBLL_L_X54Y133_SLICE_X83Y133_D = CLBLL_L_X54Y133_SLICE_X83Y133_DO6;
  assign CLBLL_L_X54Y138_SLICE_X82Y138_A = CLBLL_L_X54Y138_SLICE_X82Y138_AO6;
  assign CLBLL_L_X54Y138_SLICE_X82Y138_B = CLBLL_L_X54Y138_SLICE_X82Y138_BO6;
  assign CLBLL_L_X54Y138_SLICE_X82Y138_C = CLBLL_L_X54Y138_SLICE_X82Y138_CO6;
  assign CLBLL_L_X54Y138_SLICE_X82Y138_D = CLBLL_L_X54Y138_SLICE_X82Y138_DO6;
  assign CLBLL_L_X54Y138_SLICE_X83Y138_A = CLBLL_L_X54Y138_SLICE_X83Y138_AO6;
  assign CLBLL_L_X54Y138_SLICE_X83Y138_B = CLBLL_L_X54Y138_SLICE_X83Y138_BO6;
  assign CLBLL_L_X54Y138_SLICE_X83Y138_C = CLBLL_L_X54Y138_SLICE_X83Y138_CO6;
  assign CLBLL_L_X54Y138_SLICE_X83Y138_D = CLBLL_L_X54Y138_SLICE_X83Y138_DO6;
  assign CLBLL_L_X54Y141_SLICE_X82Y141_A = CLBLL_L_X54Y141_SLICE_X82Y141_AO6;
  assign CLBLL_L_X54Y141_SLICE_X82Y141_B = CLBLL_L_X54Y141_SLICE_X82Y141_BO6;
  assign CLBLL_L_X54Y141_SLICE_X82Y141_C = CLBLL_L_X54Y141_SLICE_X82Y141_CO6;
  assign CLBLL_L_X54Y141_SLICE_X82Y141_D = CLBLL_L_X54Y141_SLICE_X82Y141_DO6;
  assign CLBLL_L_X54Y141_SLICE_X83Y141_A = CLBLL_L_X54Y141_SLICE_X83Y141_AO6;
  assign CLBLL_L_X54Y141_SLICE_X83Y141_B = CLBLL_L_X54Y141_SLICE_X83Y141_BO6;
  assign CLBLL_L_X54Y141_SLICE_X83Y141_C = CLBLL_L_X54Y141_SLICE_X83Y141_CO6;
  assign CLBLL_L_X54Y141_SLICE_X83Y141_D = CLBLL_L_X54Y141_SLICE_X83Y141_DO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A = CLBLM_L_X8Y127_SLICE_X10Y127_AO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B = CLBLM_L_X8Y127_SLICE_X10Y127_BO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C = CLBLM_L_X8Y127_SLICE_X10Y127_CO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D = CLBLM_L_X8Y127_SLICE_X10Y127_DO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A = CLBLM_L_X8Y127_SLICE_X11Y127_AO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B = CLBLM_L_X8Y127_SLICE_X11Y127_BO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C = CLBLM_L_X8Y127_SLICE_X11Y127_CO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D = CLBLM_L_X8Y127_SLICE_X11Y127_DO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A = CLBLM_L_X8Y129_SLICE_X10Y129_AO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B = CLBLM_L_X8Y129_SLICE_X10Y129_BO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C = CLBLM_L_X8Y129_SLICE_X10Y129_CO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D = CLBLM_L_X8Y129_SLICE_X10Y129_DO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A = CLBLM_L_X8Y129_SLICE_X11Y129_AO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B = CLBLM_L_X8Y129_SLICE_X11Y129_BO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C = CLBLM_L_X8Y129_SLICE_X11Y129_CO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D = CLBLM_L_X8Y129_SLICE_X11Y129_DO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A = CLBLM_L_X8Y130_SLICE_X10Y130_AO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B = CLBLM_L_X8Y130_SLICE_X10Y130_BO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C = CLBLM_L_X8Y130_SLICE_X10Y130_CO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D = CLBLM_L_X8Y130_SLICE_X10Y130_DO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_AMUX = CLBLM_L_X8Y130_SLICE_X10Y130_A5Q;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_BMUX = CLBLM_L_X8Y130_SLICE_X10Y130_B5Q;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A = CLBLM_L_X8Y130_SLICE_X11Y130_AO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B = CLBLM_L_X8Y130_SLICE_X11Y130_BO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C = CLBLM_L_X8Y130_SLICE_X11Y130_CO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D = CLBLM_L_X8Y130_SLICE_X11Y130_DO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_AMUX = CLBLM_L_X8Y130_SLICE_X11Y130_AO5;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A = CLBLM_L_X8Y131_SLICE_X10Y131_AO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B = CLBLM_L_X8Y131_SLICE_X10Y131_BO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C = CLBLM_L_X8Y131_SLICE_X10Y131_CO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D = CLBLM_L_X8Y131_SLICE_X10Y131_DO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A = CLBLM_L_X8Y131_SLICE_X11Y131_AO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B = CLBLM_L_X8Y131_SLICE_X11Y131_BO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C = CLBLM_L_X8Y131_SLICE_X11Y131_CO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D = CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A = CLBLM_L_X8Y132_SLICE_X10Y132_AO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B = CLBLM_L_X8Y132_SLICE_X10Y132_BO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C = CLBLM_L_X8Y132_SLICE_X10Y132_CO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D = CLBLM_L_X8Y132_SLICE_X10Y132_DO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A = CLBLM_L_X8Y132_SLICE_X11Y132_AO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B = CLBLM_L_X8Y132_SLICE_X11Y132_BO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C = CLBLM_L_X8Y132_SLICE_X11Y132_CO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D = CLBLM_L_X8Y132_SLICE_X11Y132_DO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_AMUX = CLBLM_L_X8Y132_SLICE_X11Y132_A5Q;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A = CLBLM_L_X8Y133_SLICE_X10Y133_AO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B = CLBLM_L_X8Y133_SLICE_X10Y133_BO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C = CLBLM_L_X8Y133_SLICE_X10Y133_CO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D = CLBLM_L_X8Y133_SLICE_X10Y133_DO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A = CLBLM_L_X8Y133_SLICE_X11Y133_AO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B = CLBLM_L_X8Y133_SLICE_X11Y133_BO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C = CLBLM_L_X8Y133_SLICE_X11Y133_CO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D = CLBLM_L_X8Y133_SLICE_X11Y133_DO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_AMUX = CLBLM_L_X8Y133_SLICE_X11Y133_AO5;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A = CLBLM_L_X8Y134_SLICE_X10Y134_AO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B = CLBLM_L_X8Y134_SLICE_X10Y134_BO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C = CLBLM_L_X8Y134_SLICE_X10Y134_CO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D = CLBLM_L_X8Y134_SLICE_X10Y134_DO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A = CLBLM_L_X8Y134_SLICE_X11Y134_AO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B = CLBLM_L_X8Y134_SLICE_X11Y134_BO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C = CLBLM_L_X8Y134_SLICE_X11Y134_CO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D = CLBLM_L_X8Y134_SLICE_X11Y134_DO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A = CLBLM_L_X8Y135_SLICE_X10Y135_AO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B = CLBLM_L_X8Y135_SLICE_X10Y135_BO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C = CLBLM_L_X8Y135_SLICE_X10Y135_CO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D = CLBLM_L_X8Y135_SLICE_X10Y135_DO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_AMUX = CLBLM_L_X8Y135_SLICE_X10Y135_A5Q;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_BMUX = CLBLM_L_X8Y135_SLICE_X10Y135_BO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_CMUX = CLBLM_L_X8Y135_SLICE_X10Y135_CO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A = CLBLM_L_X8Y135_SLICE_X11Y135_AO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B = CLBLM_L_X8Y135_SLICE_X11Y135_BO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C = CLBLM_L_X8Y135_SLICE_X11Y135_CO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D = CLBLM_L_X8Y135_SLICE_X11Y135_DO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A = CLBLM_L_X8Y136_SLICE_X10Y136_AO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B = CLBLM_L_X8Y136_SLICE_X10Y136_BO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C = CLBLM_L_X8Y136_SLICE_X10Y136_CO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D = CLBLM_L_X8Y136_SLICE_X10Y136_DO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_AMUX = CLBLM_L_X8Y136_SLICE_X10Y136_A5Q;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_BMUX = CLBLM_L_X8Y136_SLICE_X10Y136_BO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A = CLBLM_L_X8Y136_SLICE_X11Y136_AO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B = CLBLM_L_X8Y136_SLICE_X11Y136_BO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C = CLBLM_L_X8Y136_SLICE_X11Y136_CO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D = CLBLM_L_X8Y136_SLICE_X11Y136_DO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_A = CLBLM_L_X8Y137_SLICE_X10Y137_AO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_B = CLBLM_L_X8Y137_SLICE_X10Y137_BO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_C = CLBLM_L_X8Y137_SLICE_X10Y137_CO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_D = CLBLM_L_X8Y137_SLICE_X10Y137_DO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_AMUX = CLBLM_L_X8Y137_SLICE_X10Y137_A5Q;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_BMUX = CLBLM_L_X8Y137_SLICE_X10Y137_B5Q;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_A = CLBLM_L_X8Y137_SLICE_X11Y137_AO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_B = CLBLM_L_X8Y137_SLICE_X11Y137_BO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_C = CLBLM_L_X8Y137_SLICE_X11Y137_CO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_D = CLBLM_L_X8Y137_SLICE_X11Y137_DO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_A = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_B = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_C = CLBLM_L_X8Y138_SLICE_X10Y138_CO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_D = CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_A = CLBLM_L_X8Y138_SLICE_X11Y138_AO6;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_B = CLBLM_L_X8Y138_SLICE_X11Y138_BO6;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_C = CLBLM_L_X8Y138_SLICE_X11Y138_CO6;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_D = CLBLM_L_X8Y138_SLICE_X11Y138_DO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A = CLBLM_L_X10Y130_SLICE_X12Y130_AO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B = CLBLM_L_X10Y130_SLICE_X12Y130_BO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C = CLBLM_L_X10Y130_SLICE_X12Y130_CO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D = CLBLM_L_X10Y130_SLICE_X12Y130_DO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A = CLBLM_L_X10Y130_SLICE_X13Y130_AO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B = CLBLM_L_X10Y130_SLICE_X13Y130_BO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C = CLBLM_L_X10Y130_SLICE_X13Y130_CO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D = CLBLM_L_X10Y130_SLICE_X13Y130_DO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A = CLBLM_L_X10Y131_SLICE_X12Y131_AO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B = CLBLM_L_X10Y131_SLICE_X12Y131_BO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C = CLBLM_L_X10Y131_SLICE_X12Y131_CO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D = CLBLM_L_X10Y131_SLICE_X12Y131_DO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A = CLBLM_L_X10Y131_SLICE_X13Y131_AO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B = CLBLM_L_X10Y131_SLICE_X13Y131_BO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C = CLBLM_L_X10Y131_SLICE_X13Y131_CO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D = CLBLM_L_X10Y131_SLICE_X13Y131_DO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A = CLBLM_L_X10Y132_SLICE_X12Y132_AO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B = CLBLM_L_X10Y132_SLICE_X12Y132_BO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C = CLBLM_L_X10Y132_SLICE_X12Y132_CO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D = CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A = CLBLM_L_X10Y132_SLICE_X13Y132_AO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B = CLBLM_L_X10Y132_SLICE_X13Y132_BO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C = CLBLM_L_X10Y132_SLICE_X13Y132_CO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D = CLBLM_L_X10Y132_SLICE_X13Y132_DO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A = CLBLM_L_X10Y133_SLICE_X12Y133_AO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B = CLBLM_L_X10Y133_SLICE_X12Y133_BO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C = CLBLM_L_X10Y133_SLICE_X12Y133_CO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D = CLBLM_L_X10Y133_SLICE_X12Y133_DO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A = CLBLM_L_X10Y133_SLICE_X13Y133_AO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B = CLBLM_L_X10Y133_SLICE_X13Y133_BO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C = CLBLM_L_X10Y133_SLICE_X13Y133_CO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A = CLBLM_L_X10Y134_SLICE_X12Y134_AO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B = CLBLM_L_X10Y134_SLICE_X12Y134_BO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C = CLBLM_L_X10Y134_SLICE_X12Y134_CO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D = CLBLM_L_X10Y134_SLICE_X12Y134_DO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A = CLBLM_L_X10Y134_SLICE_X13Y134_AO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B = CLBLM_L_X10Y134_SLICE_X13Y134_BO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C = CLBLM_L_X10Y134_SLICE_X13Y134_CO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D = CLBLM_L_X10Y134_SLICE_X13Y134_DO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A = CLBLM_L_X10Y135_SLICE_X12Y135_AO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B = CLBLM_L_X10Y135_SLICE_X12Y135_BO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C = CLBLM_L_X10Y135_SLICE_X12Y135_CO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D = CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_AMUX = CLBLM_L_X10Y135_SLICE_X12Y135_A5Q;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A = CLBLM_L_X10Y135_SLICE_X13Y135_AO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B = CLBLM_L_X10Y135_SLICE_X13Y135_BO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C = CLBLM_L_X10Y135_SLICE_X13Y135_CO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D = CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A = CLBLM_L_X10Y136_SLICE_X12Y136_AO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B = CLBLM_L_X10Y136_SLICE_X12Y136_BO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C = CLBLM_L_X10Y136_SLICE_X12Y136_CO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D = CLBLM_L_X10Y136_SLICE_X12Y136_DO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A = CLBLM_L_X10Y136_SLICE_X13Y136_AO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B = CLBLM_L_X10Y136_SLICE_X13Y136_BO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C = CLBLM_L_X10Y136_SLICE_X13Y136_CO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D = CLBLM_L_X10Y136_SLICE_X13Y136_DO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_AMUX = CLBLM_L_X10Y136_SLICE_X13Y136_AO5;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_BMUX = CLBLM_L_X10Y136_SLICE_X13Y136_BO5;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A = CLBLM_L_X10Y137_SLICE_X12Y137_AO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B = CLBLM_L_X10Y137_SLICE_X12Y137_BO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C = CLBLM_L_X10Y137_SLICE_X12Y137_CO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D = CLBLM_L_X10Y137_SLICE_X12Y137_DO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_AMUX = CLBLM_L_X10Y137_SLICE_X12Y137_AO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A = CLBLM_L_X10Y137_SLICE_X13Y137_AO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B = CLBLM_L_X10Y137_SLICE_X13Y137_BO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C = CLBLM_L_X10Y137_SLICE_X13Y137_CO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D = CLBLM_L_X10Y137_SLICE_X13Y137_DO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A = CLBLM_L_X10Y138_SLICE_X12Y138_AO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B = CLBLM_L_X10Y138_SLICE_X12Y138_BO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C = CLBLM_L_X10Y138_SLICE_X12Y138_CO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D = CLBLM_L_X10Y138_SLICE_X12Y138_DO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A = CLBLM_L_X10Y138_SLICE_X13Y138_AO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B = CLBLM_L_X10Y138_SLICE_X13Y138_BO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C = CLBLM_L_X10Y138_SLICE_X13Y138_CO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D = CLBLM_L_X10Y138_SLICE_X13Y138_DO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A = CLBLM_L_X12Y130_SLICE_X16Y130_AO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B = CLBLM_L_X12Y130_SLICE_X16Y130_BO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C = CLBLM_L_X12Y130_SLICE_X16Y130_CO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D = CLBLM_L_X12Y130_SLICE_X16Y130_DO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A = CLBLM_L_X12Y130_SLICE_X17Y130_AO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B = CLBLM_L_X12Y130_SLICE_X17Y130_BO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C = CLBLM_L_X12Y130_SLICE_X17Y130_CO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D = CLBLM_L_X12Y130_SLICE_X17Y130_DO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A = CLBLM_L_X12Y132_SLICE_X16Y132_AO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B = CLBLM_L_X12Y132_SLICE_X16Y132_BO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C = CLBLM_L_X12Y132_SLICE_X16Y132_CO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D = CLBLM_L_X12Y132_SLICE_X16Y132_DO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A = CLBLM_L_X12Y132_SLICE_X17Y132_AO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B = CLBLM_L_X12Y132_SLICE_X17Y132_BO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C = CLBLM_L_X12Y132_SLICE_X17Y132_CO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D = CLBLM_L_X12Y132_SLICE_X17Y132_DO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A = CLBLM_L_X12Y135_SLICE_X16Y135_AO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B = CLBLM_L_X12Y135_SLICE_X16Y135_BO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C = CLBLM_L_X12Y135_SLICE_X16Y135_CO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D = CLBLM_L_X12Y135_SLICE_X16Y135_DO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A = CLBLM_L_X12Y135_SLICE_X17Y135_AO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B = CLBLM_L_X12Y135_SLICE_X17Y135_BO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C = CLBLM_L_X12Y135_SLICE_X17Y135_CO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D = CLBLM_L_X12Y135_SLICE_X17Y135_DO6;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_A = CLBLM_L_X16Y135_SLICE_X22Y135_AO6;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_B = CLBLM_L_X16Y135_SLICE_X22Y135_BO6;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_C = CLBLM_L_X16Y135_SLICE_X22Y135_CO6;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_D = CLBLM_L_X16Y135_SLICE_X22Y135_DO6;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_A = CLBLM_L_X16Y135_SLICE_X23Y135_AO6;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_B = CLBLM_L_X16Y135_SLICE_X23Y135_BO6;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_C = CLBLM_L_X16Y135_SLICE_X23Y135_CO6;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_D = CLBLM_L_X16Y135_SLICE_X23Y135_DO6;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_A = CLBLM_L_X16Y136_SLICE_X22Y136_AO6;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_B = CLBLM_L_X16Y136_SLICE_X22Y136_BO6;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_C = CLBLM_L_X16Y136_SLICE_X22Y136_CO6;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_D = CLBLM_L_X16Y136_SLICE_X22Y136_DO6;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_A = CLBLM_L_X16Y136_SLICE_X23Y136_AO6;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_B = CLBLM_L_X16Y136_SLICE_X23Y136_BO6;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_C = CLBLM_L_X16Y136_SLICE_X23Y136_CO6;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_D = CLBLM_L_X16Y136_SLICE_X23Y136_DO6;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_A = CLBLM_L_X16Y137_SLICE_X22Y137_AO6;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_B = CLBLM_L_X16Y137_SLICE_X22Y137_BO6;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_C = CLBLM_L_X16Y137_SLICE_X22Y137_CO6;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_D = CLBLM_L_X16Y137_SLICE_X22Y137_DO6;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_A = CLBLM_L_X16Y137_SLICE_X23Y137_AO6;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_B = CLBLM_L_X16Y137_SLICE_X23Y137_BO6;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_C = CLBLM_L_X16Y137_SLICE_X23Y137_CO6;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_D = CLBLM_L_X16Y137_SLICE_X23Y137_DO6;
  assign CLBLM_L_X16Y149_SLICE_X22Y149_A = CLBLM_L_X16Y149_SLICE_X22Y149_AO6;
  assign CLBLM_L_X16Y149_SLICE_X22Y149_B = CLBLM_L_X16Y149_SLICE_X22Y149_BO6;
  assign CLBLM_L_X16Y149_SLICE_X22Y149_C = CLBLM_L_X16Y149_SLICE_X22Y149_CO6;
  assign CLBLM_L_X16Y149_SLICE_X22Y149_D = CLBLM_L_X16Y149_SLICE_X22Y149_DO6;
  assign CLBLM_L_X16Y149_SLICE_X23Y149_A = CLBLM_L_X16Y149_SLICE_X23Y149_AO6;
  assign CLBLM_L_X16Y149_SLICE_X23Y149_B = CLBLM_L_X16Y149_SLICE_X23Y149_BO6;
  assign CLBLM_L_X16Y149_SLICE_X23Y149_C = CLBLM_L_X16Y149_SLICE_X23Y149_CO6;
  assign CLBLM_L_X16Y149_SLICE_X23Y149_D = CLBLM_L_X16Y149_SLICE_X23Y149_DO6;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_A = CLBLM_L_X16Y151_SLICE_X22Y151_AO6;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_B = CLBLM_L_X16Y151_SLICE_X22Y151_BO6;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_C = CLBLM_L_X16Y151_SLICE_X22Y151_CO6;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_D = CLBLM_L_X16Y151_SLICE_X22Y151_DO6;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_A = CLBLM_L_X16Y151_SLICE_X23Y151_AO6;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_B = CLBLM_L_X16Y151_SLICE_X23Y151_BO6;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_C = CLBLM_L_X16Y151_SLICE_X23Y151_CO6;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_D = CLBLM_L_X16Y151_SLICE_X23Y151_DO6;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_A = CLBLM_L_X16Y152_SLICE_X22Y152_AO6;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_B = CLBLM_L_X16Y152_SLICE_X22Y152_BO6;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_C = CLBLM_L_X16Y152_SLICE_X22Y152_CO6;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_D = CLBLM_L_X16Y152_SLICE_X22Y152_DO6;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_A = CLBLM_L_X16Y152_SLICE_X23Y152_AO6;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_B = CLBLM_L_X16Y152_SLICE_X23Y152_BO6;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_C = CLBLM_L_X16Y152_SLICE_X23Y152_CO6;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_D = CLBLM_L_X16Y152_SLICE_X23Y152_DO6;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_A = CLBLM_L_X16Y153_SLICE_X22Y153_AO6;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_B = CLBLM_L_X16Y153_SLICE_X22Y153_BO6;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_C = CLBLM_L_X16Y153_SLICE_X22Y153_CO6;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_D = CLBLM_L_X16Y153_SLICE_X22Y153_DO6;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_A = CLBLM_L_X16Y153_SLICE_X23Y153_AO6;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_B = CLBLM_L_X16Y153_SLICE_X23Y153_BO6;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_C = CLBLM_L_X16Y153_SLICE_X23Y153_CO6;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_D = CLBLM_L_X16Y153_SLICE_X23Y153_DO6;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_A = CLBLM_L_X16Y154_SLICE_X22Y154_AO6;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_B = CLBLM_L_X16Y154_SLICE_X22Y154_BO6;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_C = CLBLM_L_X16Y154_SLICE_X22Y154_CO6;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_D = CLBLM_L_X16Y154_SLICE_X22Y154_DO6;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_A = CLBLM_L_X16Y154_SLICE_X23Y154_AO6;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_B = CLBLM_L_X16Y154_SLICE_X23Y154_BO6;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_C = CLBLM_L_X16Y154_SLICE_X23Y154_CO6;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_D = CLBLM_L_X16Y154_SLICE_X23Y154_DO6;
  assign CLBLM_L_X16Y155_SLICE_X22Y155_A = CLBLM_L_X16Y155_SLICE_X22Y155_AO6;
  assign CLBLM_L_X16Y155_SLICE_X22Y155_B = CLBLM_L_X16Y155_SLICE_X22Y155_BO6;
  assign CLBLM_L_X16Y155_SLICE_X22Y155_C = CLBLM_L_X16Y155_SLICE_X22Y155_CO6;
  assign CLBLM_L_X16Y155_SLICE_X22Y155_D = CLBLM_L_X16Y155_SLICE_X22Y155_DO6;
  assign CLBLM_L_X16Y155_SLICE_X23Y155_A = CLBLM_L_X16Y155_SLICE_X23Y155_AO6;
  assign CLBLM_L_X16Y155_SLICE_X23Y155_B = CLBLM_L_X16Y155_SLICE_X23Y155_BO6;
  assign CLBLM_L_X16Y155_SLICE_X23Y155_C = CLBLM_L_X16Y155_SLICE_X23Y155_CO6;
  assign CLBLM_L_X16Y155_SLICE_X23Y155_D = CLBLM_L_X16Y155_SLICE_X23Y155_DO6;
  assign CLBLM_L_X16Y157_SLICE_X22Y157_A = CLBLM_L_X16Y157_SLICE_X22Y157_AO6;
  assign CLBLM_L_X16Y157_SLICE_X22Y157_B = CLBLM_L_X16Y157_SLICE_X22Y157_BO6;
  assign CLBLM_L_X16Y157_SLICE_X22Y157_C = CLBLM_L_X16Y157_SLICE_X22Y157_CO6;
  assign CLBLM_L_X16Y157_SLICE_X22Y157_D = CLBLM_L_X16Y157_SLICE_X22Y157_DO6;
  assign CLBLM_L_X16Y157_SLICE_X23Y157_A = CLBLM_L_X16Y157_SLICE_X23Y157_AO6;
  assign CLBLM_L_X16Y157_SLICE_X23Y157_B = CLBLM_L_X16Y157_SLICE_X23Y157_BO6;
  assign CLBLM_L_X16Y157_SLICE_X23Y157_C = CLBLM_L_X16Y157_SLICE_X23Y157_CO6;
  assign CLBLM_L_X16Y157_SLICE_X23Y157_D = CLBLM_L_X16Y157_SLICE_X23Y157_DO6;
  assign CLBLM_L_X56Y151_SLICE_X84Y151_A = CLBLM_L_X56Y151_SLICE_X84Y151_AO6;
  assign CLBLM_L_X56Y151_SLICE_X84Y151_B = CLBLM_L_X56Y151_SLICE_X84Y151_BO6;
  assign CLBLM_L_X56Y151_SLICE_X84Y151_C = CLBLM_L_X56Y151_SLICE_X84Y151_CO6;
  assign CLBLM_L_X56Y151_SLICE_X84Y151_D = CLBLM_L_X56Y151_SLICE_X84Y151_DO6;
  assign CLBLM_L_X56Y151_SLICE_X85Y151_A = CLBLM_L_X56Y151_SLICE_X85Y151_AO6;
  assign CLBLM_L_X56Y151_SLICE_X85Y151_B = CLBLM_L_X56Y151_SLICE_X85Y151_BO6;
  assign CLBLM_L_X56Y151_SLICE_X85Y151_C = CLBLM_L_X56Y151_SLICE_X85Y151_CO6;
  assign CLBLM_L_X56Y151_SLICE_X85Y151_D = CLBLM_L_X56Y151_SLICE_X85Y151_DO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A = CLBLM_R_X3Y129_SLICE_X2Y129_AO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B = CLBLM_R_X3Y129_SLICE_X2Y129_BO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C = CLBLM_R_X3Y129_SLICE_X2Y129_CO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D = CLBLM_R_X3Y129_SLICE_X2Y129_DO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_AMUX = CLBLM_R_X3Y129_SLICE_X2Y129_A5Q;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A = CLBLM_R_X3Y129_SLICE_X3Y129_AO6;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B = CLBLM_R_X3Y129_SLICE_X3Y129_BO6;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C = CLBLM_R_X3Y129_SLICE_X3Y129_CO6;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D = CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A = CLBLM_R_X3Y130_SLICE_X2Y130_AO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B = CLBLM_R_X3Y130_SLICE_X2Y130_BO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C = CLBLM_R_X3Y130_SLICE_X2Y130_CO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D = CLBLM_R_X3Y130_SLICE_X2Y130_DO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A = CLBLM_R_X3Y130_SLICE_X3Y130_AO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B = CLBLM_R_X3Y130_SLICE_X3Y130_BO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C = CLBLM_R_X3Y130_SLICE_X3Y130_CO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D = CLBLM_R_X3Y130_SLICE_X3Y130_DO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_AMUX = CLBLM_R_X3Y130_SLICE_X3Y130_AO5;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A = CLBLM_R_X3Y131_SLICE_X2Y131_AO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B = CLBLM_R_X3Y131_SLICE_X2Y131_BO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C = CLBLM_R_X3Y131_SLICE_X2Y131_CO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D = CLBLM_R_X3Y131_SLICE_X2Y131_DO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_AMUX = CLBLM_R_X3Y131_SLICE_X2Y131_A5Q;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_BMUX = CLBLM_R_X3Y131_SLICE_X2Y131_B5Q;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_CMUX = CLBLM_R_X3Y131_SLICE_X2Y131_C5Q;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_DMUX = CLBLM_R_X3Y131_SLICE_X2Y131_DO5;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A = CLBLM_R_X3Y131_SLICE_X3Y131_AO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B = CLBLM_R_X3Y131_SLICE_X3Y131_BO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C = CLBLM_R_X3Y131_SLICE_X3Y131_CO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D = CLBLM_R_X3Y131_SLICE_X3Y131_DO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_AMUX = CLBLM_R_X3Y131_SLICE_X3Y131_AO5;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_BMUX = CLBLM_R_X3Y131_SLICE_X3Y131_B5Q;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A = CLBLM_R_X3Y132_SLICE_X2Y132_AO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B = CLBLM_R_X3Y132_SLICE_X2Y132_BO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C = CLBLM_R_X3Y132_SLICE_X2Y132_CO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D = CLBLM_R_X3Y132_SLICE_X2Y132_DO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_AMUX = CLBLM_R_X3Y132_SLICE_X2Y132_AO5;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_BMUX = CLBLM_R_X3Y132_SLICE_X2Y132_BO5;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A = CLBLM_R_X3Y132_SLICE_X3Y132_AO6;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B = CLBLM_R_X3Y132_SLICE_X3Y132_BO6;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C = CLBLM_R_X3Y132_SLICE_X3Y132_CO6;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D = CLBLM_R_X3Y132_SLICE_X3Y132_DO6;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_AMUX = CLBLM_R_X3Y132_SLICE_X3Y132_AO5;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A = CLBLM_R_X3Y133_SLICE_X2Y133_AO6;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B = CLBLM_R_X3Y133_SLICE_X2Y133_BO6;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C = CLBLM_R_X3Y133_SLICE_X2Y133_CO6;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D = CLBLM_R_X3Y133_SLICE_X2Y133_DO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A = CLBLM_R_X3Y133_SLICE_X3Y133_AO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B = CLBLM_R_X3Y133_SLICE_X3Y133_BO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C = CLBLM_R_X3Y133_SLICE_X3Y133_CO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D = CLBLM_R_X3Y133_SLICE_X3Y133_DO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_AMUX = CLBLM_R_X3Y133_SLICE_X3Y133_AO5;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_A = CLBLM_R_X3Y134_SLICE_X2Y134_AO6;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_B = CLBLM_R_X3Y134_SLICE_X2Y134_BO6;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_C = CLBLM_R_X3Y134_SLICE_X2Y134_CO6;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_D = CLBLM_R_X3Y134_SLICE_X2Y134_DO6;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_AMUX = CLBLM_R_X3Y134_SLICE_X2Y134_AO5;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_A = CLBLM_R_X3Y134_SLICE_X3Y134_AO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_B = CLBLM_R_X3Y134_SLICE_X3Y134_BO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_C = CLBLM_R_X3Y134_SLICE_X3Y134_CO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_D = CLBLM_R_X3Y134_SLICE_X3Y134_DO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_AMUX = CLBLM_R_X3Y134_SLICE_X3Y134_AO6;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_A = CLBLM_R_X3Y135_SLICE_X2Y135_AO6;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_B = CLBLM_R_X3Y135_SLICE_X2Y135_BO6;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_C = CLBLM_R_X3Y135_SLICE_X2Y135_CO6;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_D = CLBLM_R_X3Y135_SLICE_X2Y135_DO6;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_A = CLBLM_R_X3Y135_SLICE_X3Y135_AO6;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_B = CLBLM_R_X3Y135_SLICE_X3Y135_BO6;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_C = CLBLM_R_X3Y135_SLICE_X3Y135_CO6;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_D = CLBLM_R_X3Y135_SLICE_X3Y135_DO6;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_AMUX = CLBLM_R_X3Y135_SLICE_X3Y135_AO6;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_BMUX = CLBLM_R_X3Y135_SLICE_X3Y135_BO6;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_A = CLBLM_R_X3Y137_SLICE_X2Y137_AO6;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_B = CLBLM_R_X3Y137_SLICE_X2Y137_BO6;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_C = CLBLM_R_X3Y137_SLICE_X2Y137_CO6;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_D = CLBLM_R_X3Y137_SLICE_X2Y137_DO6;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_A = CLBLM_R_X3Y137_SLICE_X3Y137_AO6;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_B = CLBLM_R_X3Y137_SLICE_X3Y137_BO6;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_C = CLBLM_R_X3Y137_SLICE_X3Y137_CO6;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_D = CLBLM_R_X3Y137_SLICE_X3Y137_DO6;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_AMUX = CLBLM_R_X3Y137_SLICE_X3Y137_AO5;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_A = CLBLM_R_X3Y138_SLICE_X2Y138_AO6;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_B = CLBLM_R_X3Y138_SLICE_X2Y138_BO6;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_C = CLBLM_R_X3Y138_SLICE_X2Y138_CO6;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_D = CLBLM_R_X3Y138_SLICE_X2Y138_DO6;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_A = CLBLM_R_X3Y138_SLICE_X3Y138_AO6;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_B = CLBLM_R_X3Y138_SLICE_X3Y138_BO6;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_C = CLBLM_R_X3Y138_SLICE_X3Y138_CO6;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_D = CLBLM_R_X3Y138_SLICE_X3Y138_DO6;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_A = CLBLM_R_X3Y139_SLICE_X2Y139_AO6;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_B = CLBLM_R_X3Y139_SLICE_X2Y139_BO6;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_C = CLBLM_R_X3Y139_SLICE_X2Y139_CO6;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_D = CLBLM_R_X3Y139_SLICE_X2Y139_DO6;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_A = CLBLM_R_X3Y139_SLICE_X3Y139_AO6;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_B = CLBLM_R_X3Y139_SLICE_X3Y139_BO6;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_C = CLBLM_R_X3Y139_SLICE_X3Y139_CO6;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_D = CLBLM_R_X3Y139_SLICE_X3Y139_DO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A = CLBLM_R_X3Y141_SLICE_X2Y141_AO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B = CLBLM_R_X3Y141_SLICE_X2Y141_BO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C = CLBLM_R_X3Y141_SLICE_X2Y141_CO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D = CLBLM_R_X3Y141_SLICE_X2Y141_DO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A = CLBLM_R_X3Y141_SLICE_X3Y141_AO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B = CLBLM_R_X3Y141_SLICE_X3Y141_BO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C = CLBLM_R_X3Y141_SLICE_X3Y141_CO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D = CLBLM_R_X3Y141_SLICE_X3Y141_DO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A = CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B = CLBLM_R_X3Y142_SLICE_X2Y142_BO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C = CLBLM_R_X3Y142_SLICE_X2Y142_CO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D = CLBLM_R_X3Y142_SLICE_X2Y142_DO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A = CLBLM_R_X3Y142_SLICE_X3Y142_AO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B = CLBLM_R_X3Y142_SLICE_X3Y142_BO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C = CLBLM_R_X3Y142_SLICE_X3Y142_CO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D = CLBLM_R_X3Y142_SLICE_X3Y142_DO6;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A = CLBLM_R_X3Y145_SLICE_X2Y145_AO6;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B = CLBLM_R_X3Y145_SLICE_X2Y145_BO6;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C = CLBLM_R_X3Y145_SLICE_X2Y145_CO6;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D = CLBLM_R_X3Y145_SLICE_X2Y145_DO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A = CLBLM_R_X3Y145_SLICE_X3Y145_AO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B = CLBLM_R_X3Y145_SLICE_X3Y145_BO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C = CLBLM_R_X3Y145_SLICE_X3Y145_CO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D = CLBLM_R_X3Y145_SLICE_X3Y145_DO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A = CLBLM_R_X3Y147_SLICE_X2Y147_AO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B = CLBLM_R_X3Y147_SLICE_X2Y147_BO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C = CLBLM_R_X3Y147_SLICE_X2Y147_CO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D = CLBLM_R_X3Y147_SLICE_X2Y147_DO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A = CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B = CLBLM_R_X3Y147_SLICE_X3Y147_BO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C = CLBLM_R_X3Y147_SLICE_X3Y147_CO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D = CLBLM_R_X3Y147_SLICE_X3Y147_DO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A = CLBLM_R_X3Y149_SLICE_X2Y149_AO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B = CLBLM_R_X3Y149_SLICE_X2Y149_BO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C = CLBLM_R_X3Y149_SLICE_X2Y149_CO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D = CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A = CLBLM_R_X3Y149_SLICE_X3Y149_AO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B = CLBLM_R_X3Y149_SLICE_X3Y149_BO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C = CLBLM_R_X3Y149_SLICE_X3Y149_CO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A = CLBLM_R_X3Y151_SLICE_X2Y151_AO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B = CLBLM_R_X3Y151_SLICE_X2Y151_BO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C = CLBLM_R_X3Y151_SLICE_X2Y151_CO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D = CLBLM_R_X3Y151_SLICE_X2Y151_DO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A = CLBLM_R_X3Y151_SLICE_X3Y151_AO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B = CLBLM_R_X3Y151_SLICE_X3Y151_BO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C = CLBLM_R_X3Y151_SLICE_X3Y151_CO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D = CLBLM_R_X3Y151_SLICE_X3Y151_DO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A = CLBLM_R_X3Y153_SLICE_X2Y153_AO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B = CLBLM_R_X3Y153_SLICE_X2Y153_BO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C = CLBLM_R_X3Y153_SLICE_X2Y153_CO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D = CLBLM_R_X3Y153_SLICE_X2Y153_DO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A = CLBLM_R_X3Y153_SLICE_X3Y153_AO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B = CLBLM_R_X3Y153_SLICE_X3Y153_BO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C = CLBLM_R_X3Y153_SLICE_X3Y153_CO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D = CLBLM_R_X3Y153_SLICE_X3Y153_DO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_A = CLBLM_R_X3Y155_SLICE_X2Y155_AO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_B = CLBLM_R_X3Y155_SLICE_X2Y155_BO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_C = CLBLM_R_X3Y155_SLICE_X2Y155_CO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_D = CLBLM_R_X3Y155_SLICE_X2Y155_DO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_A = CLBLM_R_X3Y155_SLICE_X3Y155_AO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_B = CLBLM_R_X3Y155_SLICE_X3Y155_BO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_C = CLBLM_R_X3Y155_SLICE_X3Y155_CO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_D = CLBLM_R_X3Y155_SLICE_X3Y155_DO6;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_A = CLBLM_R_X3Y157_SLICE_X2Y157_AO6;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_B = CLBLM_R_X3Y157_SLICE_X2Y157_BO6;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_C = CLBLM_R_X3Y157_SLICE_X2Y157_CO6;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_D = CLBLM_R_X3Y157_SLICE_X2Y157_DO6;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_A = CLBLM_R_X3Y157_SLICE_X3Y157_AO6;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_B = CLBLM_R_X3Y157_SLICE_X3Y157_BO6;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_C = CLBLM_R_X3Y157_SLICE_X3Y157_CO6;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_D = CLBLM_R_X3Y157_SLICE_X3Y157_DO6;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_A = CLBLM_R_X3Y158_SLICE_X2Y158_AO6;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_B = CLBLM_R_X3Y158_SLICE_X2Y158_BO6;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_C = CLBLM_R_X3Y158_SLICE_X2Y158_CO6;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_D = CLBLM_R_X3Y158_SLICE_X2Y158_DO6;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_A = CLBLM_R_X3Y158_SLICE_X3Y158_AO6;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_B = CLBLM_R_X3Y158_SLICE_X3Y158_BO6;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_C = CLBLM_R_X3Y158_SLICE_X3Y158_CO6;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_D = CLBLM_R_X3Y158_SLICE_X3Y158_DO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A = CLBLM_R_X5Y125_SLICE_X6Y125_AO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B = CLBLM_R_X5Y125_SLICE_X6Y125_BO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C = CLBLM_R_X5Y125_SLICE_X6Y125_CO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D = CLBLM_R_X5Y125_SLICE_X6Y125_DO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A = CLBLM_R_X5Y125_SLICE_X7Y125_AO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B = CLBLM_R_X5Y125_SLICE_X7Y125_BO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C = CLBLM_R_X5Y125_SLICE_X7Y125_CO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D = CLBLM_R_X5Y125_SLICE_X7Y125_DO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_AMUX = CLBLM_R_X5Y125_SLICE_X7Y125_AO5;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_BMUX = CLBLM_R_X5Y125_SLICE_X7Y125_BO5;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A = CLBLM_R_X5Y126_SLICE_X6Y126_AO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B = CLBLM_R_X5Y126_SLICE_X6Y126_BO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C = CLBLM_R_X5Y126_SLICE_X6Y126_CO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D = CLBLM_R_X5Y126_SLICE_X6Y126_DO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_AMUX = CLBLM_R_X5Y126_SLICE_X6Y126_AO5;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_CMUX = CLBLM_R_X5Y126_SLICE_X6Y126_CO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A = CLBLM_R_X5Y126_SLICE_X7Y126_AO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B = CLBLM_R_X5Y126_SLICE_X7Y126_BO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C = CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D = CLBLM_R_X5Y126_SLICE_X7Y126_DO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_AMUX = CLBLM_R_X5Y126_SLICE_X7Y126_AO5;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_BMUX = CLBLM_R_X5Y126_SLICE_X7Y126_B5Q;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A = CLBLM_R_X5Y127_SLICE_X6Y127_AO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B = CLBLM_R_X5Y127_SLICE_X6Y127_BO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C = CLBLM_R_X5Y127_SLICE_X6Y127_CO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D = CLBLM_R_X5Y127_SLICE_X6Y127_DO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_AMUX = CLBLM_R_X5Y127_SLICE_X6Y127_AO5;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_BMUX = CLBLM_R_X5Y127_SLICE_X6Y127_B5Q;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_CMUX = CLBLM_R_X5Y127_SLICE_X6Y127_CO5;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A = CLBLM_R_X5Y127_SLICE_X7Y127_AO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B = CLBLM_R_X5Y127_SLICE_X7Y127_BO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C = CLBLM_R_X5Y127_SLICE_X7Y127_CO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D = CLBLM_R_X5Y127_SLICE_X7Y127_DO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_AMUX = CLBLM_R_X5Y127_SLICE_X7Y127_AO5;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_BMUX = CLBLM_R_X5Y127_SLICE_X7Y127_B5Q;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A = CLBLM_R_X5Y128_SLICE_X6Y128_AO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B = CLBLM_R_X5Y128_SLICE_X6Y128_BO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C = CLBLM_R_X5Y128_SLICE_X6Y128_CO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D = CLBLM_R_X5Y128_SLICE_X6Y128_DO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_AMUX = CLBLM_R_X5Y128_SLICE_X6Y128_AO5;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A = CLBLM_R_X5Y128_SLICE_X7Y128_AO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B = CLBLM_R_X5Y128_SLICE_X7Y128_BO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C = CLBLM_R_X5Y128_SLICE_X7Y128_CO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D = CLBLM_R_X5Y128_SLICE_X7Y128_DO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A = CLBLM_R_X5Y129_SLICE_X6Y129_AO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B = CLBLM_R_X5Y129_SLICE_X6Y129_BO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C = CLBLM_R_X5Y129_SLICE_X6Y129_CO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D = CLBLM_R_X5Y129_SLICE_X6Y129_DO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_AMUX = CLBLM_R_X5Y129_SLICE_X6Y129_A5Q;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A = CLBLM_R_X5Y129_SLICE_X7Y129_AO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B = CLBLM_R_X5Y129_SLICE_X7Y129_BO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C = CLBLM_R_X5Y129_SLICE_X7Y129_CO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D = CLBLM_R_X5Y129_SLICE_X7Y129_DO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_AMUX = CLBLM_R_X5Y129_SLICE_X7Y129_AO5;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_BMUX = CLBLM_R_X5Y129_SLICE_X7Y129_B5Q;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A = CLBLM_R_X5Y130_SLICE_X6Y130_AO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B = CLBLM_R_X5Y130_SLICE_X6Y130_BO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C = CLBLM_R_X5Y130_SLICE_X6Y130_CO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D = CLBLM_R_X5Y130_SLICE_X6Y130_DO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_AMUX = CLBLM_R_X5Y130_SLICE_X6Y130_AO5;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_BMUX = CLBLM_R_X5Y130_SLICE_X6Y130_B5Q;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_DMUX = CLBLM_R_X5Y130_SLICE_X6Y130_DO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A = CLBLM_R_X5Y130_SLICE_X7Y130_AO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B = CLBLM_R_X5Y130_SLICE_X7Y130_BO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C = CLBLM_R_X5Y130_SLICE_X7Y130_CO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D = CLBLM_R_X5Y130_SLICE_X7Y130_DO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_AMUX = CLBLM_R_X5Y130_SLICE_X7Y130_A5Q;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A = CLBLM_R_X5Y131_SLICE_X6Y131_AO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B = CLBLM_R_X5Y131_SLICE_X6Y131_BO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C = CLBLM_R_X5Y131_SLICE_X6Y131_CO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D = CLBLM_R_X5Y131_SLICE_X6Y131_DO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_AMUX = CLBLM_R_X5Y131_SLICE_X6Y131_A5Q;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_BMUX = CLBLM_R_X5Y131_SLICE_X6Y131_BO5;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A = CLBLM_R_X5Y131_SLICE_X7Y131_AO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B = CLBLM_R_X5Y131_SLICE_X7Y131_BO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C = CLBLM_R_X5Y131_SLICE_X7Y131_CO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D = CLBLM_R_X5Y131_SLICE_X7Y131_DO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_AMUX = CLBLM_R_X5Y131_SLICE_X7Y131_A5Q;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_BMUX = CLBLM_R_X5Y131_SLICE_X7Y131_BO5;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A = CLBLM_R_X5Y132_SLICE_X6Y132_AO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B = CLBLM_R_X5Y132_SLICE_X6Y132_BO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C = CLBLM_R_X5Y132_SLICE_X6Y132_CO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D = CLBLM_R_X5Y132_SLICE_X6Y132_DO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_AMUX = CLBLM_R_X5Y132_SLICE_X6Y132_AO5;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_BMUX = CLBLM_R_X5Y132_SLICE_X6Y132_B5Q;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A = CLBLM_R_X5Y132_SLICE_X7Y132_AO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B = CLBLM_R_X5Y132_SLICE_X7Y132_BO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C = CLBLM_R_X5Y132_SLICE_X7Y132_CO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_AMUX = CLBLM_R_X5Y132_SLICE_X7Y132_A5Q;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_BMUX = CLBLM_R_X5Y132_SLICE_X7Y132_B5Q;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A = CLBLM_R_X5Y133_SLICE_X6Y133_AO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B = CLBLM_R_X5Y133_SLICE_X6Y133_BO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C = CLBLM_R_X5Y133_SLICE_X6Y133_CO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D = CLBLM_R_X5Y133_SLICE_X6Y133_DO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_AMUX = CLBLM_R_X5Y133_SLICE_X6Y133_AO5;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A = CLBLM_R_X5Y133_SLICE_X7Y133_AO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B = CLBLM_R_X5Y133_SLICE_X7Y133_BO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C = CLBLM_R_X5Y133_SLICE_X7Y133_CO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D = CLBLM_R_X5Y133_SLICE_X7Y133_DO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A = CLBLM_R_X5Y134_SLICE_X6Y134_AO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B = CLBLM_R_X5Y134_SLICE_X6Y134_BO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C = CLBLM_R_X5Y134_SLICE_X6Y134_CO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D = CLBLM_R_X5Y134_SLICE_X6Y134_DO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_AMUX = CLBLM_R_X5Y134_SLICE_X6Y134_AO5;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_BMUX = CLBLM_R_X5Y134_SLICE_X6Y134_BO5;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_DMUX = CLBLM_R_X5Y134_SLICE_X6Y134_DO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A = CLBLM_R_X5Y134_SLICE_X7Y134_AO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B = CLBLM_R_X5Y134_SLICE_X7Y134_BO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C = CLBLM_R_X5Y134_SLICE_X7Y134_CO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D = CLBLM_R_X5Y134_SLICE_X7Y134_DO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_AMUX = CLBLM_R_X5Y134_SLICE_X7Y134_A5Q;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A = CLBLM_R_X5Y135_SLICE_X6Y135_AO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B = CLBLM_R_X5Y135_SLICE_X6Y135_BO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C = CLBLM_R_X5Y135_SLICE_X6Y135_CO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D = CLBLM_R_X5Y135_SLICE_X6Y135_DO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A = CLBLM_R_X5Y135_SLICE_X7Y135_AO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B = CLBLM_R_X5Y135_SLICE_X7Y135_BO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C = CLBLM_R_X5Y135_SLICE_X7Y135_CO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D = CLBLM_R_X5Y135_SLICE_X7Y135_DO6;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A = CLBLM_R_X5Y136_SLICE_X6Y136_AO6;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B = CLBLM_R_X5Y136_SLICE_X6Y136_BO6;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C = CLBLM_R_X5Y136_SLICE_X6Y136_CO6;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D = CLBLM_R_X5Y136_SLICE_X6Y136_DO6;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_CMUX = CLBLM_R_X5Y136_SLICE_X6Y136_CO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A = CLBLM_R_X5Y136_SLICE_X7Y136_AO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B = CLBLM_R_X5Y136_SLICE_X7Y136_BO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C = CLBLM_R_X5Y136_SLICE_X7Y136_CO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D = CLBLM_R_X5Y136_SLICE_X7Y136_DO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_A = CLBLM_R_X5Y137_SLICE_X6Y137_AO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_B = CLBLM_R_X5Y137_SLICE_X6Y137_BO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_C = CLBLM_R_X5Y137_SLICE_X6Y137_CO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_D = CLBLM_R_X5Y137_SLICE_X6Y137_DO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_AMUX = CLBLM_R_X5Y137_SLICE_X6Y137_AO6;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_A = CLBLM_R_X5Y137_SLICE_X7Y137_AO6;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_B = CLBLM_R_X5Y137_SLICE_X7Y137_BO6;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_C = CLBLM_R_X5Y137_SLICE_X7Y137_CO6;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_D = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A = CLBLM_R_X5Y138_SLICE_X6Y138_AO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C = CLBLM_R_X5Y138_SLICE_X6Y138_CO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D = CLBLM_R_X5Y138_SLICE_X6Y138_DO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A = CLBLM_R_X5Y138_SLICE_X7Y138_AO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B = CLBLM_R_X5Y138_SLICE_X7Y138_BO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C = CLBLM_R_X5Y138_SLICE_X7Y138_CO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D = CLBLM_R_X5Y138_SLICE_X7Y138_DO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A = CLBLM_R_X5Y139_SLICE_X6Y139_AO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B = CLBLM_R_X5Y139_SLICE_X6Y139_BO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C = CLBLM_R_X5Y139_SLICE_X6Y139_CO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D = CLBLM_R_X5Y139_SLICE_X6Y139_DO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_BMUX = CLBLM_R_X5Y139_SLICE_X6Y139_BO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A = CLBLM_R_X5Y139_SLICE_X7Y139_AO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B = CLBLM_R_X5Y139_SLICE_X7Y139_BO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C = CLBLM_R_X5Y139_SLICE_X7Y139_CO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D = CLBLM_R_X5Y139_SLICE_X7Y139_DO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A = CLBLM_R_X5Y140_SLICE_X6Y140_AO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B = CLBLM_R_X5Y140_SLICE_X6Y140_BO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C = CLBLM_R_X5Y140_SLICE_X6Y140_CO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D = CLBLM_R_X5Y140_SLICE_X6Y140_DO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A = CLBLM_R_X5Y140_SLICE_X7Y140_AO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B = CLBLM_R_X5Y140_SLICE_X7Y140_BO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C = CLBLM_R_X5Y140_SLICE_X7Y140_CO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D = CLBLM_R_X5Y140_SLICE_X7Y140_DO6;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_A = CLBLM_R_X5Y158_SLICE_X6Y158_AO6;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_B = CLBLM_R_X5Y158_SLICE_X6Y158_BO6;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_C = CLBLM_R_X5Y158_SLICE_X6Y158_CO6;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_D = CLBLM_R_X5Y158_SLICE_X6Y158_DO6;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_A = CLBLM_R_X5Y158_SLICE_X7Y158_AO6;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_B = CLBLM_R_X5Y158_SLICE_X7Y158_BO6;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_C = CLBLM_R_X5Y158_SLICE_X7Y158_CO6;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_D = CLBLM_R_X5Y158_SLICE_X7Y158_DO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A = CLBLM_R_X7Y125_SLICE_X8Y125_AO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B = CLBLM_R_X7Y125_SLICE_X8Y125_BO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C = CLBLM_R_X7Y125_SLICE_X8Y125_CO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D = CLBLM_R_X7Y125_SLICE_X8Y125_DO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_BMUX = CLBLM_R_X7Y125_SLICE_X8Y125_B5Q;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_CMUX = CLBLM_R_X7Y125_SLICE_X8Y125_C5Q;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A = CLBLM_R_X7Y125_SLICE_X9Y125_AO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B = CLBLM_R_X7Y125_SLICE_X9Y125_BO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C = CLBLM_R_X7Y125_SLICE_X9Y125_CO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D = CLBLM_R_X7Y125_SLICE_X9Y125_DO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A = CLBLM_R_X7Y126_SLICE_X8Y126_AO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B = CLBLM_R_X7Y126_SLICE_X8Y126_BO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C = CLBLM_R_X7Y126_SLICE_X8Y126_CO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D = CLBLM_R_X7Y126_SLICE_X8Y126_DO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_DMUX = CLBLM_R_X7Y126_SLICE_X8Y126_D5Q;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A = CLBLM_R_X7Y126_SLICE_X9Y126_AO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B = CLBLM_R_X7Y126_SLICE_X9Y126_BO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C = CLBLM_R_X7Y126_SLICE_X9Y126_CO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D = CLBLM_R_X7Y126_SLICE_X9Y126_DO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A = CLBLM_R_X7Y127_SLICE_X8Y127_AO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B = CLBLM_R_X7Y127_SLICE_X8Y127_BO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C = CLBLM_R_X7Y127_SLICE_X8Y127_CO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D = CLBLM_R_X7Y127_SLICE_X8Y127_DO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_AMUX = CLBLM_R_X7Y127_SLICE_X8Y127_A5Q;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A = CLBLM_R_X7Y127_SLICE_X9Y127_AO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B = CLBLM_R_X7Y127_SLICE_X9Y127_BO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C = CLBLM_R_X7Y127_SLICE_X9Y127_CO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D = CLBLM_R_X7Y127_SLICE_X9Y127_DO6;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A = CLBLM_R_X7Y128_SLICE_X8Y128_AO6;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B = CLBLM_R_X7Y128_SLICE_X8Y128_BO6;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C = CLBLM_R_X7Y128_SLICE_X8Y128_CO6;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D = CLBLM_R_X7Y128_SLICE_X8Y128_DO6;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_AMUX = CLBLM_R_X7Y128_SLICE_X8Y128_A5Q;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A = CLBLM_R_X7Y128_SLICE_X9Y128_AO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B = CLBLM_R_X7Y128_SLICE_X9Y128_BO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C = CLBLM_R_X7Y128_SLICE_X9Y128_CO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D = CLBLM_R_X7Y128_SLICE_X9Y128_DO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A = CLBLM_R_X7Y129_SLICE_X8Y129_AO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B = CLBLM_R_X7Y129_SLICE_X8Y129_BO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C = CLBLM_R_X7Y129_SLICE_X8Y129_CO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D = CLBLM_R_X7Y129_SLICE_X8Y129_DO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_AMUX = CLBLM_R_X7Y129_SLICE_X8Y129_A5Q;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_BMUX = CLBLM_R_X7Y129_SLICE_X8Y129_B5Q;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A = CLBLM_R_X7Y129_SLICE_X9Y129_AO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B = CLBLM_R_X7Y129_SLICE_X9Y129_BO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C = CLBLM_R_X7Y129_SLICE_X9Y129_CO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D = CLBLM_R_X7Y129_SLICE_X9Y129_DO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_AMUX = CLBLM_R_X7Y129_SLICE_X9Y129_A5Q;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_BMUX = CLBLM_R_X7Y129_SLICE_X9Y129_B5Q;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A = CLBLM_R_X7Y130_SLICE_X8Y130_AO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B = CLBLM_R_X7Y130_SLICE_X8Y130_BO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C = CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D = CLBLM_R_X7Y130_SLICE_X8Y130_DO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_AMUX = CLBLM_R_X7Y130_SLICE_X8Y130_AO5;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_BMUX = CLBLM_R_X7Y130_SLICE_X8Y130_B5Q;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A = CLBLM_R_X7Y130_SLICE_X9Y130_AO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B = CLBLM_R_X7Y130_SLICE_X9Y130_BO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C = CLBLM_R_X7Y130_SLICE_X9Y130_CO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D = CLBLM_R_X7Y130_SLICE_X9Y130_DO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A = CLBLM_R_X7Y131_SLICE_X8Y131_AO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B = CLBLM_R_X7Y131_SLICE_X8Y131_BO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C = CLBLM_R_X7Y131_SLICE_X8Y131_CO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D = CLBLM_R_X7Y131_SLICE_X8Y131_DO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_AMUX = CLBLM_R_X7Y131_SLICE_X8Y131_AO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A = CLBLM_R_X7Y131_SLICE_X9Y131_AO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B = CLBLM_R_X7Y131_SLICE_X9Y131_BO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C = CLBLM_R_X7Y131_SLICE_X9Y131_CO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D = CLBLM_R_X7Y131_SLICE_X9Y131_DO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_AMUX = CLBLM_R_X7Y131_SLICE_X9Y131_A5Q;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A = CLBLM_R_X7Y132_SLICE_X8Y132_AO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B = CLBLM_R_X7Y132_SLICE_X8Y132_BO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C = CLBLM_R_X7Y132_SLICE_X8Y132_CO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D = CLBLM_R_X7Y132_SLICE_X8Y132_DO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_AMUX = CLBLM_R_X7Y132_SLICE_X8Y132_A5Q;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A = CLBLM_R_X7Y132_SLICE_X9Y132_AO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B = CLBLM_R_X7Y132_SLICE_X9Y132_BO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C = CLBLM_R_X7Y132_SLICE_X9Y132_CO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D = CLBLM_R_X7Y132_SLICE_X9Y132_DO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_BMUX = CLBLM_R_X7Y132_SLICE_X9Y132_BO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A = CLBLM_R_X7Y133_SLICE_X8Y133_AO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B = CLBLM_R_X7Y133_SLICE_X8Y133_BO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C = CLBLM_R_X7Y133_SLICE_X8Y133_CO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D = CLBLM_R_X7Y133_SLICE_X8Y133_DO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A = CLBLM_R_X7Y133_SLICE_X9Y133_AO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C = CLBLM_R_X7Y133_SLICE_X9Y133_CO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D = CLBLM_R_X7Y133_SLICE_X9Y133_DO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A = CLBLM_R_X7Y134_SLICE_X8Y134_AO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B = CLBLM_R_X7Y134_SLICE_X8Y134_BO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C = CLBLM_R_X7Y134_SLICE_X8Y134_CO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D = CLBLM_R_X7Y134_SLICE_X8Y134_DO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_AMUX = CLBLM_R_X7Y134_SLICE_X8Y134_AO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_DMUX = CLBLM_R_X7Y134_SLICE_X8Y134_DO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A = CLBLM_R_X7Y134_SLICE_X9Y134_AO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B = CLBLM_R_X7Y134_SLICE_X9Y134_BO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C = CLBLM_R_X7Y134_SLICE_X9Y134_CO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D = CLBLM_R_X7Y134_SLICE_X9Y134_DO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_AMUX = CLBLM_R_X7Y134_SLICE_X9Y134_A5Q;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_BMUX = CLBLM_R_X7Y134_SLICE_X9Y134_B5Q;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A = CLBLM_R_X7Y135_SLICE_X8Y135_AO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B = CLBLM_R_X7Y135_SLICE_X8Y135_BO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C = CLBLM_R_X7Y135_SLICE_X8Y135_CO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D = CLBLM_R_X7Y135_SLICE_X8Y135_DO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A = CLBLM_R_X7Y135_SLICE_X9Y135_AO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B = CLBLM_R_X7Y135_SLICE_X9Y135_BO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C = CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D = CLBLM_R_X7Y135_SLICE_X9Y135_DO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_CMUX = CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A = CLBLM_R_X7Y136_SLICE_X8Y136_AO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B = CLBLM_R_X7Y136_SLICE_X8Y136_BO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C = CLBLM_R_X7Y136_SLICE_X8Y136_CO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D = CLBLM_R_X7Y136_SLICE_X8Y136_DO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_AMUX = CLBLM_R_X7Y136_SLICE_X8Y136_A5Q;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A = CLBLM_R_X7Y136_SLICE_X9Y136_AO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B = CLBLM_R_X7Y136_SLICE_X9Y136_BO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C = CLBLM_R_X7Y136_SLICE_X9Y136_CO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D = CLBLM_R_X7Y136_SLICE_X9Y136_DO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_AMUX = CLBLM_R_X7Y136_SLICE_X9Y136_AO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_BMUX = CLBLM_R_X7Y136_SLICE_X9Y136_BO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A = CLBLM_R_X7Y137_SLICE_X8Y137_AO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B = CLBLM_R_X7Y137_SLICE_X8Y137_BO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C = CLBLM_R_X7Y137_SLICE_X8Y137_CO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D = CLBLM_R_X7Y137_SLICE_X8Y137_DO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_AMUX = CLBLM_R_X7Y137_SLICE_X8Y137_A5Q;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A = CLBLM_R_X7Y137_SLICE_X9Y137_AO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B = CLBLM_R_X7Y137_SLICE_X9Y137_BO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C = CLBLM_R_X7Y137_SLICE_X9Y137_CO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D = CLBLM_R_X7Y137_SLICE_X9Y137_DO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_A = CLBLM_R_X7Y138_SLICE_X8Y138_AO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_B = CLBLM_R_X7Y138_SLICE_X8Y138_BO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_C = CLBLM_R_X7Y138_SLICE_X8Y138_CO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_D = CLBLM_R_X7Y138_SLICE_X8Y138_DO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_AMUX = CLBLM_R_X7Y138_SLICE_X8Y138_AO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_A = CLBLM_R_X7Y138_SLICE_X9Y138_AO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_B = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_C = CLBLM_R_X7Y138_SLICE_X9Y138_CO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_D = CLBLM_R_X7Y138_SLICE_X9Y138_DO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A = CLBLM_R_X7Y139_SLICE_X8Y139_AO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B = CLBLM_R_X7Y139_SLICE_X8Y139_BO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C = CLBLM_R_X7Y139_SLICE_X8Y139_CO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D = CLBLM_R_X7Y139_SLICE_X8Y139_DO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_DMUX = CLBLM_R_X7Y139_SLICE_X8Y139_DO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A = CLBLM_R_X7Y139_SLICE_X9Y139_AO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B = CLBLM_R_X7Y139_SLICE_X9Y139_BO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C = CLBLM_R_X7Y139_SLICE_X9Y139_CO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A = CLBLM_R_X7Y140_SLICE_X8Y140_AO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B = CLBLM_R_X7Y140_SLICE_X8Y140_BO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C = CLBLM_R_X7Y140_SLICE_X8Y140_CO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D = CLBLM_R_X7Y140_SLICE_X8Y140_DO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A = CLBLM_R_X7Y140_SLICE_X9Y140_AO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B = CLBLM_R_X7Y140_SLICE_X9Y140_BO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C = CLBLM_R_X7Y140_SLICE_X9Y140_CO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D = CLBLM_R_X7Y140_SLICE_X9Y140_DO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A = CLBLM_R_X11Y130_SLICE_X14Y130_AO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B = CLBLM_R_X11Y130_SLICE_X14Y130_BO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C = CLBLM_R_X11Y130_SLICE_X14Y130_CO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D = CLBLM_R_X11Y130_SLICE_X14Y130_DO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A = CLBLM_R_X11Y130_SLICE_X15Y130_AO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B = CLBLM_R_X11Y130_SLICE_X15Y130_BO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C = CLBLM_R_X11Y130_SLICE_X15Y130_CO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D = CLBLM_R_X11Y130_SLICE_X15Y130_DO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A = CLBLM_R_X11Y131_SLICE_X14Y131_AO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B = CLBLM_R_X11Y131_SLICE_X14Y131_BO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D = CLBLM_R_X11Y131_SLICE_X14Y131_DO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A = CLBLM_R_X11Y131_SLICE_X15Y131_AO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B = CLBLM_R_X11Y131_SLICE_X15Y131_BO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C = CLBLM_R_X11Y131_SLICE_X15Y131_CO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D = CLBLM_R_X11Y131_SLICE_X15Y131_DO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A = CLBLM_R_X11Y133_SLICE_X14Y133_AO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B = CLBLM_R_X11Y133_SLICE_X14Y133_BO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C = CLBLM_R_X11Y133_SLICE_X14Y133_CO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D = CLBLM_R_X11Y133_SLICE_X14Y133_DO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A = CLBLM_R_X11Y133_SLICE_X15Y133_AO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B = CLBLM_R_X11Y133_SLICE_X15Y133_BO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C = CLBLM_R_X11Y133_SLICE_X15Y133_CO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D = CLBLM_R_X11Y133_SLICE_X15Y133_DO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A = CLBLM_R_X11Y135_SLICE_X14Y135_AO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B = CLBLM_R_X11Y135_SLICE_X14Y135_BO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C = CLBLM_R_X11Y135_SLICE_X14Y135_CO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D = CLBLM_R_X11Y135_SLICE_X14Y135_DO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A = CLBLM_R_X11Y135_SLICE_X15Y135_AO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B = CLBLM_R_X11Y135_SLICE_X15Y135_BO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C = CLBLM_R_X11Y135_SLICE_X15Y135_CO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D = CLBLM_R_X11Y135_SLICE_X15Y135_DO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A = CLBLM_R_X11Y136_SLICE_X14Y136_AO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B = CLBLM_R_X11Y136_SLICE_X14Y136_BO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C = CLBLM_R_X11Y136_SLICE_X14Y136_CO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D = CLBLM_R_X11Y136_SLICE_X14Y136_DO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A = CLBLM_R_X11Y136_SLICE_X15Y136_AO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B = CLBLM_R_X11Y136_SLICE_X15Y136_BO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C = CLBLM_R_X11Y136_SLICE_X15Y136_CO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D = CLBLM_R_X11Y136_SLICE_X15Y136_DO6;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_A = CLBLM_R_X13Y135_SLICE_X18Y135_AO6;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_B = CLBLM_R_X13Y135_SLICE_X18Y135_BO6;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_C = CLBLM_R_X13Y135_SLICE_X18Y135_CO6;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_D = CLBLM_R_X13Y135_SLICE_X18Y135_DO6;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_AMUX = CLBLM_R_X13Y135_SLICE_X18Y135_AO6;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_A = CLBLM_R_X13Y135_SLICE_X19Y135_AO6;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_B = CLBLM_R_X13Y135_SLICE_X19Y135_BO6;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_C = CLBLM_R_X13Y135_SLICE_X19Y135_CO6;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_D = CLBLM_R_X13Y135_SLICE_X19Y135_DO6;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_A = CLBLM_R_X13Y136_SLICE_X18Y136_AO6;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_B = CLBLM_R_X13Y136_SLICE_X18Y136_BO6;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_C = CLBLM_R_X13Y136_SLICE_X18Y136_CO6;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_D = CLBLM_R_X13Y136_SLICE_X18Y136_DO6;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_A = CLBLM_R_X13Y136_SLICE_X19Y136_AO6;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_B = CLBLM_R_X13Y136_SLICE_X19Y136_BO6;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_C = CLBLM_R_X13Y136_SLICE_X19Y136_CO6;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_D = CLBLM_R_X13Y136_SLICE_X19Y136_DO6;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_A = CLBLM_R_X15Y135_SLICE_X20Y135_AO6;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_B = CLBLM_R_X15Y135_SLICE_X20Y135_BO6;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_C = CLBLM_R_X15Y135_SLICE_X20Y135_CO6;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_D = CLBLM_R_X15Y135_SLICE_X20Y135_DO6;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_A = CLBLM_R_X15Y135_SLICE_X21Y135_AO6;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_B = CLBLM_R_X15Y135_SLICE_X21Y135_BO6;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_C = CLBLM_R_X15Y135_SLICE_X21Y135_CO6;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_D = CLBLM_R_X15Y135_SLICE_X21Y135_DO6;
  assign CLBLM_R_X25Y149_SLICE_X36Y149_A = CLBLM_R_X25Y149_SLICE_X36Y149_AO6;
  assign CLBLM_R_X25Y149_SLICE_X36Y149_B = CLBLM_R_X25Y149_SLICE_X36Y149_BO6;
  assign CLBLM_R_X25Y149_SLICE_X36Y149_C = CLBLM_R_X25Y149_SLICE_X36Y149_CO6;
  assign CLBLM_R_X25Y149_SLICE_X36Y149_D = CLBLM_R_X25Y149_SLICE_X36Y149_DO6;
  assign CLBLM_R_X25Y149_SLICE_X37Y149_A = CLBLM_R_X25Y149_SLICE_X37Y149_AO6;
  assign CLBLM_R_X25Y149_SLICE_X37Y149_B = CLBLM_R_X25Y149_SLICE_X37Y149_BO6;
  assign CLBLM_R_X25Y149_SLICE_X37Y149_C = CLBLM_R_X25Y149_SLICE_X37Y149_CO6;
  assign CLBLM_R_X25Y149_SLICE_X37Y149_D = CLBLM_R_X25Y149_SLICE_X37Y149_DO6;
  assign CLBLM_R_X25Y151_SLICE_X36Y151_A = CLBLM_R_X25Y151_SLICE_X36Y151_AO6;
  assign CLBLM_R_X25Y151_SLICE_X36Y151_B = CLBLM_R_X25Y151_SLICE_X36Y151_BO6;
  assign CLBLM_R_X25Y151_SLICE_X36Y151_C = CLBLM_R_X25Y151_SLICE_X36Y151_CO6;
  assign CLBLM_R_X25Y151_SLICE_X36Y151_D = CLBLM_R_X25Y151_SLICE_X36Y151_DO6;
  assign CLBLM_R_X25Y151_SLICE_X37Y151_A = CLBLM_R_X25Y151_SLICE_X37Y151_AO6;
  assign CLBLM_R_X25Y151_SLICE_X37Y151_B = CLBLM_R_X25Y151_SLICE_X37Y151_BO6;
  assign CLBLM_R_X25Y151_SLICE_X37Y151_C = CLBLM_R_X25Y151_SLICE_X37Y151_CO6;
  assign CLBLM_R_X25Y151_SLICE_X37Y151_D = CLBLM_R_X25Y151_SLICE_X37Y151_DO6;
  assign CLBLM_R_X25Y153_SLICE_X36Y153_A = CLBLM_R_X25Y153_SLICE_X36Y153_AO6;
  assign CLBLM_R_X25Y153_SLICE_X36Y153_B = CLBLM_R_X25Y153_SLICE_X36Y153_BO6;
  assign CLBLM_R_X25Y153_SLICE_X36Y153_C = CLBLM_R_X25Y153_SLICE_X36Y153_CO6;
  assign CLBLM_R_X25Y153_SLICE_X36Y153_D = CLBLM_R_X25Y153_SLICE_X36Y153_DO6;
  assign CLBLM_R_X25Y153_SLICE_X37Y153_A = CLBLM_R_X25Y153_SLICE_X37Y153_AO6;
  assign CLBLM_R_X25Y153_SLICE_X37Y153_B = CLBLM_R_X25Y153_SLICE_X37Y153_BO6;
  assign CLBLM_R_X25Y153_SLICE_X37Y153_C = CLBLM_R_X25Y153_SLICE_X37Y153_CO6;
  assign CLBLM_R_X25Y153_SLICE_X37Y153_D = CLBLM_R_X25Y153_SLICE_X37Y153_DO6;
  assign CLBLM_R_X25Y154_SLICE_X36Y154_A = CLBLM_R_X25Y154_SLICE_X36Y154_AO6;
  assign CLBLM_R_X25Y154_SLICE_X36Y154_B = CLBLM_R_X25Y154_SLICE_X36Y154_BO6;
  assign CLBLM_R_X25Y154_SLICE_X36Y154_C = CLBLM_R_X25Y154_SLICE_X36Y154_CO6;
  assign CLBLM_R_X25Y154_SLICE_X36Y154_D = CLBLM_R_X25Y154_SLICE_X36Y154_DO6;
  assign CLBLM_R_X25Y154_SLICE_X37Y154_A = CLBLM_R_X25Y154_SLICE_X37Y154_AO6;
  assign CLBLM_R_X25Y154_SLICE_X37Y154_B = CLBLM_R_X25Y154_SLICE_X37Y154_BO6;
  assign CLBLM_R_X25Y154_SLICE_X37Y154_C = CLBLM_R_X25Y154_SLICE_X37Y154_CO6;
  assign CLBLM_R_X25Y154_SLICE_X37Y154_D = CLBLM_R_X25Y154_SLICE_X37Y154_DO6;
  assign CLBLM_R_X25Y157_SLICE_X36Y157_A = CLBLM_R_X25Y157_SLICE_X36Y157_AO6;
  assign CLBLM_R_X25Y157_SLICE_X36Y157_B = CLBLM_R_X25Y157_SLICE_X36Y157_BO6;
  assign CLBLM_R_X25Y157_SLICE_X36Y157_C = CLBLM_R_X25Y157_SLICE_X36Y157_CO6;
  assign CLBLM_R_X25Y157_SLICE_X36Y157_D = CLBLM_R_X25Y157_SLICE_X36Y157_DO6;
  assign CLBLM_R_X25Y157_SLICE_X37Y157_A = CLBLM_R_X25Y157_SLICE_X37Y157_AO6;
  assign CLBLM_R_X25Y157_SLICE_X37Y157_B = CLBLM_R_X25Y157_SLICE_X37Y157_BO6;
  assign CLBLM_R_X25Y157_SLICE_X37Y157_C = CLBLM_R_X25Y157_SLICE_X37Y157_CO6;
  assign CLBLM_R_X25Y157_SLICE_X37Y157_D = CLBLM_R_X25Y157_SLICE_X37Y157_DO6;
  assign LIOI3_X0Y1_ILOGIC_X0Y2_O = LIOB33_X0Y1_IOB_X0Y2_I;
  assign LIOI3_X0Y1_ILOGIC_X0Y1_O = LIOB33_X0Y1_IOB_X0Y1_I;
  assign LIOI3_X0Y3_ILOGIC_X0Y4_O = LIOB33_X0Y3_IOB_X0Y4_I;
  assign LIOI3_X0Y3_ILOGIC_X0Y3_O = LIOB33_X0Y3_IOB_X0Y3_I;
  assign LIOI3_X0Y5_ILOGIC_X0Y6_O = LIOB33_X0Y5_IOB_X0Y6_I;
  assign LIOI3_X0Y5_ILOGIC_X0Y5_O = LIOB33_X0Y5_IOB_X0Y5_I;
  assign LIOI3_X0Y9_ILOGIC_X0Y10_O = LIOB33_X0Y9_IOB_X0Y10_I;
  assign LIOI3_X0Y9_ILOGIC_X0Y9_O = LIOB33_X0Y9_IOB_X0Y9_I;
  assign LIOI3_X0Y11_ILOGIC_X0Y12_O = LIOB33_X0Y11_IOB_X0Y12_I;
  assign LIOI3_X0Y11_ILOGIC_X0Y11_O = LIOB33_X0Y11_IOB_X0Y11_I;
  assign LIOI3_X0Y15_ILOGIC_X0Y16_O = LIOB33_X0Y15_IOB_X0Y16_I;
  assign LIOI3_X0Y15_ILOGIC_X0Y15_O = LIOB33_X0Y15_IOB_X0Y15_I;
  assign LIOI3_X0Y17_ILOGIC_X0Y18_O = LIOB33_X0Y17_IOB_X0Y18_I;
  assign LIOI3_X0Y17_ILOGIC_X0Y17_O = LIOB33_X0Y17_IOB_X0Y17_I;
  assign LIOI3_X0Y21_ILOGIC_X0Y22_O = LIOB33_X0Y21_IOB_X0Y22_I;
  assign LIOI3_X0Y21_ILOGIC_X0Y21_O = LIOB33_X0Y21_IOB_X0Y21_I;
  assign LIOI3_X0Y23_ILOGIC_X0Y24_O = LIOB33_X0Y23_IOB_X0Y24_I;
  assign LIOI3_X0Y23_ILOGIC_X0Y23_O = LIOB33_X0Y23_IOB_X0Y23_I;
  assign LIOI3_X0Y25_ILOGIC_X0Y26_O = LIOB33_X0Y25_IOB_X0Y26_I;
  assign LIOI3_X0Y25_ILOGIC_X0Y25_O = LIOB33_X0Y25_IOB_X0Y25_I;
  assign LIOI3_X0Y27_ILOGIC_X0Y28_O = LIOB33_X0Y27_IOB_X0Y28_I;
  assign LIOI3_X0Y27_ILOGIC_X0Y27_O = LIOB33_X0Y27_IOB_X0Y27_I;
  assign LIOI3_X0Y29_ILOGIC_X0Y30_O = LIOB33_X0Y29_IOB_X0Y30_I;
  assign LIOI3_X0Y29_ILOGIC_X0Y29_O = LIOB33_X0Y29_IOB_X0Y29_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_O = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_O = LIOB33_X0Y51_IOB_X0Y51_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_O = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_O = LIOB33_X0Y53_IOB_X0Y53_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_O = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_O = LIOB33_X0Y55_IOB_X0Y55_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_O = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_O = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_O = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_O = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y66_O = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y65_O = LIOB33_X0Y65_IOB_X0Y65_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y68_O = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y67_O = LIOB33_X0Y67_IOB_X0Y67_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y72_O = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y71_O = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y74_O = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y73_O = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y76_O = LIOB33_X0Y75_IOB_X0Y76_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y75_O = LIOB33_X0Y75_IOB_X0Y75_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_O = LIOB33_X0Y77_IOB_X0Y78_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y77_O = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y79_ILOGIC_X0Y80_O = LIOB33_X0Y79_IOB_X0Y80_I;
  assign LIOI3_X0Y79_ILOGIC_X0Y79_O = LIOB33_X0Y79_IOB_X0Y79_I;
  assign LIOI3_X0Y83_ILOGIC_X0Y84_O = LIOB33_X0Y83_IOB_X0Y84_I;
  assign LIOI3_X0Y83_ILOGIC_X0Y83_O = LIOB33_X0Y83_IOB_X0Y83_I;
  assign LIOI3_X0Y85_ILOGIC_X0Y86_O = LIOB33_X0Y85_IOB_X0Y86_I;
  assign LIOI3_X0Y85_ILOGIC_X0Y85_O = LIOB33_X0Y85_IOB_X0Y85_I;
  assign LIOI3_X0Y89_ILOGIC_X0Y90_O = LIOB33_X0Y89_IOB_X0Y90_I;
  assign LIOI3_X0Y89_ILOGIC_X0Y89_O = LIOB33_X0Y89_IOB_X0Y89_I;
  assign LIOI3_X0Y91_ILOGIC_X0Y92_O = LIOB33_X0Y91_IOB_X0Y92_I;
  assign LIOI3_X0Y91_ILOGIC_X0Y91_O = LIOB33_X0Y91_IOB_X0Y91_I;
  assign LIOI3_X0Y95_ILOGIC_X0Y96_O = LIOB33_X0Y95_IOB_X0Y96_I;
  assign LIOI3_X0Y95_ILOGIC_X0Y95_O = LIOB33_X0Y95_IOB_X0Y95_I;
  assign LIOI3_X0Y97_ILOGIC_X0Y98_O = LIOB33_X0Y97_IOB_X0Y98_I;
  assign LIOI3_X0Y97_ILOGIC_X0Y97_O = LIOB33_X0Y97_IOB_X0Y97_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_O = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_O = LIOB33_X0Y101_IOB_X0Y101_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_O = LIOB33_X0Y103_IOB_X0Y104_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_O = LIOB33_X0Y103_IOB_X0Y103_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_O = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_O = LIOB33_X0Y105_IOB_X0Y105_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_O = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_O = LIOB33_X0Y109_IOB_X0Y109_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_O = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_O = LIOB33_X0Y111_IOB_X0Y111_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_O = LIOB33_X0Y115_IOB_X0Y116_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_O = LIOB33_X0Y115_IOB_X0Y115_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y118_O = LIOB33_X0Y117_IOB_X0Y118_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_O = LIOB33_X0Y117_IOB_X0Y117_I;
  assign LIOI3_X0Y121_ILOGIC_X0Y122_O = LIOB33_X0Y121_IOB_X0Y122_I;
  assign LIOI3_X0Y121_ILOGIC_X0Y121_O = LIOB33_X0Y121_IOB_X0Y121_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y124_O = LIOB33_X0Y123_IOB_X0Y124_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y123_O = LIOB33_X0Y123_IOB_X0Y123_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y126_O = LIOB33_X0Y125_IOB_X0Y126_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y125_O = LIOB33_X0Y125_IOB_X0Y125_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y128_O = LIOB33_X0Y127_IOB_X0Y128_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y127_O = LIOB33_X0Y127_IOB_X0Y127_I;
  assign LIOI3_X0Y129_ILOGIC_X0Y130_O = LIOB33_X0Y129_IOB_X0Y130_I;
  assign LIOI3_X0Y129_ILOGIC_X0Y129_O = LIOB33_X0Y129_IOB_X0Y129_I;
  assign LIOI3_X0Y133_ILOGIC_X0Y134_O = LIOB33_X0Y133_IOB_X0Y134_I;
  assign LIOI3_X0Y133_ILOGIC_X0Y133_O = LIOB33_X0Y133_IOB_X0Y133_I;
  assign LIOI3_X0Y135_ILOGIC_X0Y136_O = LIOB33_X0Y135_IOB_X0Y136_I;
  assign LIOI3_X0Y135_ILOGIC_X0Y135_O = LIOB33_X0Y135_IOB_X0Y135_I;
  assign LIOI3_X0Y139_ILOGIC_X0Y140_O = LIOB33_X0Y139_IOB_X0Y140_I;
  assign LIOI3_X0Y139_ILOGIC_X0Y139_O = LIOB33_X0Y139_IOB_X0Y139_I;
  assign LIOI3_X0Y141_ILOGIC_X0Y142_O = LIOB33_X0Y141_IOB_X0Y142_I;
  assign LIOI3_X0Y141_ILOGIC_X0Y141_O = LIOB33_X0Y141_IOB_X0Y141_I;
  assign LIOI3_X0Y145_ILOGIC_X0Y146_O = LIOB33_X0Y145_IOB_X0Y146_I;
  assign LIOI3_X0Y145_ILOGIC_X0Y145_O = LIOB33_X0Y145_IOB_X0Y145_I;
  assign LIOI3_X0Y147_ILOGIC_X0Y148_O = LIOB33_X0Y147_IOB_X0Y148_I;
  assign LIOI3_X0Y147_ILOGIC_X0Y147_O = LIOB33_X0Y147_IOB_X0Y147_I;
  assign LIOI3_X0Y151_ILOGIC_X0Y152_O = LIOB33_X0Y151_IOB_X0Y152_I;
  assign LIOI3_X0Y151_ILOGIC_X0Y151_O = LIOB33_X0Y151_IOB_X0Y151_I;
  assign LIOI3_X0Y153_ILOGIC_X0Y154_O = LIOB33_X0Y153_IOB_X0Y154_I;
  assign LIOI3_X0Y153_ILOGIC_X0Y153_O = LIOB33_X0Y153_IOB_X0Y153_I;
  assign LIOI3_X0Y155_ILOGIC_X0Y156_O = LIOB33_X0Y155_IOB_X0Y156_I;
  assign LIOI3_X0Y155_ILOGIC_X0Y155_O = LIOB33_X0Y155_IOB_X0Y155_I;
  assign LIOI3_X0Y159_ILOGIC_X0Y160_O = LIOB33_X0Y159_IOB_X0Y160_I;
  assign LIOI3_X0Y159_ILOGIC_X0Y159_O = LIOB33_X0Y159_IOB_X0Y159_I;
  assign LIOI3_X0Y161_ILOGIC_X0Y162_O = LIOB33_X0Y161_IOB_X0Y162_I;
  assign LIOI3_X0Y161_ILOGIC_X0Y161_O = LIOB33_X0Y161_IOB_X0Y161_I;
  assign LIOI3_X0Y165_ILOGIC_X0Y166_O = LIOB33_X0Y165_IOB_X0Y166_I;
  assign LIOI3_X0Y165_ILOGIC_X0Y165_O = LIOB33_X0Y165_IOB_X0Y165_I;
  assign LIOI3_X0Y167_ILOGIC_X0Y168_O = LIOB33_X0Y167_IOB_X0Y168_I;
  assign LIOI3_X0Y167_ILOGIC_X0Y167_O = LIOB33_X0Y167_IOB_X0Y167_I;
  assign LIOI3_X0Y171_ILOGIC_X0Y172_O = LIOB33_X0Y171_IOB_X0Y172_I;
  assign LIOI3_X0Y171_ILOGIC_X0Y171_O = LIOB33_X0Y171_IOB_X0Y171_I;
  assign LIOI3_X0Y173_ILOGIC_X0Y174_O = LIOB33_X0Y173_IOB_X0Y174_I;
  assign LIOI3_X0Y173_ILOGIC_X0Y173_O = LIOB33_X0Y173_IOB_X0Y173_I;
  assign LIOI3_X0Y175_ILOGIC_X0Y176_O = LIOB33_X0Y175_IOB_X0Y176_I;
  assign LIOI3_X0Y175_ILOGIC_X0Y175_O = LIOB33_X0Y175_IOB_X0Y175_I;
  assign LIOI3_X0Y177_ILOGIC_X0Y178_O = LIOB33_X0Y177_IOB_X0Y178_I;
  assign LIOI3_X0Y177_ILOGIC_X0Y177_O = LIOB33_X0Y177_IOB_X0Y177_I;
  assign LIOI3_X0Y179_ILOGIC_X0Y180_O = LIOB33_X0Y179_IOB_X0Y180_I;
  assign LIOI3_X0Y179_ILOGIC_X0Y179_O = LIOB33_X0Y179_IOB_X0Y179_I;
  assign LIOI3_X0Y183_ILOGIC_X0Y184_O = LIOB33_X0Y183_IOB_X0Y184_I;
  assign LIOI3_X0Y183_ILOGIC_X0Y183_O = LIOB33_X0Y183_IOB_X0Y183_I;
  assign LIOI3_X0Y185_ILOGIC_X0Y186_O = LIOB33_X0Y185_IOB_X0Y186_I;
  assign LIOI3_X0Y185_ILOGIC_X0Y185_O = LIOB33_X0Y185_IOB_X0Y185_I;
  assign LIOI3_X0Y189_ILOGIC_X0Y190_O = LIOB33_X0Y189_IOB_X0Y190_I;
  assign LIOI3_X0Y189_ILOGIC_X0Y189_O = LIOB33_X0Y189_IOB_X0Y189_I;
  assign LIOI3_X0Y191_ILOGIC_X0Y192_O = LIOB33_X0Y191_IOB_X0Y192_I;
  assign LIOI3_X0Y191_ILOGIC_X0Y191_O = LIOB33_X0Y191_IOB_X0Y191_I;
  assign LIOI3_X0Y195_ILOGIC_X0Y196_O = LIOB33_X0Y195_IOB_X0Y196_I;
  assign LIOI3_X0Y195_ILOGIC_X0Y195_O = LIOB33_X0Y195_IOB_X0Y195_I;
  assign LIOI3_X0Y197_ILOGIC_X0Y198_O = LIOB33_X0Y197_IOB_X0Y198_I;
  assign LIOI3_X0Y197_ILOGIC_X0Y197_O = LIOB33_X0Y197_IOB_X0Y197_I;
  assign LIOI3_X0Y201_ILOGIC_X0Y202_O = LIOB33_X0Y201_IOB_X0Y202_I;
  assign LIOI3_X0Y201_ILOGIC_X0Y201_O = LIOB33_X0Y201_IOB_X0Y201_I;
  assign LIOI3_X0Y203_ILOGIC_X0Y204_O = LIOB33_X0Y203_IOB_X0Y204_I;
  assign LIOI3_X0Y203_ILOGIC_X0Y203_O = LIOB33_X0Y203_IOB_X0Y203_I;
  assign LIOI3_X0Y205_ILOGIC_X0Y206_O = LIOB33_X0Y205_IOB_X0Y206_I;
  assign LIOI3_X0Y205_ILOGIC_X0Y205_O = LIOB33_X0Y205_IOB_X0Y205_I;
  assign LIOI3_X0Y209_ILOGIC_X0Y210_O = LIOB33_X0Y209_IOB_X0Y210_I;
  assign LIOI3_X0Y209_ILOGIC_X0Y209_O = LIOB33_X0Y209_IOB_X0Y209_I;
  assign LIOI3_X0Y211_ILOGIC_X0Y212_O = LIOB33_X0Y211_IOB_X0Y212_I;
  assign LIOI3_X0Y211_ILOGIC_X0Y211_O = LIOB33_X0Y211_IOB_X0Y211_I;
  assign LIOI3_X0Y215_ILOGIC_X0Y216_O = LIOB33_X0Y215_IOB_X0Y216_I;
  assign LIOI3_X0Y215_ILOGIC_X0Y215_O = LIOB33_X0Y215_IOB_X0Y215_I;
  assign LIOI3_X0Y217_ILOGIC_X0Y218_O = LIOB33_X0Y217_IOB_X0Y218_I;
  assign LIOI3_X0Y217_ILOGIC_X0Y217_O = LIOB33_X0Y217_IOB_X0Y217_I;
  assign LIOI3_X0Y221_ILOGIC_X0Y222_O = LIOB33_X0Y221_IOB_X0Y222_I;
  assign LIOI3_X0Y221_ILOGIC_X0Y221_O = LIOB33_X0Y221_IOB_X0Y221_I;
  assign LIOI3_X0Y223_ILOGIC_X0Y224_O = LIOB33_X0Y223_IOB_X0Y224_I;
  assign LIOI3_X0Y223_ILOGIC_X0Y223_O = LIOB33_X0Y223_IOB_X0Y223_I;
  assign LIOI3_X0Y225_ILOGIC_X0Y226_O = LIOB33_X0Y225_IOB_X0Y226_I;
  assign LIOI3_X0Y225_ILOGIC_X0Y225_O = LIOB33_X0Y225_IOB_X0Y225_I;
  assign LIOI3_X0Y227_ILOGIC_X0Y228_O = LIOB33_X0Y227_IOB_X0Y228_I;
  assign LIOI3_X0Y227_ILOGIC_X0Y227_O = LIOB33_X0Y227_IOB_X0Y227_I;
  assign LIOI3_X0Y229_ILOGIC_X0Y230_O = LIOB33_X0Y229_IOB_X0Y230_I;
  assign LIOI3_X0Y229_ILOGIC_X0Y229_O = LIOB33_X0Y229_IOB_X0Y229_I;
  assign LIOI3_X0Y233_ILOGIC_X0Y234_O = LIOB33_X0Y233_IOB_X0Y234_I;
  assign LIOI3_X0Y233_ILOGIC_X0Y233_O = LIOB33_X0Y233_IOB_X0Y233_I;
  assign LIOI3_X0Y235_ILOGIC_X0Y236_O = LIOB33_X0Y235_IOB_X0Y236_I;
  assign LIOI3_X0Y235_ILOGIC_X0Y235_O = LIOB33_X0Y235_IOB_X0Y235_I;
  assign LIOI3_X0Y239_ILOGIC_X0Y240_O = LIOB33_X0Y239_IOB_X0Y240_I;
  assign LIOI3_X0Y239_ILOGIC_X0Y239_O = LIOB33_X0Y239_IOB_X0Y239_I;
  assign LIOI3_X0Y241_ILOGIC_X0Y242_O = LIOB33_X0Y241_IOB_X0Y242_I;
  assign LIOI3_X0Y241_ILOGIC_X0Y241_O = LIOB33_X0Y241_IOB_X0Y241_I;
  assign LIOI3_X0Y245_ILOGIC_X0Y246_O = LIOB33_X0Y245_IOB_X0Y246_I;
  assign LIOI3_X0Y245_ILOGIC_X0Y245_O = LIOB33_X0Y245_IOB_X0Y245_I;
  assign LIOI3_X0Y247_ILOGIC_X0Y248_O = LIOB33_X0Y247_IOB_X0Y248_I;
  assign LIOI3_X0Y247_ILOGIC_X0Y247_O = LIOB33_X0Y247_IOB_X0Y247_I;
  assign LIOI3_SING_X0Y0_ILOGIC_X0Y0_O = LIOB33_SING_X0Y0_IOB_X0Y0_I;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_SING_X0Y99_ILOGIC_X0Y99_O = LIOB33_SING_X0Y99_IOB_X0Y99_I;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ = CLBLL_L_X2Y141_SLICE_X0Y141_AQ;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ = 1'b1;
  assign LIOI3_SING_X0Y149_ILOGIC_X0Y149_O = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign LIOI3_SING_X0Y150_ILOGIC_X0Y150_O = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign LIOI3_SING_X0Y199_ILOGIC_X0Y199_O = LIOB33_SING_X0Y199_IOB_X0Y199_I;
  assign LIOI3_SING_X0Y200_ILOGIC_X0Y200_O = LIOB33_SING_X0Y200_IOB_X0Y200_I;
  assign LIOI3_SING_X0Y249_ILOGIC_X0Y249_O = LIOB33_SING_X0Y249_IOB_X0Y249_I;
  assign LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y8_O = LIOB33_X0Y7_IOB_X0Y8_I;
  assign LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y7_O = LIOB33_X0Y7_IOB_X0Y7_I;
  assign LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y20_O = LIOB33_X0Y19_IOB_X0Y20_I;
  assign LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y19_O = LIOB33_X0Y19_IOB_X0Y19_I;
  assign LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y31_O = LIOB33_X0Y31_IOB_X0Y31_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_O = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_O = LIOB33_X0Y69_IOB_X0Y69_I;
  assign LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y82_O = LIOB33_X0Y81_IOB_X0Y82_I;
  assign LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y81_O = LIOB33_X0Y81_IOB_X0Y81_I;
  assign LIOI3_TBYTESRC_X0Y93_ILOGIC_X0Y94_O = LIOB33_X0Y93_IOB_X0Y94_I;
  assign LIOI3_TBYTESRC_X0Y93_ILOGIC_X0Y93_O = LIOB33_X0Y93_IOB_X0Y93_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O = LIOB33_X0Y107_IOB_X0Y107_I;
  assign LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_O = LIOB33_X0Y119_IOB_X0Y120_I;
  assign LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y119_O = LIOB33_X0Y119_IOB_X0Y119_I;
  assign LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y132_O = LIOB33_X0Y131_IOB_X0Y132_I;
  assign LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y131_O = LIOB33_X0Y131_IOB_X0Y131_I;
  assign LIOI3_TBYTESRC_X0Y143_ILOGIC_X0Y144_O = LIOI3_TBYTESRC_X0Y143_ILOGIC_X0Y144_D;
  assign LIOI3_TBYTESRC_X0Y143_ILOGIC_X0Y143_O = LIOB33_X0Y143_IOB_X0Y143_I;
  assign LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y158_O = LIOB33_X0Y157_IOB_X0Y158_I;
  assign LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y157_O = LIOB33_X0Y157_IOB_X0Y157_I;
  assign LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y170_O = LIOB33_X0Y169_IOB_X0Y170_I;
  assign LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y169_O = LIOB33_X0Y169_IOB_X0Y169_I;
  assign LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y182_O = LIOB33_X0Y181_IOB_X0Y182_I;
  assign LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y181_O = LIOB33_X0Y181_IOB_X0Y181_I;
  assign LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y194_O = LIOB33_X0Y193_IOB_X0Y194_I;
  assign LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y193_O = LIOB33_X0Y193_IOB_X0Y193_I;
  assign LIOI3_TBYTESRC_X0Y207_ILOGIC_X0Y208_O = LIOB33_X0Y207_IOB_X0Y208_I;
  assign LIOI3_TBYTESRC_X0Y207_ILOGIC_X0Y207_O = LIOB33_X0Y207_IOB_X0Y207_I;
  assign LIOI3_TBYTESRC_X0Y219_ILOGIC_X0Y220_O = LIOB33_X0Y219_IOB_X0Y220_I;
  assign LIOI3_TBYTESRC_X0Y219_ILOGIC_X0Y219_O = LIOB33_X0Y219_IOB_X0Y219_I;
  assign LIOI3_TBYTESRC_X0Y231_ILOGIC_X0Y232_O = LIOB33_X0Y231_IOB_X0Y232_I;
  assign LIOI3_TBYTESRC_X0Y231_ILOGIC_X0Y231_O = LIOB33_X0Y231_IOB_X0Y231_I;
  assign LIOI3_TBYTESRC_X0Y243_ILOGIC_X0Y244_O = LIOB33_X0Y243_IOB_X0Y244_I;
  assign LIOI3_TBYTESRC_X0Y243_ILOGIC_X0Y243_O = LIOB33_X0Y243_IOB_X0Y243_I;
  assign LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y14_O = LIOB33_X0Y13_IOB_X0Y14_I;
  assign LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y13_O = LIOB33_X0Y13_IOB_X0Y13_I;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_O = LIOB33_X0Y63_IOB_X0Y64_I;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_TBYTETERM_X0Y87_ILOGIC_X0Y88_O = LIOB33_X0Y87_IOB_X0Y88_I;
  assign LIOI3_TBYTETERM_X0Y87_ILOGIC_X0Y87_O = LIOB33_X0Y87_IOB_X0Y87_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O = LIOB33_X0Y113_IOB_X0Y114_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O = LIOB33_X0Y113_IOB_X0Y113_I;
  assign LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y138_O = LIOB33_X0Y137_IOB_X0Y138_I;
  assign LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_O = LIOB33_X0Y137_IOB_X0Y137_I;
  assign LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y164_O = LIOB33_X0Y163_IOB_X0Y164_I;
  assign LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y163_O = LIOB33_X0Y163_IOB_X0Y163_I;
  assign LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y188_O = LIOB33_X0Y187_IOB_X0Y188_I;
  assign LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y187_O = LIOB33_X0Y187_IOB_X0Y187_I;
  assign LIOI3_TBYTETERM_X0Y213_ILOGIC_X0Y214_O = LIOB33_X0Y213_IOB_X0Y214_I;
  assign LIOI3_TBYTETERM_X0Y213_ILOGIC_X0Y213_O = LIOB33_X0Y213_IOB_X0Y213_I;
  assign LIOI3_TBYTETERM_X0Y237_ILOGIC_X0Y238_O = LIOB33_X0Y237_IOB_X0Y238_I;
  assign LIOI3_TBYTETERM_X0Y237_ILOGIC_X0Y237_O = LIOB33_X0Y237_IOB_X0Y237_I;
  assign RIOI3_X105Y51_OLOGIC_X1Y52_OQ = CLBLM_R_X5Y134_SLICE_X7Y134_CQ;
  assign RIOI3_X105Y51_OLOGIC_X1Y52_TQ = 1'b1;
  assign RIOI3_X105Y51_OLOGIC_X1Y51_OQ = CLBLM_R_X5Y132_SLICE_X7Y132_BQ;
  assign RIOI3_X105Y51_OLOGIC_X1Y51_TQ = 1'b1;
  assign RIOI3_X105Y53_OLOGIC_X1Y54_OQ = CLBLM_R_X7Y132_SLICE_X9Y132_AQ;
  assign RIOI3_X105Y53_OLOGIC_X1Y54_TQ = 1'b1;
  assign RIOI3_X105Y53_OLOGIC_X1Y53_OQ = CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  assign RIOI3_X105Y53_OLOGIC_X1Y53_TQ = 1'b1;
  assign RIOI3_X105Y55_OLOGIC_X1Y56_OQ = CLBLM_R_X5Y133_SLICE_X7Y133_CQ;
  assign RIOI3_X105Y55_OLOGIC_X1Y56_TQ = 1'b1;
  assign RIOI3_X105Y55_OLOGIC_X1Y55_OQ = CLBLL_L_X4Y134_SLICE_X5Y134_AQ;
  assign RIOI3_X105Y55_OLOGIC_X1Y55_TQ = 1'b1;
  assign RIOI3_X105Y59_OLOGIC_X1Y60_OQ = CLBLM_R_X7Y136_SLICE_X8Y136_BQ;
  assign RIOI3_X105Y59_OLOGIC_X1Y60_TQ = 1'b1;
  assign RIOI3_X105Y59_OLOGIC_X1Y59_OQ = CLBLM_R_X5Y131_SLICE_X6Y131_AQ;
  assign RIOI3_X105Y59_OLOGIC_X1Y59_TQ = 1'b1;
  assign RIOI3_X105Y61_OLOGIC_X1Y62_OQ = CLBLL_L_X4Y134_SLICE_X5Y134_BQ;
  assign RIOI3_X105Y61_OLOGIC_X1Y62_TQ = 1'b1;
  assign RIOI3_X105Y61_OLOGIC_X1Y61_OQ = CLBLL_L_X4Y135_SLICE_X5Y135_BQ;
  assign RIOI3_X105Y61_OLOGIC_X1Y61_TQ = 1'b1;
  assign RIOI3_X105Y65_OLOGIC_X1Y66_OQ = CLBLM_R_X7Y125_SLICE_X8Y125_AQ;
  assign RIOI3_X105Y65_OLOGIC_X1Y66_TQ = 1'b1;
  assign RIOI3_X105Y65_OLOGIC_X1Y65_OQ = CLBLM_L_X8Y127_SLICE_X10Y127_AQ;
  assign RIOI3_X105Y65_OLOGIC_X1Y65_TQ = 1'b1;
  assign RIOI3_X105Y67_OLOGIC_X1Y68_OQ = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign RIOI3_X105Y67_OLOGIC_X1Y68_TQ = 1'b1;
  assign RIOI3_X105Y67_OLOGIC_X1Y67_OQ = CLBLM_L_X8Y127_SLICE_X10Y127_BQ;
  assign RIOI3_X105Y67_OLOGIC_X1Y67_TQ = 1'b1;
  assign RIOI3_X105Y71_OLOGIC_X1Y72_OQ = CLBLM_R_X7Y128_SLICE_X9Y128_AQ;
  assign RIOI3_X105Y71_OLOGIC_X1Y72_TQ = 1'b1;
  assign RIOI3_X105Y71_OLOGIC_X1Y71_OQ = CLBLL_L_X54Y101_SLICE_X82Y101_AQ;
  assign RIOI3_X105Y71_OLOGIC_X1Y71_TQ = 1'b1;
  assign RIOI3_X105Y73_OLOGIC_X1Y74_OQ = CLBLM_R_X7Y130_SLICE_X9Y130_DQ;
  assign RIOI3_X105Y73_OLOGIC_X1Y74_TQ = 1'b1;
  assign RIOI3_X105Y73_OLOGIC_X1Y73_OQ = CLBLM_L_X8Y130_SLICE_X11Y130_BQ;
  assign RIOI3_X105Y73_OLOGIC_X1Y73_TQ = 1'b1;
  assign RIOI3_X105Y75_OLOGIC_X1Y76_OQ = CLBLM_L_X10Y132_SLICE_X12Y132_AQ;
  assign RIOI3_X105Y75_OLOGIC_X1Y76_TQ = 1'b1;
  assign RIOI3_X105Y75_OLOGIC_X1Y75_OQ = CLBLM_L_X8Y130_SLICE_X10Y130_DQ;
  assign RIOI3_X105Y75_OLOGIC_X1Y75_TQ = 1'b1;
  assign RIOI3_X105Y77_OLOGIC_X1Y78_OQ = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign RIOI3_X105Y77_OLOGIC_X1Y78_TQ = 1'b1;
  assign RIOI3_X105Y77_OLOGIC_X1Y77_OQ = CLBLM_L_X8Y130_SLICE_X11Y130_CQ;
  assign RIOI3_X105Y77_OLOGIC_X1Y77_TQ = 1'b1;
  assign RIOI3_X105Y79_OLOGIC_X1Y80_OQ = CLBLM_L_X8Y131_SLICE_X11Y131_BQ;
  assign RIOI3_X105Y79_OLOGIC_X1Y80_TQ = 1'b1;
  assign RIOI3_X105Y79_OLOGIC_X1Y79_OQ = CLBLL_L_X54Y105_SLICE_X82Y105_AQ;
  assign RIOI3_X105Y79_OLOGIC_X1Y79_TQ = 1'b1;
  assign RIOI3_X105Y83_OLOGIC_X1Y84_OQ = CLBLM_L_X10Y132_SLICE_X12Y132_BQ;
  assign RIOI3_X105Y83_OLOGIC_X1Y84_TQ = 1'b1;
  assign RIOI3_X105Y83_OLOGIC_X1Y83_OQ = CLBLM_L_X8Y131_SLICE_X10Y131_BQ;
  assign RIOI3_X105Y83_OLOGIC_X1Y83_TQ = 1'b1;
  assign RIOI3_X105Y85_OLOGIC_X1Y86_OQ = CLBLM_L_X8Y132_SLICE_X11Y132_CQ;
  assign RIOI3_X105Y85_OLOGIC_X1Y86_TQ = 1'b1;
  assign RIOI3_X105Y85_OLOGIC_X1Y85_OQ = CLBLM_L_X10Y132_SLICE_X12Y132_CQ;
  assign RIOI3_X105Y85_OLOGIC_X1Y85_TQ = 1'b1;
  assign RIOI3_X105Y89_OLOGIC_X1Y90_OQ = CLBLM_L_X10Y130_SLICE_X12Y130_BQ;
  assign RIOI3_X105Y89_OLOGIC_X1Y90_TQ = 1'b1;
  assign RIOI3_X105Y89_OLOGIC_X1Y89_OQ = CLBLM_R_X11Y130_SLICE_X14Y130_AQ;
  assign RIOI3_X105Y89_OLOGIC_X1Y89_TQ = 1'b1;
  assign RIOI3_X105Y91_OLOGIC_X1Y92_OQ = CLBLM_R_X11Y131_SLICE_X14Y131_AQ;
  assign RIOI3_X105Y91_OLOGIC_X1Y92_TQ = 1'b1;
  assign RIOI3_X105Y91_OLOGIC_X1Y91_OQ = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign RIOI3_X105Y91_OLOGIC_X1Y91_TQ = 1'b1;
  assign RIOI3_X105Y95_OLOGIC_X1Y96_OQ = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign RIOI3_X105Y95_OLOGIC_X1Y96_TQ = 1'b1;
  assign RIOI3_X105Y95_OLOGIC_X1Y95_OQ = CLBLM_R_X11Y131_SLICE_X14Y131_BQ;
  assign RIOI3_X105Y95_OLOGIC_X1Y95_TQ = 1'b1;
  assign RIOI3_X105Y97_OLOGIC_X1Y98_OQ = CLBLM_R_X7Y125_SLICE_X8Y125_CQ;
  assign RIOI3_X105Y97_OLOGIC_X1Y98_TQ = 1'b1;
  assign RIOI3_X105Y97_OLOGIC_X1Y97_OQ = CLBLM_R_X7Y125_SLICE_X8Y125_BQ;
  assign RIOI3_X105Y97_OLOGIC_X1Y97_TQ = 1'b1;
  assign RIOI3_X105Y101_OLOGIC_X1Y102_OQ = CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  assign RIOI3_X105Y101_OLOGIC_X1Y102_TQ = 1'b1;
  assign RIOI3_X105Y101_OLOGIC_X1Y101_OQ = CLBLM_R_X7Y126_SLICE_X8Y126_AQ;
  assign RIOI3_X105Y101_OLOGIC_X1Y101_TQ = 1'b1;
  assign RIOI3_X105Y103_OLOGIC_X1Y104_OQ = CLBLM_R_X7Y128_SLICE_X8Y128_BQ;
  assign RIOI3_X105Y103_OLOGIC_X1Y104_TQ = 1'b1;
  assign RIOI3_X105Y103_OLOGIC_X1Y103_OQ = CLBLM_R_X7Y126_SLICE_X8Y126_CQ;
  assign RIOI3_X105Y103_OLOGIC_X1Y103_TQ = 1'b1;
  assign RIOI3_X105Y105_OLOGIC_X1Y106_OQ = CLBLM_R_X5Y131_SLICE_X7Y131_AQ;
  assign RIOI3_X105Y105_OLOGIC_X1Y106_TQ = 1'b1;
  assign RIOI3_X105Y105_OLOGIC_X1Y105_OQ = CLBLM_R_X7Y129_SLICE_X9Y129_CQ;
  assign RIOI3_X105Y105_OLOGIC_X1Y105_TQ = 1'b1;
  assign RIOI3_X105Y109_OLOGIC_X1Y110_OQ = CLBLM_R_X7Y129_SLICE_X8Y129_DQ;
  assign RIOI3_X105Y109_OLOGIC_X1Y110_TQ = 1'b1;
  assign RIOI3_X105Y109_OLOGIC_X1Y109_OQ = CLBLM_R_X7Y129_SLICE_X8Y129_CQ;
  assign RIOI3_X105Y109_OLOGIC_X1Y109_TQ = 1'b1;
  assign RIOI3_X105Y111_OLOGIC_X1Y112_OQ = CLBLM_R_X7Y131_SLICE_X9Y131_BQ;
  assign RIOI3_X105Y111_OLOGIC_X1Y112_TQ = 1'b1;
  assign RIOI3_X105Y111_OLOGIC_X1Y111_OQ = CLBLM_R_X7Y130_SLICE_X9Y130_AQ;
  assign RIOI3_X105Y111_OLOGIC_X1Y111_TQ = 1'b1;
  assign RIOI3_X105Y115_OLOGIC_X1Y116_OQ = CLBLM_L_X10Y133_SLICE_X13Y133_AQ;
  assign RIOI3_X105Y115_OLOGIC_X1Y116_TQ = 1'b1;
  assign RIOI3_X105Y115_OLOGIC_X1Y115_OQ = CLBLL_L_X54Y123_SLICE_X82Y123_AQ;
  assign RIOI3_X105Y115_OLOGIC_X1Y115_TQ = 1'b1;
  assign RIOI3_X105Y117_OLOGIC_X1Y118_OQ = CLBLM_L_X10Y131_SLICE_X12Y131_AQ;
  assign RIOI3_X105Y117_OLOGIC_X1Y118_TQ = 1'b1;
  assign RIOI3_X105Y117_OLOGIC_X1Y117_OQ = CLBLM_L_X12Y132_SLICE_X16Y132_AQ;
  assign RIOI3_X105Y117_OLOGIC_X1Y117_TQ = 1'b1;
  assign RIOI3_X105Y121_OLOGIC_X1Y122_OQ = CLBLM_L_X10Y133_SLICE_X13Y133_CQ;
  assign RIOI3_X105Y121_OLOGIC_X1Y122_TQ = 1'b1;
  assign RIOI3_X105Y121_OLOGIC_X1Y121_OQ = CLBLM_R_X11Y133_SLICE_X14Y133_BQ;
  assign RIOI3_X105Y121_OLOGIC_X1Y121_TQ = 1'b1;
  assign RIOI3_X105Y123_OLOGIC_X1Y124_OQ = CLBLM_R_X7Y130_SLICE_X9Y130_BQ;
  assign RIOI3_X105Y123_OLOGIC_X1Y124_TQ = 1'b1;
  assign RIOI3_X105Y123_OLOGIC_X1Y123_OQ = CLBLM_L_X12Y132_SLICE_X16Y132_BQ;
  assign RIOI3_X105Y123_OLOGIC_X1Y123_TQ = 1'b1;
  assign RIOI3_X105Y125_OLOGIC_X1Y126_OQ = CLBLM_R_X7Y130_SLICE_X9Y130_CQ;
  assign RIOI3_X105Y125_OLOGIC_X1Y126_TQ = 1'b1;
  assign RIOI3_X105Y125_OLOGIC_X1Y125_OQ = CLBLM_R_X5Y132_SLICE_X7Y132_AQ;
  assign RIOI3_X105Y125_OLOGIC_X1Y125_TQ = 1'b1;
  assign RIOI3_X105Y127_OLOGIC_X1Y128_OQ = CLBLM_L_X8Y134_SLICE_X10Y134_AQ;
  assign RIOI3_X105Y127_OLOGIC_X1Y128_TQ = 1'b1;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_OQ = CLBLM_R_X5Y133_SLICE_X7Y133_AQ;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_TQ = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_OQ = CLBLM_L_X8Y132_SLICE_X11Y132_BQ;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_TQ = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_OQ = CLBLM_R_X7Y133_SLICE_X9Y133_AQ;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_TQ = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_OQ = CLBLM_R_X5Y133_SLICE_X7Y133_BQ;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_TQ = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_OQ = CLBLM_R_X7Y133_SLICE_X9Y133_BQ;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_TQ = 1'b1;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_OQ = CLBLM_R_X5Y135_SLICE_X7Y135_AQ;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_TQ = 1'b1;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_OQ = CLBLM_R_X7Y137_SLICE_X9Y137_AQ;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_TQ = 1'b1;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_OQ = CLBLM_R_X7Y138_SLICE_X9Y138_AQ;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_TQ = 1'b1;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_OQ = CLBLL_L_X54Y138_SLICE_X82Y138_AQ;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_TQ = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_OQ = CLBLM_R_X7Y138_SLICE_X9Y138_CQ;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_TQ = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_OQ = CLBLM_R_X7Y138_SLICE_X9Y138_BQ;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_TQ = 1'b1;
  assign RIOI3_X105Y145_OLOGIC_X1Y146_OQ = CLBLM_R_X5Y138_SLICE_X7Y138_AQ;
  assign RIOI3_X105Y145_OLOGIC_X1Y146_TQ = 1'b1;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_OQ = CLBLM_R_X5Y138_SLICE_X6Y138_BQ;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_TQ = 1'b1;
  assign RIOI3_X105Y147_OLOGIC_X1Y148_OQ = CLBLM_R_X7Y137_SLICE_X9Y137_BQ;
  assign RIOI3_X105Y147_OLOGIC_X1Y148_TQ = 1'b1;
  assign RIOI3_X105Y147_OLOGIC_X1Y147_OQ = CLBLL_L_X54Y141_SLICE_X82Y141_AQ;
  assign RIOI3_X105Y147_OLOGIC_X1Y147_TQ = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_OQ = CLBLM_R_X7Y129_SLICE_X9Y129_BQ;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_TQ = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_OQ = CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_OQ = CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_OQ = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_OQ = CLBLM_R_X7Y129_SLICE_X8Y129_BQ;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_OQ = CLBLM_R_X7Y136_SLICE_X8Y136_AQ;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_OQ = CLBLM_R_X7Y137_SLICE_X8Y137_AQ;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_OQ = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_OQ = CLBLM_L_X8Y132_SLICE_X11Y132_AQ;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_OQ = CLBLM_R_X5Y134_SLICE_X7Y134_AQ;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_OQ = CLBLM_L_X8Y136_SLICE_X10Y136_AQ;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_OQ = CLBLM_R_X7Y134_SLICE_X9Y134_BQ;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_OQ = CLBLM_L_X8Y137_SLICE_X10Y137_AQ;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_OQ = CLBLM_L_X10Y135_SLICE_X12Y135_AQ;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_OQ = CLBLM_L_X16Y136_SLICE_X22Y136_AQ;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_OQ = CLBLM_R_X15Y135_SLICE_X21Y135_AQ;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_OQ = CLBLM_L_X16Y135_SLICE_X22Y135_BQ;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_OQ = CLBLM_L_X16Y135_SLICE_X22Y135_AQ;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_OQ = CLBLM_L_X16Y137_SLICE_X22Y137_AQ;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_OQ = CLBLM_R_X13Y136_SLICE_X18Y136_AQ;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_TQ = 1'b1;
  assign RIOI3_X105Y177_ILOGIC_X1Y178_O = RIOB33_X105Y177_IOB_X1Y178_I;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_OQ = CLBLM_L_X16Y137_SLICE_X22Y137_BQ;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_TQ = 1'b1;
  assign RIOI3_X105Y179_ILOGIC_X1Y180_O = RIOB33_X105Y179_IOB_X1Y180_I;
  assign RIOI3_X105Y179_ILOGIC_X1Y179_O = RIOB33_X105Y179_IOB_X1Y179_I;
  assign RIOI3_X105Y183_ILOGIC_X1Y184_O = RIOB33_X105Y183_IOB_X1Y184_I;
  assign RIOI3_X105Y183_ILOGIC_X1Y183_O = RIOB33_X105Y183_IOB_X1Y183_I;
  assign RIOI3_X105Y185_ILOGIC_X1Y186_O = RIOB33_X105Y185_IOB_X1Y186_I;
  assign RIOI3_X105Y185_ILOGIC_X1Y185_O = RIOB33_X105Y185_IOB_X1Y185_I;
  assign RIOI3_X105Y189_ILOGIC_X1Y190_O = RIOB33_X105Y189_IOB_X1Y190_I;
  assign RIOI3_X105Y189_ILOGIC_X1Y189_O = RIOB33_X105Y189_IOB_X1Y189_I;
  assign RIOI3_X105Y191_ILOGIC_X1Y192_O = RIOB33_X105Y191_IOB_X1Y192_I;
  assign RIOI3_X105Y191_ILOGIC_X1Y191_O = RIOB33_X105Y191_IOB_X1Y191_I;
  assign RIOI3_X105Y195_ILOGIC_X1Y196_O = RIOB33_X105Y195_IOB_X1Y196_I;
  assign RIOI3_X105Y195_ILOGIC_X1Y195_O = RIOB33_X105Y195_IOB_X1Y195_I;
  assign RIOI3_X105Y197_ILOGIC_X1Y198_O = RIOB33_X105Y197_IOB_X1Y198_I;
  assign RIOI3_X105Y197_ILOGIC_X1Y197_O = RIOB33_X105Y197_IOB_X1Y197_I;
  assign RIOI3_X105Y201_ILOGIC_X1Y202_O = RIOB33_X105Y201_IOB_X1Y202_I;
  assign RIOI3_X105Y201_ILOGIC_X1Y201_O = RIOB33_X105Y201_IOB_X1Y201_I;
  assign RIOI3_X105Y203_ILOGIC_X1Y204_O = RIOB33_X105Y203_IOB_X1Y204_I;
  assign RIOI3_X105Y203_ILOGIC_X1Y203_O = RIOB33_X105Y203_IOB_X1Y203_I;
  assign RIOI3_X105Y205_ILOGIC_X1Y205_O = RIOB33_X105Y205_IOB_X1Y205_I;
  assign RIOI3_SING_X105Y50_OLOGIC_X1Y50_OQ = CLBLM_R_X5Y130_SLICE_X7Y130_AQ;
  assign RIOI3_SING_X105Y50_OLOGIC_X1Y50_TQ = 1'b1;
  assign RIOI3_SING_X105Y99_OLOGIC_X1Y99_OQ = CLBLM_R_X7Y126_SLICE_X8Y126_DQ;
  assign RIOI3_SING_X105Y99_OLOGIC_X1Y99_TQ = 1'b1;
  assign RIOI3_SING_X105Y100_OLOGIC_X1Y100_OQ = CLBLL_L_X54Y116_SLICE_X82Y116_AQ;
  assign RIOI3_SING_X105Y100_OLOGIC_X1Y100_TQ = 1'b1;
  assign RIOI3_SING_X105Y149_OLOGIC_X1Y149_OQ = CLBLM_R_X7Y138_SLICE_X9Y138_DQ;
  assign RIOI3_SING_X105Y149_OLOGIC_X1Y149_TQ = 1'b1;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ = CLBLM_R_X7Y129_SLICE_X9Y129_AQ;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ = 1'b1;
  assign RIOI3_SING_X105Y199_ILOGIC_X1Y199_O = RIOB33_SING_X105Y199_IOB_X1Y199_I;
  assign RIOI3_SING_X105Y200_ILOGIC_X1Y200_O = RIOB33_SING_X105Y200_IOB_X1Y200_I;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_OQ = CLBLM_L_X8Y130_SLICE_X10Y130_CQ;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_OQ = CLBLM_R_X7Y137_SLICE_X9Y137_CQ;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_OQ = CLBLM_L_X8Y129_SLICE_X10Y129_CQ;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_OQ = CLBLM_L_X8Y129_SLICE_X10Y129_BQ;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_OQ = CLBLM_L_X8Y130_SLICE_X11Y130_DQ;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_OQ = CLBLM_L_X8Y131_SLICE_X11Y131_CQ;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_OQ = CLBLM_L_X10Y131_SLICE_X13Y131_AQ;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_OQ = CLBLM_L_X12Y132_SLICE_X16Y132_CQ;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_OQ = CLBLM_R_X7Y130_SLICE_X8Y130_BQ;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_OQ = CLBLL_L_X54Y119_SLICE_X82Y119_AQ;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_OQ = CLBLM_L_X10Y133_SLICE_X13Y133_BQ;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_OQ = CLBLM_R_X11Y133_SLICE_X14Y133_AQ;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_OQ = CLBLL_L_X54Y133_SLICE_X82Y133_AQ;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_OQ = CLBLM_R_X5Y134_SLICE_X7Y134_BQ;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_OQ = CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_OQ = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ = CLBLM_L_X8Y130_SLICE_X10Y130_BQ;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ = CLBLM_L_X56Y151_SLICE_X84Y151_AQ;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ = CLBLM_L_X8Y137_SLICE_X10Y137_BQ;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_ILOGIC_X1Y182_O = RIOB33_X105Y181_IOB_X1Y182_I;
  assign RIOI3_TBYTESRC_X105Y181_ILOGIC_X1Y181_O = RIOB33_X105Y181_IOB_X1Y181_I;
  assign RIOI3_TBYTESRC_X105Y193_ILOGIC_X1Y194_O = RIOB33_X105Y193_IOB_X1Y194_I;
  assign RIOI3_TBYTESRC_X105Y193_ILOGIC_X1Y193_O = RIOB33_X105Y193_IOB_X1Y193_I;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_OQ = CLBLL_L_X54Y96_SLICE_X82Y96_AQ;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_OQ = CLBLM_R_X7Y137_SLICE_X9Y137_DQ;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_OQ = CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_OQ = CLBLM_L_X10Y132_SLICE_X12Y132_DQ;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_OQ = CLBLM_R_X7Y131_SLICE_X9Y131_DQ;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_OQ = CLBLM_R_X7Y131_SLICE_X9Y131_CQ;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_OQ = CLBLM_R_X7Y137_SLICE_X8Y137_BQ;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_OQ = CLBLM_R_X5Y137_SLICE_X7Y137_AQ;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ = CLBLM_R_X7Y134_SLICE_X9Y134_AQ;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ = CLBLM_L_X8Y135_SLICE_X10Y135_AQ;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_ILOGIC_X1Y188_O = RIOB33_X105Y187_IOB_X1Y188_I;
  assign RIOI3_TBYTETERM_X105Y187_ILOGIC_X1Y187_O = RIOB33_X105Y187_IOB_X1Y187_I;
  assign RIOB33_SING_X105Y149_IOB_X1Y149_O = CLBLM_R_X7Y138_SLICE_X9Y138_DQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A2 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A3 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A4 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A5 = 1'b1;
  assign RIOB33_X105Y61_IOB_X1Y62_O = CLBLL_L_X4Y134_SLICE_X5Y134_BQ;
  assign RIOB33_X105Y61_IOB_X1Y61_O = CLBLL_L_X4Y135_SLICE_X5Y135_BQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B2 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B3 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B4 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B5 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A1 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A2 = BRAM_L_X6Y140_RAMB18_X0Y56_DO21;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A3 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A4 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A5 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO5;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A6 = CLBLM_R_X5Y132_SLICE_X7Y132_B5Q;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B6 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B1 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO4;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B2 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO5;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B3 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO5;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B4 = CLBLL_L_X4Y133_SLICE_X4Y133_A5Q;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B5 = BRAM_L_X6Y140_RAMB18_X0Y56_DO20;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B6 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO5;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C1 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO4;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C2 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO4;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C3 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO3;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C4 = CLBLM_R_X5Y133_SLICE_X6Y133_BQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C5 = BRAM_L_X6Y140_RAMB18_X0Y56_DO19;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C6 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO4;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_D1 = CLBLM_R_X7Y138_SLICE_X9Y138_AQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D1 = CLBLM_R_X7Y139_SLICE_X9Y139_AO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D2 = CLBLM_R_X5Y132_SLICE_X7Y132_B5Q;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D3 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D4 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D5 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D6 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_T1 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A1 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO7;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A2 = CLBLM_R_X7Y125_SLICE_X9Y125_AQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A3 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A4 = CLBLM_R_X7Y139_SLICE_X8Y139_DO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A5 = BRAM_L_X6Y140_RAMB18_X0Y56_DO23;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A6 = CLBLM_R_X3Y142_SLICE_X2Y142_BQ;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_D1 = CLBLL_L_X54Y138_SLICE_X82Y138_AQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B1 = BRAM_L_X6Y140_RAMB18_X0Y56_DO19;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B2 = CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B3 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO3;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B4 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO4;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B5 = BRAM_L_X6Y140_RAMB18_X0Y56_DO20;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B6 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO4;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_T1 = 1'b1;
  assign RIOB33_SING_X105Y150_IOB_X1Y150_O = CLBLM_R_X7Y129_SLICE_X9Y129_AQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C1 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO2;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C2 = CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C3 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO2;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C4 = BRAM_L_X6Y140_RAMB18_X0Y56_DO18;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C5 = BRAM_L_X6Y140_RAMB18_X0Y56_DO17;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C6 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D1 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D2 = BRAM_L_X6Y140_RAMB18_X0Y56_DO16;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D3 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO0;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D4 = CLBLM_R_X7Y125_SLICE_X9Y125_AQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D5 = BRAM_L_X6Y140_RAMB18_X0Y56_DO17;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D6 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D6 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A1 = CLBLL_L_X4Y131_SLICE_X5Y131_AQ;
  assign LIOI3_X0Y217_ILOGIC_X0Y218_D = LIOB33_X0Y217_IOB_X0Y218_I;
  assign LIOI3_X0Y217_ILOGIC_X0Y217_D = LIOB33_X0Y217_IOB_X0Y217_I;
  assign LIOI3_X0Y95_ILOGIC_X0Y96_D = LIOB33_X0Y95_IOB_X0Y96_I;
  assign LIOI3_X0Y95_ILOGIC_X0Y95_D = LIOB33_X0Y95_IOB_X0Y95_I;
  assign LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y14_D = LIOB33_X0Y13_IOB_X0Y14_I;
  assign LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y13_D = LIOB33_X0Y13_IOB_X0Y13_I;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_WEBWE5 = 1'b0;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A1 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A2 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A3 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A4 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A5 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A6 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B1 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B2 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B3 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B4 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B5 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B6 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C1 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C2 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C3 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C4 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C5 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C6 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D1 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D2 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D3 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D4 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D5 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D6 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A1 = BRAM_L_X6Y140_RAMB18_X0Y56_DO23;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A2 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO7;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A3 = CLBLM_R_X7Y139_SLICE_X9Y139_CO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A4 = CLBLM_R_X3Y149_SLICE_X2Y149_DQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A5 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A6 = CLBLM_R_X5Y133_SLICE_X6Y133_BQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B1 = BRAM_L_X6Y140_RAMB18_X0Y56_DO23;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B2 = CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B3 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B4 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO7;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B5 = CLBLM_R_X7Y139_SLICE_X8Y139_BO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B6 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C1 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C2 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C3 = CLBLM_R_X7Y139_SLICE_X9Y139_BO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C4 = CLBLL_L_X4Y133_SLICE_X4Y133_A5Q;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C5 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C6 = CLBLM_R_X3Y151_SLICE_X3Y151_AQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D1 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D2 = CLBLM_R_X7Y139_SLICE_X8Y139_CO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D3 = CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D4 = CLBLM_R_X3Y145_SLICE_X3Y145_BQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D5 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D6 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_DIADI11 = 1'b0;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_D1 = CLBLM_R_X7Y138_SLICE_X9Y138_CQ;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_T1 = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_D1 = CLBLM_R_X7Y138_SLICE_X9Y138_BQ;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_T1 = 1'b1;
  assign LIOI3_X0Y221_ILOGIC_X0Y222_D = LIOB33_X0Y221_IOB_X0Y222_I;
  assign LIOI3_X0Y221_ILOGIC_X0Y221_D = LIOB33_X0Y221_IOB_X0Y221_I;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_A1 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_A2 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_A3 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_A4 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_A5 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_A6 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_AX = LIOB33_X0Y193_IOB_X0Y194_I;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_B1 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_B2 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_B3 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_B4 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_B5 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_B6 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_BX = LIOB33_X0Y201_IOB_X0Y201_I;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_C1 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_C2 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_C3 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_C4 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_C5 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_C6 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign LIOI3_X0Y97_ILOGIC_X0Y98_D = LIOB33_X0Y97_IOB_X0Y98_I;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOI3_X0Y97_ILOGIC_X0Y97_D = LIOB33_X0Y97_IOB_X0Y97_I;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_CX = LIOB33_X0Y231_IOB_X0Y232_I;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_D1 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_D2 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_D3 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_D4 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_D5 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_D6 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_DX = LIOB33_X0Y243_IOB_X0Y244_I;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_A1 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_A2 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_A3 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_A4 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_A5 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_A6 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_B1 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_B2 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_B3 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_B4 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_B5 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_B6 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_C1 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_C2 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_C3 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_C4 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_C5 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_C6 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_D1 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_D2 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_D3 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_D4 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_D5 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_D6 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X82Y116_A1 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X82Y116_A2 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X82Y116_A3 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X82Y116_A4 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X82Y116_A5 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X82Y116_A6 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X82Y116_AX = CLBLL_L_X4Y135_SLICE_X5Y135_AO5;
  assign CLBLL_L_X54Y116_SLICE_X82Y116_B1 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X82Y116_B2 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X82Y116_B3 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X82Y116_B4 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X82Y116_B5 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X82Y116_B6 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X82Y116_C1 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X82Y116_C2 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X82Y116_C3 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X82Y116_C4 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X82Y116_C5 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X82Y116_C6 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X82Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X54Y116_SLICE_X82Y116_D1 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X82Y116_D2 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X82Y116_D3 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X82Y116_D4 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X82Y116_D5 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X82Y116_D6 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X83Y116_A1 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X83Y116_A2 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X83Y116_A3 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X83Y116_A4 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X83Y116_A5 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X83Y116_A6 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X83Y116_B1 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X83Y116_B2 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X83Y116_B3 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X83Y116_B4 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X83Y116_B5 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X83Y116_B6 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X83Y116_C1 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X83Y116_C2 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X83Y116_C3 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X83Y116_C4 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X83Y116_C5 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X83Y116_C6 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X83Y116_D1 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X83Y116_D2 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X83Y116_D3 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X83Y116_D4 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X83Y116_D5 = 1'b1;
  assign CLBLL_L_X54Y116_SLICE_X83Y116_D6 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_A1 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_A2 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_A3 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_A4 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_A5 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_A6 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_AX = LIOB33_X0Y207_IOB_X0Y207_I;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_B1 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_B2 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_B3 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_B4 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_B5 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_B6 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_BX = LIOB33_X0Y215_IOB_X0Y215_I;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_C1 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_C2 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_C3 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_C4 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_C5 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_C6 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_CX = LIOB33_X0Y215_IOB_X0Y216_I;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_D1 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_D2 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_D3 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_D4 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_D5 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_D6 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_DX = LIOB33_X0Y217_IOB_X0Y217_I;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_A1 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_A2 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_A3 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_A4 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_A5 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_A6 = LIOB33_X0Y237_IOB_X0Y237_I;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_AX = LIOB33_X0Y247_IOB_X0Y247_I;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_B1 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_B2 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_B3 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_B4 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_B5 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_B6 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_BX = LIOB33_X0Y241_IOB_X0Y242_I;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_C1 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_C2 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_C3 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_C4 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_C5 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_C6 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_CX = LIOB33_X0Y245_IOB_X0Y245_I;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_D1 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_D2 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_D3 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_D4 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_D5 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_D6 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_DX = LIOB33_X0Y245_IOB_X0Y246_I;
  assign RIOI3_X105Y145_OLOGIC_X1Y146_D1 = CLBLM_R_X5Y138_SLICE_X7Y138_AQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A3 = 1'b1;
  assign RIOI3_X105Y145_OLOGIC_X1Y146_T1 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A4 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A5 = 1'b1;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_D1 = CLBLM_R_X5Y138_SLICE_X6Y138_BQ;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_T1 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B1 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B2 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B3 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B6 = CLBLM_R_X5Y131_SLICE_X6Y131_A5Q;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C4 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C6 = 1'b1;
  assign LIOI3_X0Y223_ILOGIC_X0Y224_D = LIOB33_X0Y223_IOB_X0Y224_I;
  assign LIOI3_X0Y223_ILOGIC_X0Y223_D = LIOB33_X0Y223_IOB_X0Y223_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_D = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_D = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_D = LIOB33_X0Y63_IOB_X0Y64_I;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A3 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A4 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A5 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B2 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B3 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B4 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B6 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C5 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C6 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_ADDRARDADDR0 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_ADDRARDADDR1 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_ADDRARDADDR2 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_ADDRARDADDR3 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_ADDRARDADDR4 = CLBLM_L_X12Y135_SLICE_X16Y135_AO6;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_ADDRARDADDR5 = CLBLM_R_X15Y135_SLICE_X21Y135_BO6;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_ADDRARDADDR6 = CLBLM_L_X16Y136_SLICE_X22Y136_DO6;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_ADDRARDADDR7 = CLBLM_L_X16Y135_SLICE_X22Y135_DO6;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_ADDRARDADDR8 = CLBLM_L_X16Y135_SLICE_X22Y135_CO6;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_ADDRARDADDR9 = CLBLM_R_X13Y135_SLICE_X18Y135_AO6;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_ADDRARDADDR10 = CLBLM_L_X16Y136_SLICE_X22Y136_CO6;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_ADDRARDADDR11 = CLBLM_L_X16Y136_SLICE_X22Y136_BO6;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_ADDRARDADDR12 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_ADDRARDADDR13 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_ADDRATIEHIGH0 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_ADDRATIEHIGH1 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_ADDRBTIEHIGH0 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_ADDRBTIEHIGH1 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_ADDRBWRADDR0 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_ADDRBWRADDR1 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_ADDRBWRADDR2 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_ADDRBWRADDR3 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_ADDRBWRADDR4 = CLBLM_L_X8Y133_SLICE_X11Y133_DO6;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_ADDRBWRADDR5 = CLBLM_L_X8Y132_SLICE_X10Y132_BO6;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_ADDRBWRADDR6 = CLBLM_L_X10Y134_SLICE_X12Y134_CO6;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_ADDRBWRADDR7 = CLBLM_L_X8Y132_SLICE_X10Y132_AO6;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_ADDRBWRADDR8 = CLBLM_L_X8Y135_SLICE_X11Y135_AO6;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_ADDRBWRADDR9 = CLBLM_L_X8Y134_SLICE_X11Y134_DO6;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_ADDRBWRADDR10 = CLBLM_L_X8Y135_SLICE_X11Y135_CO6;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_ADDRBWRADDR11 = CLBLM_R_X7Y135_SLICE_X9Y135_DO6;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_ADDRBWRADDR12 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_ADDRBWRADDR13 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_RDCLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_WRCLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_DIADI0 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_DIADI1 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_DIADI2 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_DIADI3 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_DIADI4 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_DIADI5 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_DIADI6 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_DIADI7 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_DIADI8 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_DIADI9 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_DIADI10 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_DIADI11 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_DIADI12 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_DIADI13 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_DIADI14 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_DIADI15 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_DIBDI0 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_DIBDI1 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_DIBDI2 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_DIBDI3 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_DIBDI4 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_DIBDI5 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_DIBDI6 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_DIBDI7 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_DIBDI8 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_DIBDI9 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_DIBDI10 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_DIBDI11 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_DIBDI12 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_DIBDI13 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_DIBDI14 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_DIBDI15 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_DIPADIP0 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_DIPADIP1 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_DIPBDIP0 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_DIPBDIP1 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X82Y119_B5 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X82Y119_B6 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X82Y119_C1 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X82Y119_C2 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X82Y119_C3 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X82Y119_C4 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X82Y119_C6 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X82Y119_C5 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X82Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X54Y119_SLICE_X82Y119_D1 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X82Y119_D2 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X82Y119_D3 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X82Y119_D4 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X82Y119_D5 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X82Y119_D6 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_RDEN = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_WREN = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X83Y119_A1 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X83Y119_A2 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X83Y119_A3 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X83Y119_A4 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X83Y119_A5 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X83Y119_A6 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_REGCE = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_REGCEB = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_RDRCLK = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_REGCLKB = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_RST = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_RSTRAMB = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_RSTREG = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_RSTREGB = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_WEA0 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_WEA1 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_WEA2 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_WEA3 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_WEBWE0 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_WEBWE1 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_WEBWE2 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_WEBWE3 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_WEBWE4 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_WEBWE5 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_WEBWE6 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y54_WEBWE7 = 1'b0;
  assign CLBLL_L_X54Y119_SLICE_X83Y119_C1 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X83Y119_C2 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X83Y119_C3 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X83Y119_C4 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X83Y119_C5 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X83Y119_C6 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X83Y119_D1 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X83Y119_D2 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X83Y119_D3 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X83Y119_D4 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X83Y119_D5 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X83Y119_D6 = 1'b1;
  assign RIOI3_X105Y147_OLOGIC_X1Y148_D1 = CLBLM_R_X7Y137_SLICE_X9Y137_BQ;
  assign RIOI3_X105Y147_OLOGIC_X1Y148_T1 = 1'b1;
  assign RIOI3_X105Y147_OLOGIC_X1Y147_D1 = CLBLL_L_X54Y141_SLICE_X82Y141_AQ;
  assign RIOI3_X105Y147_OLOGIC_X1Y147_T1 = 1'b1;
  assign LIOI3_X0Y225_ILOGIC_X0Y226_D = LIOB33_X0Y225_IOB_X0Y226_I;
  assign LIOI3_X0Y225_ILOGIC_X0Y225_D = LIOB33_X0Y225_IOB_X0Y225_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_D = LIOB33_X0Y103_IOB_X0Y103_I;
  assign LIOI3_TBYTETERM_X0Y87_ILOGIC_X0Y88_D = LIOB33_X0Y87_IOB_X0Y88_I;
  assign LIOI3_TBYTETERM_X0Y87_ILOGIC_X0Y87_D = LIOB33_X0Y87_IOB_X0Y87_I;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1 = CLBLM_L_X8Y137_SLICE_X10Y137_BQ;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1 = 1'b1;
  assign RIOI3_SING_X105Y50_OLOGIC_X1Y50_D1 = CLBLM_R_X5Y130_SLICE_X7Y130_AQ;
  assign RIOI3_SING_X105Y50_OLOGIC_X1Y50_T1 = 1'b1;
  assign RIOB33_X105Y113_IOB_X1Y114_O = CLBLM_R_X7Y131_SLICE_X9Y131_DQ;
  assign RIOB33_X105Y113_IOB_X1Y113_O = CLBLM_R_X7Y131_SLICE_X9Y131_CQ;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_D1 = CLBLM_R_X7Y129_SLICE_X9Y129_BQ;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_D1 = CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_T1 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A2 = BRAM_R_X17Y135_RAMB18_X1Y54_DO3;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A3 = BRAM_R_X17Y135_RAMB18_X1Y54_DO4;
  assign LIOI3_X0Y227_ILOGIC_X0Y228_D = LIOB33_X0Y227_IOB_X0Y228_I;
  assign LIOI3_X0Y227_ILOGIC_X0Y227_D = LIOB33_X0Y227_IOB_X0Y227_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A1 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A2 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A3 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A4 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A5 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A6 = 1'b1;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_D = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_D = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B1 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B2 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B3 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B4 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B5 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B6 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C1 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C2 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C3 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C4 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C5 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C6 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C6 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D1 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D2 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D3 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D4 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D5 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D = LIOB33_X0Y113_IOB_X0Y114_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A1 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A2 = CLBLM_R_X3Y129_SLICE_X2Y129_BQ;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A3 = CLBLM_R_X3Y129_SLICE_X2Y129_AQ;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A4 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A5 = CLBLM_R_X3Y129_SLICE_X2Y129_A5Q;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A6 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X82Y123_A1 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X82Y123_A2 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X82Y123_A3 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X82Y123_A4 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X82Y123_A5 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X82Y123_A6 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B1 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X82Y123_AX = CLBLM_R_X5Y134_SLICE_X6Y134_AO5;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B2 = CLBLM_R_X3Y129_SLICE_X2Y129_BQ;
  assign CLBLL_L_X54Y123_SLICE_X82Y123_B1 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X82Y123_B2 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X82Y123_B3 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X82Y123_B4 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X82Y123_B5 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X82Y123_B6 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B4 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B5 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X82Y123_C1 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X82Y123_C2 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X82Y123_C3 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X82Y123_C4 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X82Y123_C5 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X82Y123_C6 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C3 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C4 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X82Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_ADDRARDADDR0 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_ADDRARDADDR1 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_ADDRARDADDR2 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_ADDRARDADDR3 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_ADDRARDADDR4 = CLBLM_L_X10Y136_SLICE_X13Y136_DO6;
  assign CLBLL_L_X54Y123_SLICE_X82Y123_D1 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X82Y123_D2 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X82Y123_D3 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X82Y123_D4 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X82Y123_D5 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X82Y123_D6 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_ADDRARDADDR5 = CLBLM_R_X11Y135_SLICE_X14Y135_BO6;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_ADDRARDADDR6 = CLBLM_L_X12Y135_SLICE_X16Y135_BO6;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_ADDRARDADDR7 = CLBLM_L_X10Y134_SLICE_X12Y134_BO6;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_ADDRARDADDR8 = CLBLM_L_X10Y136_SLICE_X12Y136_CO6;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_ADDRARDADDR9 = CLBLM_R_X11Y135_SLICE_X14Y135_CO6;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_ADDRARDADDR10 = CLBLM_R_X11Y136_SLICE_X14Y136_DO6;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_ADDRARDADDR11 = CLBLM_R_X13Y136_SLICE_X18Y136_BO6;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_ADDRARDADDR12 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_ADDRARDADDR13 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_ADDRATIEHIGH0 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_ADDRATIEHIGH1 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_ADDRBTIEHIGH0 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_ADDRBTIEHIGH1 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_ADDRBWRADDR0 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_ADDRBWRADDR1 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_ADDRBWRADDR2 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_ADDRBWRADDR3 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_ADDRBWRADDR4 = CLBLM_L_X8Y133_SLICE_X11Y133_CO6;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_ADDRBWRADDR5 = CLBLM_L_X8Y134_SLICE_X11Y134_BO6;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_ADDRBWRADDR6 = CLBLM_L_X8Y135_SLICE_X10Y135_DO6;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_ADDRBWRADDR7 = CLBLM_L_X8Y133_SLICE_X10Y133_BO6;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_ADDRBWRADDR8 = CLBLM_L_X8Y133_SLICE_X10Y133_AO6;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_CLKBWRCLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_ADDRBWRADDR9 = CLBLM_L_X8Y135_SLICE_X11Y135_DO6;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_ADDRBWRADDR10 = CLBLM_L_X8Y135_SLICE_X10Y135_CO6;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_ADDRBWRADDR11 = CLBLM_R_X7Y136_SLICE_X9Y136_CO6;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_ADDRBWRADDR12 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_ADDRBWRADDR13 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_CLKARDCLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_DIADI6 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X83Y123_A1 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X83Y123_A2 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X83Y123_A3 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X83Y123_A4 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X83Y123_A5 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X83Y123_A6 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_DIADI14 = 1'b0;
  assign CLBLL_L_X54Y123_SLICE_X83Y123_B1 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X83Y123_B2 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_DIBDI1 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_DIBDI2 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_DIBDI3 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_DIBDI4 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_DIBDI5 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X83Y123_B3 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X83Y123_B4 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X83Y123_B5 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X83Y123_B6 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X83Y123_C2 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X83Y123_C3 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X83Y123_C4 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X83Y123_C5 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X83Y123_C6 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_DIBDI7 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_DIBDI8 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_DIBDI9 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_DIBDI10 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_DIBDI11 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_DIBDI12 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_DIBDI13 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_DIBDI14 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_DIBDI15 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_DIPADIP0 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_DIPADIP1 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_DIPBDIP0 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_DIPBDIP1 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X83Y123_D1 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X83Y123_D2 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X83Y123_D3 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X83Y123_D4 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X83Y123_D5 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X83Y123_D6 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_C4 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_ENARDEN = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_ENBWREN = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B1 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO7;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_REGCEAREGCE = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_REGCEB = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_REGCLKARDRCLK = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_REGCLKB = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_RSTRAMARSTRAM = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_RSTRAMB = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_RSTREGARSTREG = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_RSTREGB = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_WEA0 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_WEA1 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_WEA2 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_WEA3 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_WEBWE0 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_WEBWE1 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_WEBWE2 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_WEBWE3 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_WEBWE4 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_WEBWE5 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_WEBWE6 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_WEBWE7 = 1'b0;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B4 = CLBLM_R_X7Y134_SLICE_X9Y134_B5Q;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C2 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C3 = CLBLM_R_X3Y155_SLICE_X2Y155_DQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C4 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C5 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A1 = CLBLM_R_X7Y131_SLICE_X9Y131_A5Q;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A2 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A3 = CLBLM_R_X3Y130_SLICE_X3Y130_AQ;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A4 = BRAM_L_X6Y125_RAMB18_X0Y50_DO21;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A6 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B1 = LIOB33_X0Y27_IOB_X0Y27_I;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B2 = CLBLM_R_X3Y130_SLICE_X3Y130_BQ;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B3 = CLBLM_R_X3Y130_SLICE_X3Y130_AQ;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B5 = BRAM_L_X6Y125_RAMB18_X0Y50_DO21;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B6 = CLBLM_R_X7Y131_SLICE_X9Y131_A5Q;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C1 = CLBLM_R_X3Y130_SLICE_X2Y130_AQ;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C2 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C3 = CLBLM_R_X3Y131_SLICE_X2Y131_DO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C5 = CLBLM_R_X5Y130_SLICE_X7Y130_BQ;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C6 = CLBLM_R_X3Y131_SLICE_X3Y131_BQ;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D1 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D2 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D3 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D4 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D5 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D6 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A1 = CLBLM_R_X3Y131_SLICE_X2Y131_DO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A2 = CLBLM_R_X3Y131_SLICE_X3Y131_BQ;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A3 = CLBLM_R_X3Y130_SLICE_X2Y130_AQ;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A5 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A6 = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B1 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B2 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B3 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B4 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B5 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B6 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_B4 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C1 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C2 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C3 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C4 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C5 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_B5 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C6 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D1 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D2 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D3 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D4 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D5 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D6 = 1'b1;
  assign RIOI3_SING_X105Y100_OLOGIC_X1Y100_D1 = CLBLL_L_X54Y116_SLICE_X82Y116_AQ;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_C3 = 1'b1;
  assign RIOI3_SING_X105Y100_OLOGIC_X1Y100_T1 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_C4 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_C6 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_D1 = CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_T1 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_D1 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_T1 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A1 = CLBLM_R_X3Y131_SLICE_X3Y131_B5Q;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A2 = BRAM_L_X6Y130_RAMB18_X0Y52_DO18;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A3 = LIOB33_X0Y141_IOB_X0Y142_I;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A4 = CLBLM_R_X3Y131_SLICE_X2Y131_BQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A5 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A6 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_AX = CLBLM_R_X3Y131_SLICE_X2Y131_DO5;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B1 = LIOB33_X0Y87_IOB_X0Y88_I;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B2 = CLBLM_R_X3Y131_SLICE_X3Y131_BQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B3 = CLBLM_R_X3Y131_SLICE_X3Y131_AQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B5 = BRAM_L_X6Y130_RAMB18_X0Y52_DO16;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B6 = CLBLL_L_X2Y131_SLICE_X1Y131_BQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_BX = CLBLM_R_X3Y131_SLICE_X3Y131_AO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C1 = BRAM_L_X6Y130_RAMB18_X0Y52_DO18;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C2 = CLBLM_R_X3Y131_SLICE_X3Y131_CQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C3 = LIOB33_X0Y89_IOB_X0Y90_I;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C5 = CLBLM_R_X3Y131_SLICE_X3Y131_B5Q;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C6 = CLBLM_R_X3Y131_SLICE_X2Y131_BQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D1 = CLBLM_R_X3Y132_SLICE_X3Y132_AQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D2 = CLBLM_R_X3Y131_SLICE_X2Y131_A5Q;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D3 = CLBLM_R_X3Y131_SLICE_X3Y131_DQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D4 = BRAM_L_X6Y130_RAMB18_X0Y52_DO20;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D5 = LIOB33_X0Y91_IOB_X0Y92_I;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D6 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A1 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A2 = CLBLL_L_X2Y131_SLICE_X1Y131_A5Q;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A3 = CLBLM_R_X3Y129_SLICE_X2Y129_A5Q;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A4 = CLBLM_R_X3Y129_SLICE_X2Y129_BQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A5 = CLBLM_R_X3Y129_SLICE_X2Y129_AQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A6 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B1 = CLBLL_L_X2Y131_SLICE_X1Y131_A5Q;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B2 = CLBLM_R_X3Y129_SLICE_X2Y129_BQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B3 = CLBLM_R_X3Y129_SLICE_X2Y129_AQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B4 = CLBLM_R_X3Y129_SLICE_X2Y129_A5Q;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B5 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B6 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C1 = CLBLM_R_X3Y129_SLICE_X2Y129_AQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C2 = CLBLM_R_X3Y129_SLICE_X2Y129_BQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C3 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C4 = CLBLM_R_X3Y129_SLICE_X2Y129_A5Q;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C5 = CLBLL_L_X2Y131_SLICE_X1Y131_A5Q;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C6 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y229_ILOGIC_X0Y230_D = LIOB33_X0Y229_IOB_X0Y230_I;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D1 = CLBLM_R_X3Y131_SLICE_X3Y131_AQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D2 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D3 = BRAM_L_X6Y130_RAMB18_X0Y52_DO16;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D4 = CLBLL_L_X2Y131_SLICE_X1Y131_BQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D5 = LIOB33_X0Y139_IOB_X0Y140_I;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D6 = 1'b1;
  assign LIOI3_X0Y229_ILOGIC_X0Y229_D = LIOB33_X0Y229_IOB_X0Y229_I;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_SR = LIOB33_X0Y147_IOB_X0Y148_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_D = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_D = LIOB33_X0Y109_IOB_X0Y109_I;
  assign LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y138_D = LIOB33_X0Y137_IOB_X0Y138_I;
  assign LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_D = LIOB33_X0Y137_IOB_X0Y137_I;
  assign RIOI3_SING_X105Y149_OLOGIC_X1Y149_D1 = CLBLM_R_X7Y138_SLICE_X9Y138_DQ;
  assign RIOI3_SING_X105Y149_OLOGIC_X1Y149_T1 = 1'b1;
  assign LIOI3_SING_X0Y249_ILOGIC_X0Y249_D = LIOB33_SING_X0Y249_IOB_X0Y249_I;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A1 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A2 = BRAM_L_X6Y130_RAMB18_X0Y52_DO20;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A3 = CLBLM_R_X3Y132_SLICE_X3Y132_AQ;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A5 = CLBLM_R_X3Y131_SLICE_X2Y131_A5Q;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A6 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B1 = LIOB33_X0Y93_IOB_X0Y93_I;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B2 = CLBLM_R_X3Y132_SLICE_X3Y132_BQ;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B3 = CLBLL_L_X2Y131_SLICE_X1Y131_AQ;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B5 = CLBLM_R_X3Y133_SLICE_X3Y133_AQ;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B6 = BRAM_L_X6Y130_RAMB18_X0Y52_DO21;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C1 = CLBLM_R_X3Y132_SLICE_X2Y132_DQ;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C2 = CLBLM_R_X3Y132_SLICE_X3Y132_CQ;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C3 = CLBLM_R_X3Y132_SLICE_X2Y132_BO5;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C4 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C5 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C6 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D1 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D2 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D3 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D4 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D5 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D6 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A1 = BRAM_L_X6Y130_RAMB18_X0Y52_DO22;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A2 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A3 = CLBLM_R_X3Y132_SLICE_X2Y132_AQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A4 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A5 = CLBLM_R_X3Y131_SLICE_X2Y131_CQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A6 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B1 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B2 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B3 = CLBLM_R_X3Y131_SLICE_X2Y131_C5Q;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B4 = BRAM_L_X6Y130_RAMB18_X0Y52_DO23;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B5 = CLBLM_R_X3Y132_SLICE_X2Y132_BQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B6 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C1 = CLBLM_R_X3Y132_SLICE_X2Y132_AQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C2 = CLBLM_R_X3Y132_SLICE_X2Y132_CQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C3 = BRAM_L_X6Y130_RAMB18_X0Y52_DO22;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C4 = CLBLM_R_X3Y131_SLICE_X2Y131_CQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C5 = LIOB33_X0Y93_IOB_X0Y94_I;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C6 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D1 = CLBLM_R_X3Y132_SLICE_X2Y132_BQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D2 = CLBLM_R_X3Y131_SLICE_X2Y131_C5Q;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D3 = CLBLM_R_X3Y132_SLICE_X2Y132_DQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D4 = BRAM_L_X6Y130_RAMB18_X0Y52_DO23;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D5 = LIOB33_X0Y95_IOB_X0Y95_I;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D6 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0 = LIOB33_X0Y127_IOB_X0Y128_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1 = CLBLM_R_X7Y129_SLICE_X9Y129_AQ;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A1 = LIOB33_X0Y145_IOB_X0Y145_I;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A2 = BRAM_L_X6Y130_RAMB18_X0Y52_DO21;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A3 = CLBLM_R_X3Y133_SLICE_X3Y133_AQ;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A5 = CLBLL_L_X2Y131_SLICE_X1Y131_AQ;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A6 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B1 = CLBLM_R_X3Y131_SLICE_X3Y131_DQ;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B2 = CLBLM_R_X3Y133_SLICE_X3Y133_BQ;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B3 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B5 = CLBLM_R_X3Y132_SLICE_X3Y132_AO5;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B6 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C1 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C2 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C3 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C4 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C5 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C6 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D1 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D2 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D3 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D4 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D5 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D6 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_D1 = CLBLM_R_X7Y129_SLICE_X8Y129_BQ;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A1 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A2 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A3 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A4 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A5 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A6 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_T1 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B1 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B2 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B3 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B4 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B5 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B6 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_D1 = CLBLM_R_X7Y136_SLICE_X8Y136_AQ;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C1 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C2 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C3 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C4 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C5 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C6 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_T1 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D1 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D2 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D3 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D4 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D5 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D6 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign LIOI3_X0Y233_ILOGIC_X0Y234_D = LIOB33_X0Y233_IOB_X0Y234_I;
  assign LIOI3_X0Y233_ILOGIC_X0Y233_D = LIOB33_X0Y233_IOB_X0Y233_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_D = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_D = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A1 = CLBLM_R_X3Y132_SLICE_X3Y132_AQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A2 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO3;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A3 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO4;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A5 = BRAM_R_X17Y135_RAMB18_X1Y54_DO3;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A6 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO4;
  assign LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y164_D = LIOB33_X0Y163_IOB_X0Y164_I;
  assign LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y163_D = LIOB33_X0Y163_IOB_X0Y163_I;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_A1 = LIOB33_X0Y13_IOB_X0Y14_I;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_A2 = CLBLL_L_X4Y134_SLICE_X4Y134_AQ;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_A3 = CLBLM_R_X3Y134_SLICE_X2Y134_AO5;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_A4 = CLBLM_R_X3Y134_SLICE_X2Y134_BQ;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_A5 = BRAM_L_X6Y125_RAMB18_X0Y50_DO23;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_A6 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_B1 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_B2 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_B3 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_B4 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_B5 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_B6 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_C1 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_C2 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_C3 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_C4 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_C5 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_C6 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_D1 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_D2 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_D3 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_D4 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_D5 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_D6 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C5 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO2;
  assign RIOI3_SING_X105Y199_ILOGIC_X1Y199_D = RIOB33_SING_X105Y199_IOB_X1Y199_I;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C6 = CLBLM_R_X7Y134_SLICE_X9Y134_A5Q;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_A1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_A2 = CLBLM_R_X5Y134_SLICE_X7Y134_A5Q;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_A3 = CLBLM_R_X3Y134_SLICE_X2Y134_AQ;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_A4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_A5 = BRAM_L_X6Y125_RAMB18_X0Y50_DO23;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_A6 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_B1 = CLBLM_R_X5Y134_SLICE_X7Y134_A5Q;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_B2 = CLBLM_R_X3Y134_SLICE_X2Y134_BQ;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_B3 = CLBLM_R_X3Y134_SLICE_X2Y134_AQ;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_B4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_B5 = BRAM_L_X6Y125_RAMB18_X0Y50_DO23;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_B6 = LIOB33_X0Y29_IOB_X0Y29_I;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_C1 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_C2 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_C3 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_C4 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_C5 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_C6 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_D1 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_D2 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_D3 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_D4 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_D5 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_D6 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B2 = BRAM_L_X6Y135_RAMB18_X0Y54_DO7;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D1 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO0;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D2 = BRAM_L_X6Y135_RAMB18_X0Y54_DO1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D4 = CLBLM_L_X8Y135_SLICE_X10Y135_A5Q;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D5 = BRAM_R_X17Y135_RAMB18_X1Y54_DO1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A1 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A2 = LIOB33_X0Y137_IOB_X0Y137_I;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A4 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO5;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A5 = CLBLM_L_X10Y135_SLICE_X12Y135_A5Q;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A6 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_A5 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_C5 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_A6 = CLBLL_L_X2Y142_SLICE_X0Y142_CQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B5 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO5;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A3 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A4 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_B4 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_B5 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_B6 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_A1 = CLBLM_R_X5Y135_SLICE_X6Y135_BO6;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_A2 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_A3 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_A4 = CLBLM_R_X5Y132_SLICE_X7Y132_A5Q;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_A5 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_A6 = CLBLM_R_X3Y147_SLICE_X2Y147_CQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_B1 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_B2 = CLBLM_R_X5Y135_SLICE_X7Y135_BO6;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_B3 = CLBLL_L_X2Y158_SLICE_X0Y158_BQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_B4 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_B5 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_B6 = CLBLL_L_X4Y131_SLICE_X5Y131_B5Q;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_C1 = CLBLM_R_X3Y134_SLICE_X2Y134_AQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_C2 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_C3 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_C4 = CLBLL_L_X2Y158_SLICE_X0Y158_CQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_C5 = CLBLM_R_X5Y135_SLICE_X6Y135_CO6;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_C6 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_D1 = CLBLM_R_X5Y130_SLICE_X6Y130_B5Q;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_D2 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_D3 = CLBLM_R_X5Y135_SLICE_X6Y135_DO6;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_D4 = CLBLM_R_X3Y147_SLICE_X3Y147_CQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_D5 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_D6 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_A1 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_A2 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_A3 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_A4 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_A5 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_A6 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_B1 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_B2 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_B3 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_B4 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_B5 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_B6 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_C1 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_C2 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_C3 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_C4 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_C5 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_C6 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_D1 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_D2 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_D3 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_D4 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_D5 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_D6 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D1 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A1 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A2 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A3 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A4 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A5 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A6 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D2 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B1 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B2 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B3 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B4 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B5 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B6 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C1 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C2 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C3 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C4 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C5 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C6 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D1 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D2 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D3 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D4 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D5 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D6 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_C4 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_C5 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A1 = BRAM_R_X17Y135_RAMB18_X1Y54_DO19;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A2 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A3 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A4 = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A5 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A6 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_C6 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B1 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B2 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B3 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B4 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B5 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B6 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_D1 = CLBLM_R_X7Y137_SLICE_X8Y137_AQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C1 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C2 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C3 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C4 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C5 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C6 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_T1 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A5 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_D1 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D1 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D2 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D3 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D4 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D5 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D6 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A6 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_T1 = 1'b1;
  assign RIOI3_X105Y125_OLOGIC_X1Y126_D1 = CLBLM_R_X7Y130_SLICE_X9Y130_CQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_BX = LIOB33_X0Y171_IOB_X0Y171_I;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C1 = 1'b1;
  assign RIOI3_X105Y197_ILOGIC_X1Y198_D = RIOB33_X105Y197_IOB_X1Y198_I;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C6 = 1'b1;
  assign RIOI3_X105Y197_ILOGIC_X1Y197_D = RIOB33_X105Y197_IOB_X1Y197_I;
  assign LIOI3_X0Y235_ILOGIC_X0Y236_D = LIOB33_X0Y235_IOB_X0Y236_I;
  assign LIOI3_X0Y235_ILOGIC_X0Y235_D = LIOB33_X0Y235_IOB_X0Y235_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_D = LIOB33_X0Y115_IOB_X0Y116_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_D = LIOB33_X0Y115_IOB_X0Y115_I;
  assign LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y188_D = LIOB33_X0Y187_IOB_X0Y188_I;
  assign LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y187_D = LIOB33_X0Y187_IOB_X0Y187_I;
  assign RIOI3_SING_X105Y99_OLOGIC_X1Y99_D1 = CLBLM_R_X7Y126_SLICE_X8Y126_DQ;
  assign RIOI3_SING_X105Y99_OLOGIC_X1Y99_T1 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_A1 = CLBLL_L_X4Y132_SLICE_X4Y132_AQ;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_A2 = BRAM_R_X17Y135_RAMB18_X1Y54_DO1;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_A3 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_A4 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_A5 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_A6 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_B1 = CLBLL_L_X4Y132_SLICE_X4Y132_AQ;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_B2 = BRAM_R_X17Y135_RAMB18_X1Y54_DO7;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_B3 = CLBLM_L_X10Y135_SLICE_X13Y135_BO6;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_B4 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO7;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_B5 = CLBLM_R_X25Y157_SLICE_X36Y157_AQ;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_B6 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_C1 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_C2 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_C3 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_C4 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_C5 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_C6 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_D1 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_D2 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_D3 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_D4 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_D5 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_D6 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_A1 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_A2 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_A3 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_A4 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_A5 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_A6 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_B1 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_B2 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_B3 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_B4 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_B5 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_B6 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_C1 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_C2 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_C3 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_C4 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_C5 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_C6 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_D1 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_D2 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_D3 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_D4 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_D5 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_D6 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_A1 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_A2 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO7;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_A3 = CLBLM_R_X3Y134_SLICE_X2Y134_BQ;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_A4 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO7;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_A5 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_A6 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_B1 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO7;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_B2 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO6;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_B3 = CLBLL_L_X4Y133_SLICE_X5Y133_BQ;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_B4 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO7;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_B5 = BRAM_L_X6Y140_RAMB18_X0Y56_DO7;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_B6 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO6;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_C1 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO6;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_C2 = BRAM_L_X6Y140_RAMB18_X0Y56_DO7;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_C3 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO7;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_C4 = BRAM_L_X6Y140_RAMB18_X0Y56_DO6;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_C5 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO7;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_C6 = CLBLL_L_X4Y128_SLICE_X5Y128_BQ;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_D1 = CLBLM_R_X3Y157_SLICE_X3Y157_AQ;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_D2 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_D3 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_D4 = CLBLL_L_X4Y133_SLICE_X5Y133_BQ;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_D5 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_D6 = CLBLM_R_X3Y137_SLICE_X3Y137_BO6;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_A1 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO7;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_A2 = CLBLM_R_X3Y130_SLICE_X2Y130_AQ;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_A3 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO0;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_A4 = BRAM_L_X6Y140_RAMB18_X0Y56_DO7;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_A5 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO0;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_A6 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO0;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_B1 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO7;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_B2 = BRAM_L_X6Y140_RAMB18_X0Y56_DO7;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_B3 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO6;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_B4 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO7;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_B5 = CLBLM_R_X3Y134_SLICE_X2Y134_BQ;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_B6 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO6;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_C1 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_C2 = CLBLL_L_X2Y155_SLICE_X0Y155_BQ;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_C3 = CLBLL_L_X4Y137_SLICE_X4Y137_BO6;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_C4 = CLBLL_L_X4Y131_SLICE_X4Y131_DQ;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_C5 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_C6 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_D1 = CLBLM_R_X3Y134_SLICE_X2Y134_BQ;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_D2 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_D3 = CLBLL_L_X2Y155_SLICE_X1Y155_BQ;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_D4 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_D5 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_D6 = CLBLM_R_X3Y137_SLICE_X2Y137_BO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A1 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A2 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A3 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A4 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A5 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A6 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B1 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B2 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B3 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B4 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B5 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B6 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C1 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C2 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C3 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C4 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C5 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C6 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D1 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D2 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D3 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D4 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D5 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D6 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A1 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A2 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A3 = CLBLM_R_X7Y130_SLICE_X8Y130_B5Q;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A4 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A5 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A6 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B1 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B2 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B3 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B4 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO7;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B5 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B6 = CLBLL_L_X4Y132_SLICE_X5Y132_A5Q;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C1 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C2 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C3 = CLBLM_R_X3Y132_SLICE_X3Y132_BQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C4 = BRAM_R_X17Y135_RAMB18_X1Y54_DO21;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C5 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C6 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D1 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D2 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D3 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D4 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D5 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D6 = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_D1 = CLBLM_L_X8Y132_SLICE_X11Y132_AQ;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_T1 = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_D1 = CLBLM_R_X5Y134_SLICE_X7Y134_AQ;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_T1 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_A1 = BRAM_L_X6Y140_RAMB18_X0Y56_DO7;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_A2 = CLBLM_R_X3Y133_SLICE_X3Y133_BQ;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_A3 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO7;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_A4 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_A5 = CLBLL_L_X2Y157_SLICE_X0Y157_AQ;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_A6 = CLBLL_L_X4Y138_SLICE_X5Y138_BO6;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_B1 = BRAM_L_X6Y140_RAMB18_X0Y56_DO7;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_B2 = CLBLL_L_X4Y138_SLICE_X4Y138_CO6;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_B3 = CLBLM_R_X5Y126_SLICE_X6Y126_BQ;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_B4 = CLBLM_R_X3Y153_SLICE_X3Y153_AQ;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_B5 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_B6 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO7;
  assign CLBLM_R_X25Y157_SLICE_X37Y157_A1 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_C1 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_C2 = BRAM_L_X6Y140_RAMB18_X0Y56_DO7;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_C3 = CLBLM_R_X3Y151_SLICE_X2Y151_CQ;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_C4 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO7;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_C5 = CLBLL_L_X4Y137_SLICE_X4Y137_DO6;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_C6 = CLBLM_R_X5Y125_SLICE_X7Y125_CQ;
  assign CLBLM_R_X25Y157_SLICE_X37Y157_A2 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X37Y157_A3 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X37Y157_A4 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_D1 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_D2 = CLBLL_L_X4Y128_SLICE_X5Y128_BQ;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_D3 = CLBLM_R_X3Y153_SLICE_X3Y153_DQ;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_D4 = CLBLM_R_X3Y137_SLICE_X3Y137_CO6;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_D5 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_D6 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_A1 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_A2 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_A3 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_A4 = CLBLL_L_X2Y132_SLICE_X1Y132_AQ;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_A5 = CLBLL_L_X4Y136_SLICE_X4Y136_AO6;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_A6 = CLBLL_L_X2Y157_SLICE_X0Y157_CQ;
  assign CLBLM_R_X25Y157_SLICE_X37Y157_AX = RIOB33_X105Y205_IOB_X1Y205_I;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_B1 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_B2 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_B3 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_B4 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_B5 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_B6 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_C1 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_C2 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_C3 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_C4 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_C5 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_C6 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_D1 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_D2 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_D3 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_D4 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_D5 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_D6 = 1'b1;
  assign LIOI3_X0Y239_ILOGIC_X0Y240_D = LIOB33_X0Y239_IOB_X0Y240_I;
  assign LIOI3_X0Y239_ILOGIC_X0Y239_D = LIOB33_X0Y239_IOB_X0Y239_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y118_D = LIOB33_X0Y117_IOB_X0Y118_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_D = LIOB33_X0Y117_IOB_X0Y117_I;
  assign LIOI3_TBYTETERM_X0Y213_ILOGIC_X0Y214_D = LIOB33_X0Y213_IOB_X0Y214_I;
  assign LIOI3_TBYTETERM_X0Y213_ILOGIC_X0Y213_D = LIOB33_X0Y213_IOB_X0Y213_I;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_A1 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_A2 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_A3 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_A4 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_A5 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X82Y133_A1 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X82Y133_A2 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X82Y133_A3 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X82Y133_A4 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X82Y133_A5 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X82Y133_A6 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_A6 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X82Y133_AX = CLBLL_L_X4Y135_SLICE_X4Y135_AO5;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_B1 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X82Y133_B1 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X82Y133_B2 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X82Y133_B3 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X82Y133_B4 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X82Y133_B5 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X82Y133_B6 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_B3 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_B4 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_B6 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X82Y133_C1 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X82Y133_C2 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X82Y133_C3 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X82Y133_C4 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X82Y133_C5 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X82Y133_C6 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_C3 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_C4 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X82Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_C6 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_D1 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_D2 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_D3 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X82Y133_D1 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X82Y133_D2 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X82Y133_D3 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X82Y133_D4 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X82Y133_D5 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X82Y133_D6 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_D4 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_D5 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_A1 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_A2 = CLBLM_R_X3Y130_SLICE_X2Y130_AQ;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_A3 = CLBLM_R_X3Y137_SLICE_X2Y137_AO6;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_A4 = CLBLM_R_X3Y157_SLICE_X3Y157_BQ;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_A5 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_A6 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_B1 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_B2 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_B3 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_B4 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_B5 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_B6 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_C1 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_C2 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_C3 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_C4 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_C5 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X83Y133_A1 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X83Y133_A2 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X83Y133_A3 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X83Y133_A4 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X83Y133_A5 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X83Y133_A6 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_C6 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X83Y133_B1 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X83Y133_B2 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X83Y133_B3 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X83Y133_B4 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X83Y133_B5 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X83Y133_B6 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_D1 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_D2 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_D3 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X83Y133_C1 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X83Y133_C2 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X83Y133_C3 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X83Y133_C4 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X83Y133_C5 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X83Y133_C6 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D2 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLL_L_X54Y133_SLICE_X83Y133_D1 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X83Y133_D2 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X83Y133_D3 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X83Y133_D4 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X83Y133_D5 = 1'b1;
  assign CLBLL_L_X54Y133_SLICE_X83Y133_D6 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D4 = CLBLM_L_X8Y132_SLICE_X11Y132_A5Q;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_B3 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_C1 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_C2 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_D1 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_D1 = CLBLM_L_X8Y136_SLICE_X10Y136_AQ;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_B1 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_T1 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_B3 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_B4 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_D1 = CLBLM_R_X7Y134_SLICE_X9Y134_BQ;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A1 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A2 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_B5 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A4 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A3 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A6 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A5 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B1 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B2 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B3 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B4 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B5 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B6 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_T1 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C1 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C2 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C3 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C4 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C5 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C6 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D1 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D2 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D3 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D4 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D5 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D6 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A1 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A2 = CLBLM_R_X25Y154_SLICE_X36Y154_AQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A3 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A4 = CLBLM_R_X3Y131_SLICE_X3Y131_AQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A5 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A6 = CLBLM_R_X11Y135_SLICE_X14Y135_AO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B1 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B2 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B3 = CLBLM_L_X16Y152_SLICE_X22Y152_BQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B4 = CLBLM_R_X7Y134_SLICE_X9Y134_A5Q;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B5 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B6 = CLBLM_L_X10Y135_SLICE_X13Y135_CO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C1 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C2 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C3 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C4 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C5 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C6 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D1 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D2 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D3 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D4 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D5 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D6 = 1'b1;
  assign LIOI3_X0Y241_ILOGIC_X0Y242_D = LIOB33_X0Y241_IOB_X0Y242_I;
  assign LIOI3_X0Y241_ILOGIC_X0Y241_D = LIOB33_X0Y241_IOB_X0Y241_I;
  assign LIOI3_X0Y121_ILOGIC_X0Y122_D = LIOB33_X0Y121_IOB_X0Y122_I;
  assign LIOI3_X0Y121_ILOGIC_X0Y121_D = LIOB33_X0Y121_IOB_X0Y121_I;
  assign LIOI3_TBYTETERM_X0Y237_ILOGIC_X0Y238_D = LIOB33_X0Y237_IOB_X0Y238_I;
  assign LIOI3_TBYTETERM_X0Y237_ILOGIC_X0Y237_D = LIOB33_X0Y237_IOB_X0Y237_I;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A1 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A2 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A3 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A4 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A5 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A6 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B1 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B2 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B3 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B4 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B5 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B6 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C1 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C2 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C3 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C4 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C5 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C6 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D1 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D2 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D3 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D4 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D5 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D6 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A1 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A2 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A3 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A4 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A5 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A6 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_AX = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B1 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B2 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B3 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B4 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B5 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B6 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_BX = LIOB33_X0Y159_IOB_X0Y160_I;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C1 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C2 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C3 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C4 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C5 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C6 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_CX = LIOB33_X0Y157_IOB_X0Y158_I;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D1 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D2 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D3 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D4 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D5 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D6 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A1 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A2 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A3 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A4 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A5 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A6 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B1 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B2 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B3 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B4 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B5 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B6 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C1 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C2 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C3 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C4 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C5 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C6 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D1 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D2 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D3 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D4 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D5 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D6 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A1 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A2 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A3 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A4 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A5 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A6 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_AX = LIOB33_X0Y161_IOB_X0Y161_I;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B1 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B2 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B3 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B4 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B5 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B6 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_BX = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C1 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C2 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C3 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C4 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C5 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C6 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_CX = LIOB33_X0Y153_IOB_X0Y153_I;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D1 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D2 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D3 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D4 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D5 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D6 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_DX = LIOB33_X0Y159_IOB_X0Y159_I;
  assign RIOB33_X105Y51_IOB_X1Y52_O = CLBLM_R_X5Y134_SLICE_X7Y134_CQ;
  assign RIOB33_X105Y51_IOB_X1Y51_O = CLBLM_R_X5Y132_SLICE_X7Y132_BQ;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_D1 = CLBLM_L_X8Y137_SLICE_X10Y137_AQ;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_T1 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_D1 = CLBLM_L_X10Y135_SLICE_X12Y135_AQ;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_T1 = 1'b1;
  assign LIOI3_X0Y245_ILOGIC_X0Y246_D = LIOB33_X0Y245_IOB_X0Y246_I;
  assign LIOI3_X0Y245_ILOGIC_X0Y245_D = LIOB33_X0Y245_IOB_X0Y245_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y124_D = LIOB33_X0Y123_IOB_X0Y124_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y123_D = LIOB33_X0Y123_IOB_X0Y123_I;
  assign LIOI3_X0Y1_ILOGIC_X0Y2_D = LIOB33_X0Y1_IOB_X0Y2_I;
  assign LIOI3_X0Y1_ILOGIC_X0Y1_D = LIOB33_X0Y1_IOB_X0Y1_I;
  assign RIOB33_X105Y53_IOB_X1Y54_O = CLBLM_R_X7Y132_SLICE_X9Y132_AQ;
  assign RIOB33_X105Y53_IOB_X1Y53_O = CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  assign CLBLL_L_X54Y138_SLICE_X82Y138_A1 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X82Y138_A2 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X82Y138_A3 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X82Y138_A4 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X82Y138_A5 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X82Y138_A6 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X82Y138_AX = CLBLL_L_X4Y137_SLICE_X5Y137_AO5;
  assign CLBLL_L_X54Y138_SLICE_X82Y138_B1 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X82Y138_B2 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X82Y138_B3 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X82Y138_B4 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X82Y138_B5 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X82Y138_B6 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X82Y138_C1 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X82Y138_C2 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X82Y138_C3 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X82Y138_C4 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X82Y138_C5 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X82Y138_C6 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X82Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X54Y138_SLICE_X82Y138_D1 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X82Y138_D2 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X82Y138_D3 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X82Y138_D4 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X82Y138_D5 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X82Y138_D6 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X83Y138_A1 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X83Y138_A2 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X83Y138_A3 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X83Y138_A4 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X83Y138_A5 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X83Y138_A6 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B6 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X83Y138_B1 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X83Y138_B2 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X83Y138_B3 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X83Y138_B4 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X83Y138_B5 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X83Y138_B6 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X83Y138_C1 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X83Y138_C2 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X83Y138_C3 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X83Y138_C4 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X83Y138_C5 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X83Y138_C6 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X83Y138_D1 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X83Y138_D2 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X83Y138_D3 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X83Y138_D4 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X83Y138_D5 = 1'b1;
  assign CLBLL_L_X54Y138_SLICE_X83Y138_D6 = 1'b1;
  assign RIOB33_X105Y55_IOB_X1Y56_O = CLBLM_R_X5Y133_SLICE_X7Y133_CQ;
  assign RIOB33_X105Y55_IOB_X1Y55_O = CLBLL_L_X4Y134_SLICE_X5Y134_AQ;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_B4 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_B5 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_C4 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_C5 = 1'b1;
  assign RIOI3_X105Y103_OLOGIC_X1Y104_D1 = CLBLM_R_X7Y128_SLICE_X8Y128_BQ;
  assign RIOI3_X105Y103_OLOGIC_X1Y104_T1 = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_D1 = CLBLM_L_X16Y136_SLICE_X22Y136_AQ;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_T1 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A1 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A2 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A3 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A4 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A5 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A6 = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_D1 = CLBLM_R_X15Y135_SLICE_X21Y135_AQ;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_AX = LIOB33_X0Y165_IOB_X0Y165_I;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B1 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B2 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B3 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B4 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B5 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B6 = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_T1 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_BX = LIOB33_X0Y151_IOB_X0Y152_I;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C1 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C2 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C3 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C4 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C5 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C6 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_A1 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D1 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D2 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D3 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D4 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D5 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D6 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_A3 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A1 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A2 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A3 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A4 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A5 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A6 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_AX = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B1 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B2 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B3 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B4 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B5 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B6 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_BX = LIOB33_X0Y155_IOB_X0Y155_I;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C1 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C2 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C3 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C4 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C5 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C6 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_AX = RIOB33_X105Y193_IOB_X1Y194_I;
  assign RIOB33_X105Y57_IOB_X1Y58_O = CLBLM_L_X8Y130_SLICE_X10Y130_CQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOB33_X105Y57_IOB_X1Y57_O = CLBLM_R_X7Y137_SLICE_X9Y137_CQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_CX = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_B1 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D1 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D2 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D3 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D4 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D5 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D6 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_B2 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_B3 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_DX = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_B4 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_B5 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_BX = RIOB33_X105Y197_IOB_X1Y197_I;
  assign LIOI3_X0Y247_ILOGIC_X0Y248_D = LIOB33_X0Y247_IOB_X0Y248_I;
  assign LIOI3_X0Y247_ILOGIC_X0Y247_D = LIOB33_X0Y247_IOB_X0Y247_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y126_D = LIOB33_X0Y125_IOB_X0Y126_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y125_D = LIOB33_X0Y125_IOB_X0Y125_I;
  assign LIOI3_X0Y3_ILOGIC_X0Y4_D = LIOB33_X0Y3_IOB_X0Y4_I;
  assign LIOI3_X0Y3_ILOGIC_X0Y3_D = LIOB33_X0Y3_IOB_X0Y3_I;
  assign CLBLM_L_X56Y151_SLICE_X85Y151_A1 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X85Y151_A2 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X85Y151_A3 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X85Y151_A4 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X85Y151_A5 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X85Y151_A6 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X85Y151_B1 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X85Y151_B2 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X85Y151_B3 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X85Y151_B4 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X85Y151_B5 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X85Y151_B6 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X85Y151_C1 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X85Y151_C2 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X85Y151_C3 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X85Y151_C4 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X85Y151_C5 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X85Y151_C6 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X85Y151_D1 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X85Y151_D2 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X85Y151_D3 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X85Y151_D4 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X85Y151_D5 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X85Y151_D6 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X84Y151_A1 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X84Y151_A2 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X84Y151_A3 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X84Y151_A4 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X84Y151_A5 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X84Y151_A6 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X84Y151_AX = CLBLM_L_X10Y136_SLICE_X13Y136_BO6;
  assign CLBLM_L_X56Y151_SLICE_X84Y151_B1 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X84Y151_B2 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X84Y151_B3 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X84Y151_B4 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X84Y151_B5 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X84Y151_B6 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X84Y151_C1 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X84Y151_C2 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X84Y151_C3 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X84Y151_C4 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X84Y151_C5 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X84Y151_C6 = 1'b1;
  assign RIOB33_X105Y59_IOB_X1Y59_O = CLBLM_R_X5Y131_SLICE_X6Y131_AQ;
  assign RIOB33_X105Y59_IOB_X1Y60_O = CLBLM_R_X7Y136_SLICE_X8Y136_BQ;
  assign CLBLM_L_X56Y151_SLICE_X84Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X1Y44_O;
  assign CLBLM_L_X56Y151_SLICE_X84Y151_D1 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X84Y151_D2 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X84Y151_D3 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X84Y151_D4 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X84Y151_D5 = 1'b1;
  assign CLBLM_L_X56Y151_SLICE_X84Y151_D6 = 1'b1;
  assign RIOB33_X105Y121_IOB_X1Y122_O = CLBLM_L_X10Y133_SLICE_X13Y133_CQ;
  assign RIOB33_X105Y121_IOB_X1Y121_O = CLBLM_R_X11Y133_SLICE_X14Y133_BQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C4 = BRAM_R_X17Y135_RAMB18_X1Y54_DO23;
  assign CLBLL_L_X54Y141_SLICE_X82Y141_A1 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X82Y141_A2 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X82Y141_A3 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X82Y141_A4 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X82Y141_A5 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X82Y141_A6 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X82Y141_AX = CLBLM_R_X3Y137_SLICE_X3Y137_AO5;
  assign CLBLL_L_X54Y141_SLICE_X82Y141_B1 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X82Y141_B2 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X82Y141_B3 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X82Y141_B4 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X82Y141_B5 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X82Y141_B6 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X82Y141_C1 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X82Y141_C2 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X82Y141_C3 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X82Y141_C4 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X82Y141_C5 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X82Y141_C6 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X82Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X54Y141_SLICE_X82Y141_D1 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X82Y141_D2 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X82Y141_D3 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X82Y141_D4 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X82Y141_D5 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A6 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X82Y141_D6 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A1 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A2 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B1 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B2 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B3 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A5 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B4 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B5 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B6 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_AX = LIOB33_X0Y161_IOB_X0Y162_I;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_BX = LIOB33_X0Y163_IOB_X0Y163_I;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C6 = CLBLM_R_X3Y158_SLICE_X3Y158_BQ;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C1 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C2 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C3 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C4 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C5 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C6 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_CX = LIOB33_X0Y163_IOB_X0Y164_I;
  assign CLBLL_L_X54Y141_SLICE_X83Y141_A1 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X83Y141_A2 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D3 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D4 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D5 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D6 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X83Y141_A3 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X83Y141_A4 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_DX = LIOB33_X0Y167_IOB_X0Y168_I;
  assign CLBLL_L_X54Y141_SLICE_X83Y141_A5 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X83Y141_A6 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X83Y141_B1 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X83Y141_B2 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X83Y141_B3 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A3 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A4 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X83Y141_B4 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X83Y141_B5 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X83Y141_B6 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A1 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A2 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X83Y141_C1 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X83Y141_C2 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X83Y141_C3 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X83Y141_C4 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X83Y141_C5 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B5 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B6 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X83Y141_C6 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_AX = LIOB33_X0Y169_IOB_X0Y170_I;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B1 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B2 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B3 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B4 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X83Y141_D1 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X83Y141_D2 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X83Y141_D3 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X83Y141_D4 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X83Y141_D5 = 1'b1;
  assign CLBLL_L_X54Y141_SLICE_X83Y141_D6 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C2 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C3 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C4 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C5 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_CX = LIOB33_X0Y171_IOB_X0Y172_I;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D1 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D2 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D3 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D4 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D5 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D6 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_D1 = CLBLM_L_X16Y135_SLICE_X22Y135_BQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_DX = LIOB33_X0Y173_IOB_X0Y173_I;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_T1 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_D1 = CLBLM_L_X16Y135_SLICE_X22Y135_AQ;
  assign RIOI3_X105Y51_OLOGIC_X1Y52_D1 = CLBLM_R_X5Y134_SLICE_X7Y134_CQ;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_T1 = 1'b1;
  assign RIOI3_X105Y51_OLOGIC_X1Y52_T1 = 1'b1;
  assign RIOI3_X105Y51_OLOGIC_X1Y51_D1 = CLBLM_R_X5Y132_SLICE_X7Y132_BQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A2 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO7;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_D1 = CLBLM_L_X8Y130_SLICE_X10Y130_CQ;
  assign RIOI3_X105Y51_OLOGIC_X1Y51_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_D1 = CLBLM_R_X7Y137_SLICE_X9Y137_CQ;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_T1 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B2 = LIOB33_X0Y19_IOB_X0Y19_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B3 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B5 = CLBLM_R_X5Y127_SLICE_X7Y127_BQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B6 = BRAM_L_X6Y125_RAMB18_X0Y50_DO5;
  assign LIOI3_X0Y127_ILOGIC_X0Y128_D = LIOB33_X0Y127_IOB_X0Y128_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y127_D = LIOB33_X0Y127_IOB_X0Y127_I;
  assign RIOB33_X105Y63_IOB_X1Y64_O = CLBLL_L_X54Y96_SLICE_X82Y96_AQ;
  assign RIOB33_X105Y63_IOB_X1Y63_O = CLBLM_R_X7Y137_SLICE_X9Y137_DQ;
  assign LIOI3_X0Y5_ILOGIC_X0Y6_D = LIOB33_X0Y5_IOB_X0Y6_I;
  assign LIOI3_X0Y5_ILOGIC_X0Y5_D = LIOB33_X0Y5_IOB_X0Y5_I;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B4 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO7;
  assign LIOI3_X0Y161_ILOGIC_X0Y162_D = LIOB33_X0Y161_IOB_X0Y162_I;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B5 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO7;
  assign LIOI3_X0Y161_ILOGIC_X0Y161_D = LIOB33_X0Y161_IOB_X0Y161_I;
  assign RIOB33_X105Y65_IOB_X1Y66_O = CLBLM_R_X7Y125_SLICE_X8Y125_AQ;
  assign RIOB33_X105Y65_IOB_X1Y65_O = CLBLM_L_X8Y127_SLICE_X10Y127_AQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_CX = CLBLM_R_X5Y127_SLICE_X6Y127_DO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A1 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A2 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A3 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A4 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A5 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A6 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D1 = BRAM_L_X6Y125_RAMB18_X0Y50_DO0;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_AX = LIOB33_X0Y173_IOB_X0Y174_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D2 = CLBLM_R_X5Y127_SLICE_X6Y127_CQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B1 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B2 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B3 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B4 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B5 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B6 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D3 = LIOB33_SING_X0Y0_IOB_X0Y0_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D4 = CLBLM_R_X5Y127_SLICE_X6Y127_CO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C1 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C2 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C3 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C4 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C5 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C6 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D5 = CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D6 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D1 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D2 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D3 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D4 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D5 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D6 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A1 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A2 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B3 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A3 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A4 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A5 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A6 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C1 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO7;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_AX = LIOB33_X0Y175_IOB_X0Y175_I;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B1 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B2 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B3 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B4 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B5 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B6 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B6 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C4 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_BX = LIOB33_X0Y175_IOB_X0Y176_I;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C5 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C1 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C2 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C3 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C4 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C5 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C6 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C2 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO7;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_CX = LIOB33_X0Y177_IOB_X0Y177_I;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D1 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D2 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D3 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D4 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D5 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D6 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C1 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_DX = LIOB33_X0Y177_IOB_X0Y178_I;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C2 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C3 = BRAM_L_X6Y140_RAMB18_X0Y56_DO23;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C5 = 1'b1;
  assign CLBLM_L_X16Y155_SLICE_X23Y155_A2 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C6 = 1'b1;
  assign CLBLM_L_X16Y155_SLICE_X23Y155_A3 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D3 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C5 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO6;
  assign CLBLM_L_X16Y155_SLICE_X23Y155_B1 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D1 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C6 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D2 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D3 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D4 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D5 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A3 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D6 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_D1 = CLBLM_L_X16Y137_SLICE_X22Y137_AQ;
  assign CLBLM_L_X16Y155_SLICE_X23Y155_C2 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_T1 = 1'b1;
  assign CLBLM_L_X16Y155_SLICE_X23Y155_C3 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_SR = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_L_X16Y155_SLICE_X23Y155_C4 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_D1 = CLBLM_R_X13Y136_SLICE_X18Y136_AQ;
  assign CLBLM_L_X16Y155_SLICE_X23Y155_C5 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_AX = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_L_X16Y155_SLICE_X23Y155_C6 = 1'b1;
  assign RIOB33_X105Y67_IOB_X1Y67_O = CLBLM_L_X8Y127_SLICE_X10Y127_BQ;
  assign RIOB33_X105Y67_IOB_X1Y68_O = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign RIOI3_X105Y53_OLOGIC_X1Y54_D1 = CLBLM_R_X7Y132_SLICE_X9Y132_AQ;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_T1 = 1'b1;
  assign RIOI3_X105Y53_OLOGIC_X1Y54_T1 = 1'b1;
  assign RIOI3_X105Y53_OLOGIC_X1Y53_D1 = CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_D1 = CLBLM_L_X8Y129_SLICE_X10Y129_CQ;
  assign RIOI3_X105Y53_OLOGIC_X1Y53_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_D1 = CLBLM_L_X8Y129_SLICE_X10Y129_BQ;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_T1 = 1'b1;
  assign CLBLM_L_X16Y155_SLICE_X22Y155_A1 = 1'b1;
  assign CLBLM_L_X16Y155_SLICE_X22Y155_A2 = 1'b1;
  assign CLBLM_L_X16Y155_SLICE_X22Y155_A3 = 1'b1;
  assign LIOI3_X0Y129_ILOGIC_X0Y130_D = LIOB33_X0Y129_IOB_X0Y130_I;
  assign CLBLM_L_X16Y155_SLICE_X22Y155_AX = RIOB33_X105Y201_IOB_X1Y202_I;
  assign LIOI3_X0Y129_ILOGIC_X0Y129_D = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLM_L_X16Y155_SLICE_X22Y155_B1 = 1'b1;
  assign CLBLM_L_X16Y155_SLICE_X22Y155_B2 = 1'b1;
  assign CLBLM_L_X16Y155_SLICE_X22Y155_B3 = 1'b1;
  assign CLBLM_L_X16Y155_SLICE_X22Y155_B4 = 1'b1;
  assign LIOI3_X0Y9_ILOGIC_X0Y10_D = LIOB33_X0Y9_IOB_X0Y10_I;
  assign LIOI3_X0Y9_ILOGIC_X0Y9_D = LIOB33_X0Y9_IOB_X0Y9_I;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D1 = 1'b1;
  assign CLBLM_L_X16Y155_SLICE_X22Y155_C6 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D3 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X16Y155_SLICE_X22Y155_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign RIOB33_X105Y69_IOB_X1Y70_O = CLBLM_L_X8Y129_SLICE_X10Y129_CQ;
  assign RIOB33_X105Y69_IOB_X1Y69_O = CLBLM_L_X8Y129_SLICE_X10Y129_BQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D4 = CLBLM_R_X5Y135_SLICE_X6Y135_AO6;
  assign CLBLM_L_X16Y155_SLICE_X22Y155_D1 = 1'b1;
  assign CLBLM_L_X16Y155_SLICE_X22Y155_D2 = 1'b1;
  assign CLBLM_L_X16Y155_SLICE_X22Y155_D3 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D5 = 1'b1;
  assign CLBLM_L_X16Y155_SLICE_X22Y155_D4 = 1'b1;
  assign CLBLM_L_X16Y155_SLICE_X22Y155_D5 = 1'b1;
  assign RIOB33_X105Y123_IOB_X1Y123_O = CLBLM_L_X12Y132_SLICE_X16Y132_BQ;
  assign CLBLM_L_X16Y155_SLICE_X22Y155_D6 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D6 = CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A1 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A2 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A3 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A4 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A5 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A6 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_AX = LIOB33_X0Y179_IOB_X0Y179_I;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B1 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B2 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B3 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B4 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B5 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B6 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_BX = LIOB33_X0Y179_IOB_X0Y180_I;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C1 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C2 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C3 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C4 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C5 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C6 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D1 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D2 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D3 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D4 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D5 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D6 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A1 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A2 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A3 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A4 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A5 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A6 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_AX = LIOB33_X0Y181_IOB_X0Y181_I;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B1 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B2 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B3 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B4 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B5 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B6 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_BX = LIOB33_X0Y181_IOB_X0Y182_I;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C1 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C2 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C3 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C4 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C5 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C6 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_CX = LIOB33_X0Y183_IOB_X0Y183_I;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D1 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D2 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D3 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D4 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D5 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D6 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_DX = LIOB33_X0Y183_IOB_X0Y184_I;
  assign RIOB33_X105Y71_IOB_X1Y72_O = CLBLM_R_X7Y128_SLICE_X9Y128_AQ;
  assign RIOB33_X105Y71_IOB_X1Y71_O = CLBLL_L_X54Y101_SLICE_X82Y101_AQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A1 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A2 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A3 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A4 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A5 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A6 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B1 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B2 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B3 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B4 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B5 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B6 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C1 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C2 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C3 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C4 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C5 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C6 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D1 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D2 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D3 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D4 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D5 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D6 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A1 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A2 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A3 = BRAM_R_X17Y135_RAMB18_X1Y54_DO17;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A4 = CLBLL_L_X4Y131_SLICE_X4Y131_CQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A5 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A6 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B1 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B2 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B3 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B4 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B5 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B6 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C1 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C2 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C3 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C4 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C5 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C6 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D1 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D2 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D3 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D4 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D5 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D6 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_D1 = CLBLM_L_X16Y137_SLICE_X22Y137_BQ;
  assign RIOI3_X105Y55_OLOGIC_X1Y56_D1 = CLBLM_R_X5Y133_SLICE_X7Y133_CQ;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_T1 = 1'b1;
  assign RIOI3_X105Y55_OLOGIC_X1Y56_T1 = 1'b1;
  assign RIOI3_X105Y55_OLOGIC_X1Y55_D1 = CLBLL_L_X4Y134_SLICE_X5Y134_AQ;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_D1 = CLBLM_L_X8Y130_SLICE_X11Y130_DQ;
  assign RIOI3_X105Y55_OLOGIC_X1Y55_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_D1 = CLBLM_L_X8Y131_SLICE_X11Y131_CQ;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_T1 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A1 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A2 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A3 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A4 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A5 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A6 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B1 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B2 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B3 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B4 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B5 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B6 = 1'b1;
  assign RIOB33_X105Y73_IOB_X1Y73_O = CLBLM_L_X8Y130_SLICE_X11Y130_BQ;
  assign RIOB33_X105Y73_IOB_X1Y74_O = CLBLM_R_X7Y130_SLICE_X9Y130_DQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C1 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C2 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C3 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C4 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C5 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C6 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D1 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D2 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D3 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D4 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D5 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D6 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A1 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A2 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A3 = CLBLM_R_X5Y125_SLICE_X7Y125_AQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A4 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A5 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A6 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B1 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B2 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO3;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B3 = CLBLM_R_X5Y126_SLICE_X6Y126_AQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B4 = 1'b1;
  assign LIOI3_X0Y133_ILOGIC_X0Y134_D = LIOB33_X0Y133_IOB_X0Y134_I;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B5 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B6 = 1'b1;
  assign LIOI3_X0Y133_ILOGIC_X0Y133_D = LIOB33_X0Y133_IOB_X0Y133_I;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C1 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C2 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C3 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C4 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C5 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C6 = 1'b1;
  assign RIOI3_X105Y177_ILOGIC_X1Y178_D = RIOB33_X105Y177_IOB_X1Y178_I;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D1 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D2 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D3 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D4 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D5 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D6 = 1'b1;
  assign LIOI3_X0Y11_ILOGIC_X0Y12_D = LIOB33_X0Y11_IOB_X0Y12_I;
  assign LIOI3_X0Y11_ILOGIC_X0Y11_D = LIOB33_X0Y11_IOB_X0Y11_I;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A1 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A2 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A3 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A4 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A5 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A6 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B1 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B2 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B3 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B4 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B5 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B6 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C1 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C2 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C3 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C4 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C5 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C6 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D1 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D2 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D3 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D4 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D5 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D6 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A1 = CLBLM_R_X3Y131_SLICE_X3Y131_DQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A2 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A3 = BRAM_R_X17Y135_RAMB18_X1Y54_DO20;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A4 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A5 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A6 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A1 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A2 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A3 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A4 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B2 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B3 = BRAM_R_X17Y135_RAMB18_X1Y54_DO23;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B4 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A5 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A6 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_AX = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B1 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B1 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B2 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B3 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B4 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B5 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B6 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_BX = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C1 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C2 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C3 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C4 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C5 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C6 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C5 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D1 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D3 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D4 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D5 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_CX = LIOB33_X0Y187_IOB_X0Y188_I;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D2 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D1 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D2 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D3 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D4 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D5 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D6 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_DX = LIOB33_X0Y189_IOB_X0Y189_I;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D6 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A1 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A2 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A3 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A4 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A5 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A6 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_AX = LIOB33_X0Y189_IOB_X0Y190_I;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B1 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B2 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B3 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B4 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B5 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B6 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_BX = LIOB33_X0Y191_IOB_X0Y191_I;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C1 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C2 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C3 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C4 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C5 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C6 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_CX = LIOB33_X0Y191_IOB_X0Y192_I;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D1 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D2 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D3 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D4 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D5 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D6 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_DX = LIOB33_X0Y193_IOB_X0Y193_I;
  assign RIOB33_X105Y75_IOB_X1Y76_O = CLBLM_L_X10Y132_SLICE_X12Y132_AQ;
  assign RIOB33_X105Y75_IOB_X1Y75_O = CLBLM_L_X8Y130_SLICE_X10Y130_DQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A1 = CLBLM_L_X8Y130_SLICE_X10Y130_B5Q;
  assign RIOI3_TBYTESRC_X105Y193_ILOGIC_X1Y194_D = RIOB33_X105Y193_IOB_X1Y194_I;
  assign RIOI3_TBYTESRC_X105Y193_ILOGIC_X1Y193_D = RIOB33_X105Y193_IOB_X1Y193_I;
  assign RIOB33_X105Y77_IOB_X1Y78_O = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign RIOB33_X105Y77_IOB_X1Y77_O = CLBLM_L_X8Y130_SLICE_X11Y130_CQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A1 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A2 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A3 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A4 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A5 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A6 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B1 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B2 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B3 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B4 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B5 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B6 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C1 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C2 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C3 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C4 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C5 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C6 = 1'b1;
  assign RIOI3_X105Y59_OLOGIC_X1Y60_D1 = CLBLM_R_X7Y136_SLICE_X8Y136_BQ;
  assign RIOI3_X105Y59_OLOGIC_X1Y60_T1 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D1 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D2 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D3 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D4 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D5 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D6 = 1'b1;
  assign RIOI3_X105Y59_OLOGIC_X1Y59_D1 = CLBLM_R_X5Y131_SLICE_X6Y131_AQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A1 = CLBLM_R_X5Y126_SLICE_X7Y126_AQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A2 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A3 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO4;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A4 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A5 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_D1 = CLBLM_L_X10Y131_SLICE_X13Y131_AQ;
  assign RIOI3_X105Y59_OLOGIC_X1Y59_T1 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B1 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B2 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO5;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B3 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B4 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B5 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_T1 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C1 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C2 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C3 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C4 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C5 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C6 = CLBLM_R_X5Y127_SLICE_X6Y127_B5Q;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_D1 = CLBLM_L_X12Y132_SLICE_X16Y132_CQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D1 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D2 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D3 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D4 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D5 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_T1 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A1 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A2 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A3 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A4 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A5 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A6 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B1 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B2 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B3 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B4 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B5 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B6 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C1 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C2 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C3 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C4 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C5 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C6 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D1 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D2 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D3 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D4 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D5 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D6 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A1 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO3;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A2 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A3 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A4 = CLBLM_R_X7Y132_SLICE_X8Y132_BQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A5 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A6 = 1'b1;
  assign LIOI3_X0Y135_ILOGIC_X0Y136_D = LIOB33_X0Y135_IOB_X0Y136_I;
  assign LIOI3_X0Y135_ILOGIC_X0Y135_D = LIOB33_X0Y135_IOB_X0Y135_I;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_A1 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_A2 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_A3 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_A4 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_A5 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B3 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B4 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO5;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_A6 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B1 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_AX = LIOB33_X0Y195_IOB_X0Y196_I;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B2 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_B1 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_B2 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C1 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_B3 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_B4 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C4 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_B5 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C6 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_B6 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_BX = LIOB33_X0Y197_IOB_X0Y198_I;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_C1 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_C2 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_C3 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_C4 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_C5 = 1'b1;
  assign LIOI3_X0Y15_ILOGIC_X0Y16_D = LIOB33_X0Y15_IOB_X0Y16_I;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_C6 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOI3_X0Y15_ILOGIC_X0Y15_D = LIOB33_X0Y15_IOB_X0Y15_I;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D1 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D2 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_CX = LIOB33_X0Y201_IOB_X0Y202_I;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D3 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_D1 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_D2 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_D3 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_D4 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_D5 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_D6 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_A1 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_A2 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_A3 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_A4 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_A5 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_A6 = 1'b1;
  assign RIOB33_X105Y79_IOB_X1Y79_O = CLBLL_L_X54Y105_SLICE_X82Y105_AQ;
  assign RIOB33_X105Y79_IOB_X1Y80_O = CLBLM_L_X8Y131_SLICE_X11Y131_BQ;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_AX = LIOB33_X0Y221_IOB_X0Y222_I;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_B1 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_B2 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_B3 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_B4 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_B5 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_B6 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_BX = LIOB33_X0Y225_IOB_X0Y225_I;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_C1 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_C2 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_C3 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_C4 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_C5 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_C6 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLL_L_X54Y119_SLICE_X82Y119_A1 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_CX = LIOB33_X0Y231_IOB_X0Y231_I;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_D1 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_D2 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X82Y119_A2 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_D3 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_D4 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_D5 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_D6 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X82Y119_A3 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_DX = LIOB33_X0Y239_IOB_X0Y240_I;
  assign CLBLL_L_X54Y119_SLICE_X82Y119_A4 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X82Y119_A5 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X82Y119_A6 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X82Y119_AX = CLBLM_R_X5Y134_SLICE_X6Y134_BO5;
  assign CLBLL_L_X54Y119_SLICE_X82Y119_B1 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A2 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A3 = CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A4 = BRAM_R_X17Y135_RAMB18_X1Y54_DO16;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A5 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A1 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO0;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A6 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X82Y119_B2 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X82Y119_B3 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B1 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B3 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B4 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B5 = CLBLL_L_X4Y129_SLICE_X4Y129_AQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B6 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X82Y119_B4 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B2 = BRAM_L_X6Y135_RAMB18_X0Y54_DO17;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C1 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C2 = BRAM_L_X6Y135_RAMB18_X0Y54_DO21;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C3 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C4 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C5 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C6 = CLBLM_R_X3Y130_SLICE_X3Y130_AQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D1 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO2;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D2 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D3 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D4 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D5 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D6 = CLBLL_L_X4Y131_SLICE_X4Y131_BQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A1 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO7;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A2 = CLBLM_L_X8Y130_SLICE_X10Y130_A5Q;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A3 = BRAM_L_X6Y125_RAMB18_X0Y50_DO7;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A5 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A6 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B1 = CLBLM_L_X8Y130_SLICE_X10Y130_B5Q;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B2 = BRAM_L_X6Y125_RAMB18_X0Y50_DO19;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B3 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B4 = BRAM_L_X6Y135_RAMB18_X0Y54_DO3;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B5 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B6 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C1 = CLBLL_L_X4Y130_SLICE_X5Y130_AQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C2 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C3 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C4 = BRAM_L_X6Y140_RAMB18_X0Y56_DO2;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C5 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C6 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D1 = CLBLM_R_X5Y128_SLICE_X6Y128_AQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D2 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D3 = BRAM_L_X6Y135_RAMB18_X0Y54_DO19;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D4 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D5 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D6 = 1'b1;
  assign LIOB33_SING_X0Y100_IOB_X0Y100_O = CLBLL_L_X2Y141_SLICE_X0Y141_AQ;
  assign RIOB33_X105Y81_IOB_X1Y82_O = CLBLM_L_X8Y130_SLICE_X11Y130_DQ;
  assign RIOB33_X105Y81_IOB_X1Y81_O = CLBLM_L_X8Y131_SLICE_X11Y131_CQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A1 = CLBLL_L_X4Y131_SLICE_X5Y131_B5Q;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A2 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A3 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A4 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A5 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A6 = BRAM_L_X6Y135_RAMB18_X0Y54_DO22;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B1 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B2 = CLBLM_R_X5Y131_SLICE_X7Y131_A5Q;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B3 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B4 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B5 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B6 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO0;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C1 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C2 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C3 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C4 = CLBLL_L_X4Y131_SLICE_X4Y131_AQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C5 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D1 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO0;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D2 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO0;
  assign CLBLL_L_X54Y119_SLICE_X83Y119_B1 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D3 = BRAM_R_X17Y135_RAMB18_X1Y54_DO23;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D4 = CLBLM_R_X3Y131_SLICE_X3Y131_BQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D5 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO7;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D6 = BRAM_L_X6Y135_RAMB18_X0Y54_DO16;
  assign CLBLL_L_X54Y119_SLICE_X83Y119_B2 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X83Y119_B3 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A1 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A2 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A3 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A4 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO5;
  assign CLBLL_L_X54Y119_SLICE_X83Y119_B4 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A5 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A6 = CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  assign CLBLL_L_X54Y119_SLICE_X83Y119_B5 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B1 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO3;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B2 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B3 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B4 = 1'b1;
  assign CLBLL_L_X54Y119_SLICE_X83Y119_B6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B5 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B6 = CLBLM_R_X5Y133_SLICE_X6Y133_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C1 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO2;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C2 = BRAM_R_X17Y135_RAMB18_X1Y54_DO19;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C3 = CLBLM_R_X5Y126_SLICE_X6Y126_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C4 = BRAM_R_X17Y135_RAMB18_X1Y54_DO18;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C5 = BRAM_L_X6Y135_RAMB18_X0Y54_DO19;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C6 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO3;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D1 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D2 = BRAM_R_X17Y135_RAMB18_X1Y54_DO17;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D3 = CLBLM_R_X5Y125_SLICE_X7Y125_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D4 = BRAM_L_X6Y135_RAMB18_X0Y54_DO17;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D5 = BRAM_R_X17Y135_RAMB18_X1Y54_DO16;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D6 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO0;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A1 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A2 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A3 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A4 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A5 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A6 = 1'b1;
  assign RIOI3_X105Y61_OLOGIC_X1Y62_D1 = CLBLL_L_X4Y134_SLICE_X5Y134_BQ;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B1 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B2 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B3 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B4 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B5 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B6 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C1 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C2 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C3 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C4 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C5 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C6 = 1'b1;
  assign RIOI3_X105Y61_OLOGIC_X1Y62_T1 = 1'b1;
  assign RIOI3_X105Y61_OLOGIC_X1Y61_D1 = CLBLL_L_X4Y135_SLICE_X5Y135_BQ;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D1 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D2 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D3 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D4 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D5 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_D1 = CLBLM_R_X7Y130_SLICE_X8Y130_BQ;
  assign RIOI3_X105Y61_OLOGIC_X1Y61_T1 = 1'b1;
  assign RIOB33_X105Y83_IOB_X1Y84_O = CLBLM_L_X10Y132_SLICE_X12Y132_BQ;
  assign RIOB33_X105Y83_IOB_X1Y83_O = CLBLM_L_X8Y131_SLICE_X10Y131_BQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A1 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO7;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A2 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO0;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A3 = CLBLM_R_X3Y131_SLICE_X3Y131_AQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A4 = BRAM_R_X17Y135_RAMB18_X1Y54_DO7;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A5 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO0;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A6 = BRAM_L_X6Y135_RAMB18_X0Y54_DO0;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_T1 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_A1 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_A2 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B1 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO7;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B2 = CLBLM_L_X8Y135_SLICE_X10Y135_A5Q;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B3 = CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B4 = BRAM_L_X6Y135_RAMB18_X0Y54_DO7;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B5 = CLBLM_L_X16Y151_SLICE_X22Y151_DQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B6 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_A3 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_A4 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_A5 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_A6 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C1 = CLBLM_R_X25Y153_SLICE_X36Y153_AQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C2 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C3 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C4 = CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C5 = CLBLM_L_X10Y135_SLICE_X12Y135_A5Q;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C6 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_B2 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_B3 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_B4 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_B5 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_B6 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_BX = LIOB33_X0Y205_IOB_X0Y206_I;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_C1 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_C2 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_C3 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D1 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D2 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D3 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D4 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D5 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D6 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_CX = LIOB33_X0Y219_IOB_X0Y220_I;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_D1 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_D2 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_D6 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_D3 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_D4 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_DX = LIOB33_X0Y221_IOB_X0Y221_I;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_D5 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_A1 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_A2 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_A3 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_A4 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_A5 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_A6 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_AX = LIOB33_X0Y227_IOB_X0Y227_I;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_B1 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_B2 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_B3 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_B4 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_B5 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_B6 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_BX = LIOB33_X0Y243_IOB_X0Y243_I;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_C1 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_C2 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_C3 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_C4 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_C5 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_C6 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_CX = LIOB33_X0Y247_IOB_X0Y248_I;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_D1 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_D2 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_D3 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_D4 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_D5 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_D6 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_DX = LIOB33_SING_X0Y249_IOB_X0Y249_I;
  assign LIOI3_X0Y139_ILOGIC_X0Y140_D = LIOB33_X0Y139_IOB_X0Y140_I;
  assign LIOI3_X0Y139_ILOGIC_X0Y139_D = LIOB33_X0Y139_IOB_X0Y139_I;
  assign RIOI3_X105Y183_ILOGIC_X1Y184_D = RIOB33_X105Y183_IOB_X1Y184_I;
  assign RIOI3_X105Y183_ILOGIC_X1Y183_D = RIOB33_X105Y183_IOB_X1Y183_I;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A1 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A2 = BRAM_L_X6Y130_RAMB18_X0Y52_DO0;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A3 = LIOB33_X0Y131_IOB_X0Y132_I;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A4 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO0;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A5 = CLBLM_L_X8Y132_SLICE_X11Y132_A5Q;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A6 = 1'b1;
  assign LIOI3_X0Y17_ILOGIC_X0Y18_D = LIOB33_X0Y17_IOB_X0Y18_I;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B1 = BRAM_L_X6Y140_RAMB18_X0Y56_DO22;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B2 = 1'b1;
  assign LIOI3_X0Y17_ILOGIC_X0Y17_D = LIOB33_X0Y17_IOB_X0Y17_I;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B3 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B4 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B5 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B6 = CLBLM_R_X5Y132_SLICE_X7Y132_B5Q;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C1 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C2 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C3 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C4 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C5 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C6 = CLBLL_L_X4Y132_SLICE_X4Y132_BQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D1 = CLBLL_L_X4Y131_SLICE_X4Y131_AQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D2 = BRAM_R_X17Y135_RAMB18_X1Y54_DO17;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D3 = BRAM_L_X6Y135_RAMB18_X0Y54_DO17;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D4 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D5 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO0;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D6 = BRAM_L_X6Y135_RAMB18_X0Y54_DO16;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A1 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO7;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A2 = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A3 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A4 = BRAM_R_X17Y135_RAMB18_X1Y54_DO23;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A5 = CLBLM_R_X5Y158_SLICE_X6Y158_DQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A6 = CLBLM_L_X8Y132_SLICE_X10Y132_CO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B1 = CLBLM_L_X8Y132_SLICE_X10Y132_DO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B2 = BRAM_R_X17Y135_RAMB18_X1Y54_DO23;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B4 = CLBLM_R_X5Y158_SLICE_X6Y158_CQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B5 = CLBLL_L_X4Y131_SLICE_X4Y131_CQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B6 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B3 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO7;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C1 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO2;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C2 = BRAM_R_X17Y135_RAMB18_X1Y54_DO18;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C3 = BRAM_L_X6Y135_RAMB18_X0Y54_DO19;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C4 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO3;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C5 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO3;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C6 = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D1 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D2 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D3 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO0;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D4 = CLBLL_L_X4Y131_SLICE_X4Y131_CQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D5 = BRAM_L_X6Y135_RAMB18_X0Y54_DO17;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D6 = BRAM_R_X17Y135_RAMB18_X1Y54_DO16;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A1 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A2 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A3 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A4 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A5 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A6 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B1 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B2 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B3 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B4 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B5 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B6 = 1'b1;
  assign RIOB33_X105Y85_IOB_X1Y85_O = CLBLM_L_X10Y132_SLICE_X12Y132_CQ;
  assign RIOB33_X105Y85_IOB_X1Y86_O = CLBLM_L_X8Y132_SLICE_X11Y132_CQ;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C1 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C2 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C3 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C4 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C5 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C6 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D1 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D2 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D3 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D4 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D5 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D6 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A1 = BRAM_R_X17Y135_RAMB18_X1Y54_DO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A2 = CLBLM_R_X3Y132_SLICE_X2Y132_BQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A3 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO7;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A4 = BRAM_L_X6Y135_RAMB18_X0Y54_DO7;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A5 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO7;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A6 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO6;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_A1 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_A2 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_A3 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_A4 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_A5 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_A6 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B1 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO6;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_AX = LIOB33_X0Y213_IOB_X0Y214_I;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B2 = BRAM_R_X17Y135_RAMB18_X1Y54_DO5;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_B1 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_B2 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_B3 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_B4 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_B5 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_B6 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B5 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO5;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B6 = BRAM_L_X6Y135_RAMB18_X0Y54_DO6;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_BX = LIOB33_X0Y217_IOB_X0Y218_I;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_C1 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_C2 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_C3 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_C4 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_C5 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_C6 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C5 = CLBLM_L_X8Y137_SLICE_X10Y137_B5Q;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D1 = CLBLM_L_X8Y137_SLICE_X10Y137_A5Q;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D2 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D3 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_CX = LIOB33_X0Y223_IOB_X0Y223_I;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D4 = CLBLM_R_X25Y153_SLICE_X36Y153_BQ;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_D1 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_D2 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_D3 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_D4 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_D5 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_D6 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D5 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_DX = LIOB33_X0Y223_IOB_X0Y224_I;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D6 = CLBLM_L_X10Y136_SLICE_X12Y136_AO6;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_A1 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_A2 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_A3 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_A4 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_A5 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_A6 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_AX = LIOB33_X0Y225_IOB_X0Y226_I;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_B1 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_B2 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_B3 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_B4 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_B5 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_B6 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_BX = LIOB33_X0Y233_IOB_X0Y234_I;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_C1 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_C2 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_C3 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_C4 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_C5 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_C6 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_CX = LIOB33_X0Y235_IOB_X0Y236_I;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_D1 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_D2 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_D3 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_D4 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_D5 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_D6 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C3 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_DX = LIOB33_X0Y237_IOB_X0Y238_I;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C4 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C6 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A1 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A2 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO7;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A3 = CLBLM_R_X3Y134_SLICE_X2Y134_AQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A4 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A5 = BRAM_L_X6Y135_RAMB18_X0Y54_DO23;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A6 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B1 = BRAM_R_X17Y135_RAMB18_X1Y54_DO19;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B2 = BRAM_L_X6Y135_RAMB18_X0Y54_DO20;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B3 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO4;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B4 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO3;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B5 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO4;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B6 = CLBLM_R_X3Y131_SLICE_X3Y131_DQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C1 = CLBLM_L_X8Y133_SLICE_X11Y133_AO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C2 = BRAM_L_X6Y135_RAMB18_X0Y54_DO16;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C3 = CLBLM_R_X5Y158_SLICE_X6Y158_AQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C4 = CLBLM_R_X5Y131_SLICE_X7Y131_A5Q;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C5 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C6 = CLBLM_L_X8Y130_SLICE_X11Y130_AO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D1 = CLBLM_R_X3Y158_SLICE_X2Y158_DQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D2 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D3 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D4 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D5 = CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D6 = CLBLM_R_X3Y131_SLICE_X3Y131_BQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A1 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A2 = CLBLM_R_X3Y158_SLICE_X2Y158_BQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A3 = BRAM_L_X6Y135_RAMB18_X0Y54_DO23;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A4 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO7;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A5 = CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A6 = CLBLM_L_X8Y133_SLICE_X10Y133_CO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B1 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B2 = CLBLM_R_X5Y158_SLICE_X6Y158_BQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B3 = CLBLM_L_X8Y133_SLICE_X10Y133_DO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B4 = CLBLM_R_X5Y133_SLICE_X6Y133_AQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B5 = BRAM_L_X6Y135_RAMB18_X0Y54_DO23;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B6 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO7;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C1 = CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C2 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO4;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C3 = BRAM_L_X6Y135_RAMB18_X0Y54_DO19;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C4 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO3;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C5 = BRAM_R_X17Y135_RAMB18_X1Y54_DO20;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C6 = BRAM_L_X6Y135_RAMB18_X0Y54_DO20;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D1 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO2;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D2 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO3;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D3 = BRAM_R_X17Y135_RAMB18_X1Y54_DO19;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D4 = BRAM_L_X6Y135_RAMB18_X0Y54_DO18;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D5 = BRAM_L_X6Y135_RAMB18_X0Y54_DO19;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D6 = CLBLM_R_X5Y133_SLICE_X6Y133_AQ;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_B1 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_B2 = 1'b1;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_B3 = CLBLM_R_X3Y132_SLICE_X2Y132_BQ;
  assign RIOB33_X105Y87_IOB_X1Y88_O = CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  assign RIOB33_X105Y87_IOB_X1Y87_O = CLBLM_L_X10Y132_SLICE_X12Y132_DQ;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_B4 = CLBLM_R_X25Y154_SLICE_X36Y154_CQ;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_B5 = 1'b1;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_B6 = CLBLM_R_X11Y136_SLICE_X14Y136_AO6;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_C1 = CLBLM_R_X11Y136_SLICE_X14Y136_BO6;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_C2 = 1'b1;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_C3 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_C4 = CLBLM_R_X25Y154_SLICE_X36Y154_BQ;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_C5 = 1'b1;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_C6 = CLBLM_R_X3Y132_SLICE_X2Y132_AQ;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C1 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C2 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C3 = 1'b1;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_D2 = CLBLM_L_X10Y136_SLICE_X13Y136_CO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C4 = 1'b1;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_D3 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_D4 = 1'b1;
  assign RIOI3_X105Y65_OLOGIC_X1Y66_D1 = CLBLM_R_X7Y125_SLICE_X8Y125_AQ;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_D5 = CLBLM_R_X3Y131_SLICE_X3Y131_B5Q;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_D6 = 1'b1;
  assign RIOI3_X105Y65_OLOGIC_X1Y66_T1 = 1'b1;
  assign RIOI3_X105Y65_OLOGIC_X1Y65_D1 = CLBLM_L_X8Y127_SLICE_X10Y127_AQ;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_D1 = CLBLM_L_X10Y133_SLICE_X13Y133_BQ;
  assign RIOI3_X105Y65_OLOGIC_X1Y65_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_D1 = CLBLM_R_X11Y133_SLICE_X14Y133_AQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A1 = BRAM_R_X17Y135_RAMB18_X1Y54_DO20;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A2 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO5;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A3 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO5;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A4 = BRAM_L_X6Y135_RAMB18_X0Y54_DO21;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A5 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO4;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A6 = CLBLM_R_X3Y132_SLICE_X3Y132_BQ;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_T1 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B1 = CLBLM_L_X8Y132_SLICE_X11Y132_DO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B2 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO7;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B3 = CLBLL_L_X4Y131_SLICE_X4Y131_AQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B4 = CLBLM_R_X3Y155_SLICE_X2Y155_CQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B5 = BRAM_L_X6Y135_RAMB18_X0Y54_DO23;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B6 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X16Y157_SLICE_X23Y157_A5 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C1 = BRAM_L_X6Y135_RAMB18_X0Y54_DO21;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C2 = CLBLM_R_X5Y132_SLICE_X6Y132_AQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C3 = BRAM_L_X6Y135_RAMB18_X0Y54_DO20;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C4 = BRAM_R_X17Y135_RAMB18_X1Y54_DO21;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C5 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO4;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C6 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO5;
  assign CLBLM_L_X16Y157_SLICE_X23Y157_A6 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D1 = CLBLM_L_X8Y134_SLICE_X11Y134_AO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D2 = CLBLM_R_X3Y132_SLICE_X3Y132_BQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D3 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D4 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D5 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D6 = CLBLM_R_X3Y157_SLICE_X2Y157_BQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A1 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A2 = BRAM_L_X6Y140_RAMB18_X0Y56_DO20;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A3 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A4 = CLBLM_R_X5Y133_SLICE_X6Y133_BQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A5 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A6 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B1 = BRAM_L_X6Y135_RAMB18_X0Y54_DO18;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B2 = BRAM_R_X17Y135_RAMB18_X1Y54_DO17;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B3 = CLBLM_R_X3Y131_SLICE_X3Y131_CQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B4 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO2;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B5 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B6 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO2;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C1 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C2 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO2;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C3 = BRAM_L_X6Y135_RAMB18_X0Y54_DO17;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C4 = BRAM_R_X17Y135_RAMB18_X1Y54_DO18;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C5 = BRAM_L_X6Y135_RAMB18_X0Y54_DO18;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C6 = CLBLL_L_X4Y131_SLICE_X4Y131_BQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOB33_X105Y89_IOB_X1Y89_O = CLBLM_R_X11Y130_SLICE_X14Y130_AQ;
  assign RIOB33_X105Y89_IOB_X1Y90_O = CLBLM_L_X10Y130_SLICE_X12Y130_BQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D1 = CLBLM_R_X7Y125_SLICE_X8Y125_C5Q;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D2 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO2;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D3 = BRAM_R_X17Y135_RAMB18_X1Y54_DO1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D4 = BRAM_L_X6Y135_RAMB18_X0Y54_DO2;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D5 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D6 = BRAM_R_X17Y135_RAMB18_X1Y54_DO2;
  assign LIOI3_X0Y141_ILOGIC_X0Y142_D = LIOB33_X0Y141_IOB_X0Y142_I;
  assign LIOI3_X0Y141_ILOGIC_X0Y141_D = LIOB33_X0Y141_IOB_X0Y141_I;
  assign CLBLM_L_X16Y157_SLICE_X23Y157_C1 = 1'b1;
  assign CLBLM_L_X16Y157_SLICE_X23Y157_C2 = 1'b1;
  assign RIOI3_X105Y185_ILOGIC_X1Y186_D = RIOB33_X105Y185_IOB_X1Y186_I;
  assign CLBLM_L_X16Y157_SLICE_X23Y157_C3 = 1'b1;
  assign RIOI3_X105Y185_ILOGIC_X1Y185_D = RIOB33_X105Y185_IOB_X1Y185_I;
  assign CLBLM_L_X16Y157_SLICE_X23Y157_C5 = 1'b1;
  assign LIOI3_X0Y21_ILOGIC_X0Y22_D = LIOB33_X0Y21_IOB_X0Y22_I;
  assign CLBLM_L_X16Y157_SLICE_X23Y157_C6 = 1'b1;
  assign LIOI3_X0Y21_ILOGIC_X0Y21_D = LIOB33_X0Y21_IOB_X0Y21_I;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_T1 = 1'b1;
  assign CLBLM_L_X16Y157_SLICE_X22Y157_A5 = 1'b1;
  assign CLBLM_L_X16Y157_SLICE_X22Y157_A6 = 1'b1;
  assign CLBLM_L_X16Y157_SLICE_X22Y157_AX = RIOB33_X105Y203_IOB_X1Y203_I;
  assign CLBLM_L_X16Y157_SLICE_X22Y157_B1 = 1'b1;
  assign CLBLM_L_X16Y157_SLICE_X22Y157_B2 = 1'b1;
  assign CLBLM_L_X16Y157_SLICE_X22Y157_B3 = 1'b1;
  assign CLBLM_L_X16Y157_SLICE_X22Y157_B4 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A1 = CLBLM_R_X3Y131_SLICE_X3Y131_DQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A2 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A3 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO7;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A4 = CLBLM_L_X8Y133_SLICE_X11Y133_BO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A5 = CLBLL_L_X4Y156_SLICE_X5Y156_BQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A6 = BRAM_R_X17Y135_RAMB18_X1Y54_DO23;
  assign CLBLM_L_X16Y157_SLICE_X22Y157_B5 = 1'b1;
  assign CLBLM_L_X16Y157_SLICE_X22Y157_B6 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B1 = BRAM_R_X17Y135_RAMB18_X1Y54_DO21;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B2 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B3 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B4 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO5;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B5 = CLBLM_R_X3Y132_SLICE_X2Y132_CQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B6 = BRAM_L_X6Y135_RAMB18_X0Y54_DO22;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C1 = CLBLL_L_X4Y155_SLICE_X4Y155_DQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C2 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C3 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C4 = CLBLM_R_X3Y132_SLICE_X2Y132_CQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C5 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C6 = CLBLM_L_X8Y135_SLICE_X11Y135_BO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D1 = CLBLM_R_X5Y132_SLICE_X6Y132_AQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D2 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D3 = CLBLL_L_X2Y158_SLICE_X0Y158_DQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D4 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D5 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D6 = CLBLM_L_X8Y134_SLICE_X11Y134_CO6;
  assign CLBLM_L_X16Y157_SLICE_X22Y157_C1 = 1'b1;
  assign CLBLM_L_X16Y157_SLICE_X22Y157_C2 = 1'b1;
  assign CLBLM_L_X16Y157_SLICE_X22Y157_C3 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A1 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A2 = CLBLM_L_X8Y135_SLICE_X10Y135_A5Q;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A3 = LIOB33_X0Y133_IOB_X0Y133_I;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A5 = BRAM_L_X6Y130_RAMB18_X0Y52_DO1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A6 = 1'b1;
  assign CLBLM_L_X16Y157_SLICE_X22Y157_C4 = 1'b1;
  assign RIOB33_X105Y91_IOB_X1Y91_O = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_L_X16Y157_SLICE_X22Y157_C5 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B1 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO5;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B2 = CLBLL_L_X4Y132_SLICE_X4Y132_BQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B3 = BRAM_R_X17Y135_RAMB18_X1Y54_DO22;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B4 = BRAM_L_X6Y135_RAMB18_X0Y54_DO21;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B5 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B6 = BRAM_L_X6Y135_RAMB18_X0Y54_DO22;
  assign CLBLM_L_X16Y157_SLICE_X22Y157_C6 = 1'b1;
  assign CLBLM_L_X16Y157_SLICE_X22Y157_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y68_D = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C1 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C2 = CLBLM_R_X3Y158_SLICE_X2Y158_CQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C3 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C4 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C5 = CLBLM_L_X8Y135_SLICE_X10Y135_BO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C6 = CLBLL_L_X4Y132_SLICE_X4Y132_BQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y157_SLICE_X22Y157_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOI3_X0Y67_ILOGIC_X0Y67_D = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D1 = CLBLL_L_X4Y155_SLICE_X4Y155_CQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D2 = CLBLM_L_X8Y134_SLICE_X10Y134_CO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D3 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D4 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D5 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D6 = CLBLL_L_X4Y131_SLICE_X4Y131_BQ;
  assign CLBLM_L_X16Y157_SLICE_X22Y157_D1 = 1'b1;
  assign CLBLM_L_X16Y157_SLICE_X22Y157_D2 = 1'b1;
  assign CLBLM_L_X16Y157_SLICE_X22Y157_D3 = 1'b1;
  assign CLBLM_L_X16Y157_SLICE_X22Y157_D4 = 1'b1;
  assign CLBLM_L_X16Y157_SLICE_X22Y157_D5 = 1'b1;
  assign CLBLM_L_X16Y157_SLICE_X22Y157_D6 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A1 = CLBLM_R_X7Y132_SLICE_X8Y132_A5Q;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A2 = BRAM_L_X6Y135_RAMB18_X0Y54_DO3;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A3 = BRAM_R_X17Y135_RAMB18_X1Y54_DO4;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A4 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO4;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A5 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO4;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A6 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO3;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B1 = CLBLM_R_X7Y132_SLICE_X8Y132_A5Q;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B2 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B3 = BRAM_L_X6Y135_RAMB18_X0Y54_DO7;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B4 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO7;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B5 = CLBLM_L_X8Y136_SLICE_X11Y136_AO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B6 = CLBLM_L_X16Y151_SLICE_X22Y151_BQ;
  assign RIOB33_X105Y93_IOB_X1Y94_O = CLBLM_L_X10Y131_SLICE_X13Y131_AQ;
  assign RIOB33_X105Y93_IOB_X1Y93_O = CLBLM_L_X12Y132_SLICE_X16Y132_CQ;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C1 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C2 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO5;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C3 = BRAM_R_X17Y135_RAMB18_X1Y54_DO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C4 = BRAM_R_X17Y135_RAMB18_X1Y54_DO5;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C5 = CLBLM_R_X7Y129_SLICE_X9Y129_B5Q;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C6 = BRAM_L_X6Y135_RAMB18_X0Y54_DO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D1 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D2 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D3 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D4 = CLBLM_L_X8Y136_SLICE_X11Y136_CO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D5 = CLBLM_R_X7Y129_SLICE_X9Y129_B5Q;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D6 = CLBLM_R_X25Y149_SLICE_X36Y149_BQ;
  assign RIOI3_X105Y67_OLOGIC_X1Y68_D1 = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A1 = CLBLM_L_X8Y136_SLICE_X10Y136_A5Q;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A2 = BRAM_L_X6Y130_RAMB18_X0Y52_DO4;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A3 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO4;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A4 = LIOB33_X0Y135_IOB_X0Y136_I;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A5 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A6 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B1 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO2;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B2 = BRAM_L_X6Y135_RAMB18_X0Y54_DO2;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B3 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO3;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B4 = BRAM_R_X17Y135_RAMB18_X1Y54_DO3;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B5 = CLBLM_L_X8Y130_SLICE_X10Y130_B5Q;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B6 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO3;
  assign RIOI3_X105Y67_OLOGIC_X1Y68_T1 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C1 = CLBLM_L_X8Y130_SLICE_X10Y130_B5Q;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C2 = BRAM_L_X6Y135_RAMB18_X0Y54_DO7;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C3 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO7;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C4 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C5 = CLBLM_L_X8Y136_SLICE_X10Y136_BO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C6 = CLBLM_L_X16Y151_SLICE_X22Y151_AQ;
  assign RIOI3_X105Y67_OLOGIC_X1Y67_D1 = CLBLM_L_X8Y127_SLICE_X10Y127_BQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_D1 = CLBLL_L_X54Y133_SLICE_X82Y133_AQ;
  assign RIOI3_X105Y67_OLOGIC_X1Y67_T1 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D1 = BRAM_L_X6Y135_RAMB18_X0Y54_DO1;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D2 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO1;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D3 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO0;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D4 = BRAM_R_X17Y135_RAMB18_X1Y54_DO0;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D5 = CLBLM_R_X7Y125_SLICE_X8Y125_B5Q;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D6 = BRAM_R_X17Y135_RAMB18_X1Y54_DO1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_D1 = CLBLM_R_X5Y134_SLICE_X7Y134_BQ;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_T1 = 1'b1;
  assign LIOI3_X0Y145_ILOGIC_X0Y146_D = LIOB33_X0Y145_IOB_X0Y146_I;
  assign LIOI3_X0Y145_ILOGIC_X0Y145_D = LIOB33_X0Y145_IOB_X0Y145_I;
  assign RIOI3_X105Y189_ILOGIC_X1Y190_D = RIOB33_X105Y189_IOB_X1Y190_I;
  assign RIOI3_X105Y189_ILOGIC_X1Y189_D = RIOB33_X105Y189_IOB_X1Y189_I;
  assign LIOI3_X0Y23_ILOGIC_X0Y24_D = LIOB33_X0Y23_IOB_X0Y24_I;
  assign LIOI3_X0Y23_ILOGIC_X0Y23_D = LIOB33_X0Y23_IOB_X0Y23_I;
  assign RIOB33_X105Y95_IOB_X1Y96_O = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign RIOB33_X105Y95_IOB_X1Y95_O = CLBLM_R_X11Y131_SLICE_X14Y131_BQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_A1 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO7;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_A2 = BRAM_L_X6Y135_RAMB18_X0Y54_DO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_A3 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO7;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_A4 = BRAM_R_X17Y135_RAMB18_X1Y54_DO7;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_A5 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_A6 = CLBLM_R_X5Y134_SLICE_X7Y134_A5Q;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_B1 = BRAM_R_X17Y135_RAMB18_X1Y54_DO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_B2 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_B3 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO7;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_B4 = BRAM_R_X17Y135_RAMB18_X1Y54_DO7;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_B5 = BRAM_L_X6Y135_RAMB18_X0Y54_DO7;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_B6 = CLBLM_L_X8Y130_SLICE_X10Y130_A5Q;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_C1 = CLBLM_L_X8Y137_SLICE_X11Y137_AO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_C2 = CLBLM_R_X5Y134_SLICE_X7Y134_A5Q;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_C3 = CLBLM_R_X25Y151_SLICE_X36Y151_CQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_C4 = 1'b1;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_C5 = 1'b1;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_C6 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_D1 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_D2 = CLBLM_L_X16Y149_SLICE_X22Y149_BQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_D3 = 1'b1;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_D4 = CLBLM_L_X8Y130_SLICE_X10Y130_A5Q;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_D5 = 1'b1;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_D6 = CLBLM_L_X8Y137_SLICE_X11Y137_BO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_A1 = BRAM_L_X6Y130_RAMB18_X0Y52_DO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_A2 = CLBLM_L_X8Y137_SLICE_X10Y137_A5Q;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_A3 = LIOB33_X0Y137_IOB_X0Y138_I;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_A4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_A5 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_A6 = 1'b1;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_B1 = CLBLM_L_X8Y137_SLICE_X10Y137_B5Q;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_B2 = LIOB33_X0Y139_IOB_X0Y139_I;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_B3 = BRAM_L_X6Y130_RAMB18_X0Y52_DO7;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_B4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_B5 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO7;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_B6 = 1'b1;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_C1 = BRAM_L_X6Y135_RAMB18_X0Y54_DO0;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_C2 = BRAM_R_X17Y135_RAMB18_X1Y54_DO1;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_C3 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO1;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_C4 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO1;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_C5 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO0;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_C6 = CLBLM_R_X7Y136_SLICE_X8Y136_A5Q;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_D1 = BRAM_L_X6Y135_RAMB18_X0Y54_DO7;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_D2 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_D3 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO7;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_D4 = CLBLM_L_X8Y137_SLICE_X10Y137_CO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_D5 = CLBLM_L_X16Y151_SLICE_X23Y151_AQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_D6 = CLBLM_R_X7Y136_SLICE_X8Y136_A5Q;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_A1 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_A2 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_A3 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_A4 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_A5 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_A6 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_B1 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_B2 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_B3 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_B4 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_B5 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_B6 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_C1 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_C2 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_C3 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_C4 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_C5 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_C6 = 1'b1;
  assign RIOB33_X105Y97_IOB_X1Y98_O = CLBLM_R_X7Y125_SLICE_X8Y125_CQ;
  assign RIOB33_X105Y97_IOB_X1Y97_O = CLBLM_R_X7Y125_SLICE_X8Y125_BQ;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_D1 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_D2 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_D3 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_A1 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_A2 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_A3 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_A4 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_A5 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_A6 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_D4 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_D5 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_B1 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_D6 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_B2 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_B3 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_B4 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_B5 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_B6 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_C1 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_C2 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_C3 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_C4 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_C5 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_C6 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_D1 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_D2 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_D3 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_D4 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_D5 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_D6 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_A1 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_A2 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_A3 = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_A4 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_A5 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_A6 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO3;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_B1 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_B2 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_B3 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_B4 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_B5 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_B6 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_C1 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_C2 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_C3 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_C4 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_C5 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_C6 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_D1 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_D2 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_D3 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_D4 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_D5 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_D6 = 1'b1;
  assign LIOI3_SING_X0Y0_ILOGIC_X0Y0_D = LIOB33_SING_X0Y0_IOB_X0Y0_I;
  assign RIOI3_X105Y71_OLOGIC_X1Y72_D1 = CLBLM_R_X7Y128_SLICE_X9Y128_AQ;
  assign RIOI3_X105Y71_OLOGIC_X1Y72_T1 = 1'b1;
  assign RIOI3_X105Y71_OLOGIC_X1Y71_D1 = CLBLL_L_X54Y101_SLICE_X82Y101_AQ;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_D1 = CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  assign RIOI3_X105Y71_OLOGIC_X1Y71_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_D1 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_T1 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_C5 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_C6 = 1'b1;
  assign RIOB33_X105Y101_IOB_X1Y102_O = CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  assign RIOB33_X105Y101_IOB_X1Y101_O = CLBLM_R_X7Y126_SLICE_X8Y126_AQ;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A1 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A4 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A5 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A6 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B1 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B4 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B5 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B6 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C1 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_D1 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C4 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C5 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_D2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C6 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_D3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D1 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_D4 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D4 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D5 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_D5 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D6 = 1'b1;
  assign LIOI3_X0Y147_ILOGIC_X0Y148_D = LIOB33_X0Y147_IOB_X0Y148_I;
  assign LIOI3_X0Y147_ILOGIC_X0Y147_D = LIOB33_X0Y147_IOB_X0Y147_I;
  assign RIOI3_X105Y191_ILOGIC_X1Y192_D = RIOB33_X105Y191_IOB_X1Y192_I;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A1 = CLBLM_R_X3Y129_SLICE_X2Y129_A5Q;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A2 = CLBLL_L_X2Y131_SLICE_X1Y131_A5Q;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A3 = CLBLM_R_X3Y129_SLICE_X2Y129_BQ;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A4 = CLBLM_R_X3Y129_SLICE_X2Y129_AQ;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A5 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A6 = 1'b1;
  assign RIOI3_X105Y191_ILOGIC_X1Y191_D = RIOB33_X105Y191_IOB_X1Y191_I;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B1 = CLBLM_R_X3Y129_SLICE_X2Y129_A5Q;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B2 = CLBLM_R_X3Y129_SLICE_X2Y129_AQ;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B3 = CLBLM_R_X3Y129_SLICE_X2Y129_BQ;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B4 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B5 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B6 = 1'b1;
  assign LIOI3_X0Y25_ILOGIC_X0Y26_D = LIOB33_X0Y25_IOB_X0Y26_I;
  assign LIOI3_X0Y25_ILOGIC_X0Y25_D = LIOB33_X0Y25_IOB_X0Y25_I;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C1 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C4 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C5 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C6 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D1 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D4 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D5 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D6 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_SR = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_A5 = LIOB33_X0Y71_IOB_X0Y71_I;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_A6 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_B1 = LIOB33_X0Y21_IOB_X0Y21_I;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_B2 = CLBLL_L_X4Y128_SLICE_X5Y128_BQ;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_B3 = CLBLL_L_X4Y128_SLICE_X5Y128_AQ;
  assign RIOB33_X105Y103_IOB_X1Y103_O = CLBLM_R_X7Y126_SLICE_X8Y126_CQ;
  assign RIOB33_X105Y103_IOB_X1Y104_O = CLBLM_R_X7Y128_SLICE_X8Y128_BQ;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_B4 = CLBLM_L_X8Y130_SLICE_X10Y130_A5Q;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_B5 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_B6 = BRAM_L_X6Y125_RAMB18_X0Y50_DO7;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_C1 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_C2 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_C3 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_A1 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_A2 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_A3 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_A4 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_A5 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_A6 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_B1 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_B2 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_B3 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_B4 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_B5 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_B6 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_C1 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_C2 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_C3 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_C4 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_C5 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_C6 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_D1 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_D2 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_D3 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_D4 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_D5 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_D6 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_A1 = CLBLM_R_X3Y132_SLICE_X2Y132_CQ;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_A2 = CLBLM_R_X3Y132_SLICE_X2Y132_AO5;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_A3 = CLBLL_L_X2Y132_SLICE_X1Y132_AQ;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_A4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_A5 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_B1 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_B2 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_B3 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_B4 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_B5 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_B6 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_C1 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_C2 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_C3 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_C4 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_C5 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_C6 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_D1 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_D2 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_D3 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_D4 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_D5 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_D6 = 1'b1;
  assign RIOB33_X105Y105_IOB_X1Y106_O = CLBLM_R_X5Y131_SLICE_X7Y131_AQ;
  assign RIOB33_X105Y105_IOB_X1Y105_O = CLBLM_R_X7Y129_SLICE_X9Y129_CQ;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_D = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign RIOI3_X105Y73_OLOGIC_X1Y74_D1 = CLBLM_R_X7Y130_SLICE_X9Y130_DQ;
  assign RIOI3_X105Y73_OLOGIC_X1Y74_T1 = 1'b1;
  assign RIOI3_X105Y73_OLOGIC_X1Y73_D1 = CLBLM_L_X8Y130_SLICE_X11Y130_BQ;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1 = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign RIOI3_X105Y73_OLOGIC_X1Y73_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1 = CLBLM_L_X8Y130_SLICE_X10Y130_BQ;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1 = 1'b1;
  assign RIOI3_SING_X105Y200_ILOGIC_X1Y200_D = RIOB33_SING_X105Y200_IOB_X1Y200_I;
  assign LIOI3_X0Y151_ILOGIC_X0Y152_D = LIOB33_X0Y151_IOB_X0Y152_I;
  assign LIOI3_X0Y151_ILOGIC_X0Y151_D = LIOB33_X0Y151_IOB_X0Y151_I;
  assign RIOI3_X105Y195_ILOGIC_X1Y196_D = RIOB33_X105Y195_IOB_X1Y196_I;
  assign RIOI3_X105Y195_ILOGIC_X1Y195_D = RIOB33_X105Y195_IOB_X1Y195_I;
  assign RIOB33_X105Y107_IOB_X1Y108_O = CLBLM_R_X7Y130_SLICE_X8Y130_BQ;
  assign RIOB33_X105Y107_IOB_X1Y107_O = CLBLL_L_X54Y119_SLICE_X82Y119_AQ;
  assign LIOI3_X0Y27_ILOGIC_X0Y28_D = LIOB33_X0Y27_IOB_X0Y28_I;
  assign LIOI3_X0Y27_ILOGIC_X0Y27_D = LIOB33_X0Y27_IOB_X0Y27_I;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A1 = LIOB33_X0Y65_IOB_X0Y65_I;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A2 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A3 = CLBLM_R_X5Y125_SLICE_X7Y125_AQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A4 = BRAM_L_X6Y125_RAMB18_X0Y50_DO1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A5 = CLBLM_R_X7Y125_SLICE_X8Y125_B5Q;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A6 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B1 = BRAM_L_X6Y125_RAMB18_X0Y50_DO2;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B2 = CLBLM_R_X5Y125_SLICE_X7Y125_BQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B3 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B5 = CLBLM_R_X7Y125_SLICE_X8Y125_C5Q;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B6 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C1 = BRAM_L_X6Y125_RAMB18_X0Y50_DO1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C2 = CLBLM_R_X5Y125_SLICE_X7Y125_CQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C3 = CLBLM_R_X7Y125_SLICE_X8Y125_B5Q;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C4 = CLBLM_R_X5Y125_SLICE_X7Y125_AQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C5 = LIOB33_X0Y51_IOB_X0Y51_I;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C6 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D1 = CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D2 = LIOB33_X0Y1_IOB_X0Y2_I;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D3 = CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D4 = BRAM_L_X6Y125_RAMB18_X0Y50_DO2;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D5 = CLBLM_R_X5Y125_SLICE_X7Y125_BO5;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D6 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A1 = BRAM_L_X6Y125_RAMB18_X0Y50_DO2;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A2 = CLBLM_R_X7Y125_SLICE_X8Y125_C5Q;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A3 = CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A4 = CLBLM_R_X5Y125_SLICE_X7Y125_BQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A5 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A6 = LIOB33_X0Y17_IOB_X0Y17_I;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B1 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B2 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B3 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B4 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B5 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B6 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C1 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C2 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C3 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C4 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C5 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C6 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D1 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D2 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D3 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D4 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D5 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D6 = 1'b1;
  assign LIOI3_SING_X0Y99_ILOGIC_X0Y99_D = LIOB33_SING_X0Y99_IOB_X0Y99_I;
  assign RIOB33_X105Y109_IOB_X1Y110_O = CLBLM_R_X7Y129_SLICE_X8Y129_DQ;
  assign RIOB33_X105Y109_IOB_X1Y109_O = CLBLM_R_X7Y129_SLICE_X8Y129_CQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A1 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A2 = CLBLM_R_X7Y129_SLICE_X9Y129_A5Q;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A3 = CLBLM_R_X5Y126_SLICE_X7Y126_AQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A5 = BRAM_L_X6Y125_RAMB18_X0Y50_DO4;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A6 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B1 = CLBLM_R_X7Y129_SLICE_X9Y129_A5Q;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B2 = CLBLM_R_X5Y126_SLICE_X7Y126_BQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B3 = CLBLM_R_X5Y126_SLICE_X7Y126_AQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B5 = BRAM_L_X6Y125_RAMB18_X0Y50_DO4;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B6 = LIOB33_X0Y17_IOB_X0Y18_I;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_BX = CLBLM_R_X5Y126_SLICE_X6Y126_CO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C1 = BRAM_L_X6Y125_RAMB18_X0Y50_DO4;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C2 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C3 = CLBLM_R_X5Y126_SLICE_X7Y126_BQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C4 = CLBLM_R_X5Y126_SLICE_X7Y126_AO5;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C5 = LIOB33_X0Y3_IOB_X0Y4_I;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C6 = CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D1 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D2 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D3 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D4 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D5 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D6 = 1'b1;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1 = CLBLL_L_X2Y141_SLICE_X0Y141_AQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A1 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A2 = BRAM_L_X6Y125_RAMB18_X0Y50_DO3;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A3 = CLBLM_R_X5Y126_SLICE_X6Y126_AQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A5 = CLBLM_R_X7Y126_SLICE_X8Y126_D5Q;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A6 = 1'b1;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B1 = LIOB33_X0Y51_IOB_X0Y52_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B2 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B3 = CLBLM_R_X5Y126_SLICE_X6Y126_AQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B4 = CLBLM_R_X7Y126_SLICE_X8Y126_D5Q;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B5 = CLBLM_R_X5Y126_SLICE_X6Y126_BQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B6 = BRAM_L_X6Y125_RAMB18_X0Y50_DO3;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C1 = CLBLM_R_X5Y126_SLICE_X6Y126_BQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C2 = BRAM_L_X6Y125_RAMB18_X0Y50_DO3;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C3 = CLBLM_R_X5Y126_SLICE_X7Y126_B5Q;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C4 = CLBLM_R_X5Y126_SLICE_X6Y126_AO5;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C5 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C6 = LIOB33_X0Y3_IOB_X0Y3_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D1 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D2 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D3 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D4 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D5 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D6 = 1'b1;
  assign RIOI3_X105Y179_ILOGIC_X1Y180_D = RIOB33_X105Y179_IOB_X1Y180_I;
  assign RIOI3_X105Y75_OLOGIC_X1Y76_D1 = CLBLM_L_X10Y132_SLICE_X12Y132_AQ;
  assign RIOB33_X105Y111_IOB_X1Y112_O = CLBLM_R_X7Y131_SLICE_X9Y131_BQ;
  assign RIOB33_X105Y111_IOB_X1Y111_O = CLBLM_R_X7Y130_SLICE_X9Y130_AQ;
  assign RIOI3_X105Y75_OLOGIC_X1Y76_T1 = 1'b1;
  assign RIOI3_X105Y179_ILOGIC_X1Y179_D = RIOB33_X105Y179_IOB_X1Y179_I;
  assign RIOI3_X105Y75_OLOGIC_X1Y75_D1 = CLBLM_L_X8Y130_SLICE_X10Y130_DQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A1 = CLBLM_R_X5Y126_SLICE_X7Y126_BQ;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1 = CLBLM_L_X56Y151_SLICE_X84Y151_AQ;
  assign RIOI3_X105Y75_OLOGIC_X1Y75_T1 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B6 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_ADDRARDADDR0 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_ADDRARDADDR1 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_ADDRARDADDR2 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_ADDRARDADDR3 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_ADDRARDADDR4 = CLBLM_R_X3Y130_SLICE_X3Y130_CO6;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_ADDRARDADDR5 = CLBLL_L_X4Y132_SLICE_X5Y132_DO6;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_ADDRARDADDR6 = CLBLL_L_X4Y130_SLICE_X5Y130_DO6;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_ADDRARDADDR7 = CLBLM_R_X5Y129_SLICE_X6Y129_DO6;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_ADDRARDADDR8 = CLBLL_L_X4Y133_SLICE_X5Y133_DO6;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_ADDRARDADDR9 = CLBLL_L_X4Y133_SLICE_X4Y133_CO6;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_ADDRARDADDR10 = CLBLL_L_X4Y132_SLICE_X5Y132_CO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A2 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_ADDRARDADDR11 = CLBLL_L_X4Y132_SLICE_X5Y132_BO6;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_ADDRARDADDR12 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_ADDRARDADDR13 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_ADDRATIEHIGH0 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_ADDRATIEHIGH1 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_ADDRBTIEHIGH0 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_ADDRBTIEHIGH1 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_ADDRBWRADDR0 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_ADDRBWRADDR1 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_ADDRBWRADDR2 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_ADDRBWRADDR3 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_ADDRBWRADDR4 = CLBLM_R_X5Y127_SLICE_X6Y127_DO6;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_ADDRBWRADDR5 = CLBLM_R_X7Y125_SLICE_X8Y125_DO6;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_ADDRBWRADDR6 = CLBLM_R_X5Y125_SLICE_X7Y125_DO6;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_ADDRBWRADDR7 = CLBLM_R_X5Y126_SLICE_X6Y126_CO6;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_ADDRBWRADDR8 = CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_ADDRBWRADDR9 = CLBLM_R_X5Y127_SLICE_X7Y127_DO6;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_ADDRBWRADDR10 = CLBLM_R_X5Y127_SLICE_X7Y127_CO6;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_ADDRBWRADDR11 = CLBLL_L_X4Y127_SLICE_X5Y127_BO6;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_ADDRBWRADDR12 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_ADDRBWRADDR13 = 1'b0;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C2 = CLBLM_R_X5Y131_SLICE_X6Y131_CQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C1 = BRAM_L_X6Y130_RAMB18_X0Y52_DO0;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A3 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_RDCLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_WRCLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C3 = CLBLM_L_X8Y132_SLICE_X11Y132_A5Q;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_DIADI0 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_DIADI1 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_DIADI2 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_DIADI3 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_DIADI4 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_DIADI5 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_DIADI6 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_DIADI7 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C5 = LIOB33_X0Y29_IOB_X0Y30_I;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_DIADI8 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_DIADI9 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_DIADI10 = 1'b0;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A1 = CLBLM_R_X7Y128_SLICE_X8Y128_A5Q;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C6 = CLBLM_R_X5Y131_SLICE_X7Y131_A5Q;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A2 = BRAM_L_X6Y125_RAMB18_X0Y50_DO5;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A3 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A5 = LIOB33_X0Y69_IOB_X0Y69_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A6 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_DIBDI0 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A4 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO4;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B1 = CLBLM_R_X7Y128_SLICE_X8Y128_A5Q;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_DIBDI4 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_DIBDI5 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_DIBDI6 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_DIBDI7 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_DIBDI8 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_DIBDI9 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_DIBDI10 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_DIBDI11 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_DIBDI12 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_DIBDI13 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_DIBDI15 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_DIPADIP0 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_DIPADIP1 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_DIPBDIP0 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_DIPBDIP1 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_BX = CLBLM_R_X5Y127_SLICE_X7Y127_DO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C1 = BRAM_L_X6Y125_RAMB18_X0Y50_DO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C2 = CLBLM_R_X5Y127_SLICE_X7Y127_CQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C3 = LIOB33_X0Y5_IOB_X0Y6_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C5 = CLBLM_R_X5Y127_SLICE_X6Y127_AO5;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C6 = CLBLL_L_X4Y127_SLICE_X5Y127_AQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A5 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D1 = CLBLM_R_X5Y127_SLICE_X7Y127_BQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D2 = BRAM_L_X6Y125_RAMB18_X0Y50_DO5;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D3 = LIOB33_X0Y5_IOB_X0Y5_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D4 = CLBLM_R_X5Y127_SLICE_X7Y127_AO5;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D5 = CLBLM_R_X5Y127_SLICE_X7Y127_B5Q;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D6 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_DX = CLBLL_L_X4Y127_SLICE_X5Y127_BO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A1 = CLBLM_R_X7Y129_SLICE_X9Y129_B5Q;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A2 = CLBLM_R_X5Y127_SLICE_X6Y127_B5Q;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A3 = BRAM_L_X6Y125_RAMB18_X0Y50_DO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A5 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A6 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_RDEN = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D1 = BRAM_L_X6Y130_RAMB18_X0Y52_DO4;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_WREN = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_AX = CLBLM_R_X5Y127_SLICE_X6Y127_CO5;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B2 = CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B3 = CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B5 = BRAM_L_X6Y125_RAMB18_X0Y50_DO0;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B6 = CLBLM_R_X7Y127_SLICE_X8Y127_A5Q;
  assign LIOI3_X0Y153_ILOGIC_X0Y154_D = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D3 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO5;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A6 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_BX = CLBLM_R_X5Y127_SLICE_X6Y127_AO6;
  assign LIOI3_X0Y153_ILOGIC_X0Y153_D = LIOB33_X0Y153_IOB_X0Y153_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C1 = BRAM_L_X6Y125_RAMB18_X0Y50_DO0;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D4 = CLBLM_R_X5Y131_SLICE_X7Y131_CQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C2 = LIOB33_X0Y63_IOB_X0Y64_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C3 = CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C5 = CLBLM_R_X7Y127_SLICE_X8Y127_A5Q;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C6 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_REGCE = 1'b0;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_REGCEB = 1'b0;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D6 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_RDRCLK = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_REGCLKB = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_RST = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_RSTRAMB = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_RSTREG = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_RSTREGB = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_WEA0 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_WEA1 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_WEA2 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_WEA3 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_WEBWE0 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_WEBWE1 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_WEBWE2 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_WEBWE3 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_WEBWE4 = 1'b0;
  assign LIOI3_X0Y29_ILOGIC_X0Y30_D = LIOB33_X0Y29_IOB_X0Y30_I;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_WEBWE6 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_WEBWE7 = 1'b0;
  assign LIOI3_X0Y29_ILOGIC_X0Y29_D = LIOB33_X0Y29_IOB_X0Y29_I;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C1 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D3 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C2 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D6 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C3 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C4 = 1'b1;
  assign LIOI3_SING_X0Y149_ILOGIC_X0Y149_D = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_ILOGIC_X0Y143_D = LIOB33_X0Y143_IOB_X0Y143_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A1 = LIOB33_X0Y73_IOB_X0Y74_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A2 = BRAM_L_X6Y125_RAMB18_X0Y50_DO18;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A6 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A1 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A2 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A3 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A4 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A5 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A6 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_AX = CLBLM_R_X5Y129_SLICE_X7Y129_AO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B1 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B2 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B3 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B4 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B5 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B6 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C1 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C2 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C3 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C4 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C5 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C6 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D1 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D2 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D3 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D4 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D5 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D6 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A2 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A3 = CLBLM_R_X5Y128_SLICE_X6Y128_AQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A4 = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A5 = BRAM_L_X6Y125_RAMB18_X0Y50_DO19;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A6 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B1 = CLBLM_L_X8Y130_SLICE_X10Y130_B5Q;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B2 = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B3 = CLBLM_R_X5Y128_SLICE_X6Y128_AQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B5 = BRAM_L_X6Y125_RAMB18_X0Y50_DO19;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B6 = LIOB33_X0Y25_IOB_X0Y25_I;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C1 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C2 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C3 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C4 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C5 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C6 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D1 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D2 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D3 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D4 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D5 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D6 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A4 = CLBLM_R_X7Y133_SLICE_X8Y133_BO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C1 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO7;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A5 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C2 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO7;
  assign RIOB33_X105Y115_IOB_X1Y116_O = CLBLM_L_X10Y133_SLICE_X13Y133_AQ;
  assign RIOB33_X105Y115_IOB_X1Y115_O = CLBLL_L_X54Y123_SLICE_X82Y123_AQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C3 = CLBLM_R_X5Y129_SLICE_X6Y129_A5Q;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C4 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign LIOI3_SING_X0Y150_ILOGIC_X0Y150_D = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B1 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO3;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A1 = CLBLM_R_X7Y129_SLICE_X8Y129_A5Q;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A2 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A3 = LIOB33_X0Y71_IOB_X0Y72_I;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A4 = BRAM_L_X6Y125_RAMB18_X0Y50_DO16;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A5 = CLBLM_R_X5Y128_SLICE_X7Y128_AQ;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A6 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_AX = CLBLM_R_X5Y129_SLICE_X6Y129_DO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B1 = LIOB33_X0Y21_IOB_X0Y22_I;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B2 = CLBLM_R_X5Y129_SLICE_X7Y129_BQ;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B3 = CLBLM_R_X5Y128_SLICE_X7Y128_AQ;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B5 = BRAM_L_X6Y125_RAMB18_X0Y50_DO16;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B6 = CLBLM_R_X7Y129_SLICE_X8Y129_A5Q;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_BX = CLBLM_R_X5Y129_SLICE_X7Y129_CO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C1 = BRAM_L_X6Y125_RAMB18_X0Y50_DO17;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C2 = CLBLM_R_X5Y129_SLICE_X6Y129_BQ;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C3 = LIOB33_X0Y7_IOB_X0Y8_I;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C4 = CLBLL_L_X4Y129_SLICE_X5Y129_BO5;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C5 = CLBLM_R_X5Y129_SLICE_X7Y129_B5Q;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C6 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign RIOI3_X105Y77_OLOGIC_X1Y78_D1 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y77_OLOGIC_X1Y78_T1 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D1 = BRAM_L_X6Y125_RAMB18_X0Y50_DO16;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D2 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D3 = CLBLM_R_X5Y129_SLICE_X7Y129_BQ;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D4 = CLBLM_R_X5Y129_SLICE_X7Y129_AO5;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D5 = LIOB33_X0Y7_IOB_X0Y7_I;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D6 = CLBLM_R_X5Y130_SLICE_X7Y130_CQ;
  assign RIOI3_X105Y77_OLOGIC_X1Y77_D1 = CLBLM_L_X8Y130_SLICE_X11Y130_CQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A1 = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A2 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A3 = CLBLM_R_X5Y129_SLICE_X6Y129_AQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A4 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A5 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A6 = CLBLM_R_X5Y130_SLICE_X6Y130_AO5;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_AX = CLBLM_R_X5Y129_SLICE_X6Y129_CO6;
  assign RIOI3_X105Y77_OLOGIC_X1Y77_T1 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B1 = CLBLM_R_X7Y136_SLICE_X8Y136_A5Q;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B2 = CLBLM_R_X5Y129_SLICE_X6Y129_BQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B3 = BRAM_L_X6Y125_RAMB18_X0Y50_DO17;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B5 = LIOB33_X0Y23_IOB_X0Y23_I;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B6 = CLBLL_L_X4Y129_SLICE_X4Y129_AQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C1 = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C2 = CLBLM_R_X5Y128_SLICE_X6Y128_AO5;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C3 = LIOB33_X0Y9_IOB_X0Y10_I;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C4 = CLBLM_R_X5Y129_SLICE_X6Y129_A5Q;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C5 = BRAM_L_X6Y125_RAMB18_X0Y50_DO19;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C6 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D1 = CLBLM_R_X5Y129_SLICE_X7Y129_AQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D2 = CLBLM_R_X5Y129_SLICE_X6Y129_AQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D3 = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D4 = CLBLM_R_X5Y130_SLICE_X6Y130_AO5;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D5 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign RIOB33_X105Y117_IOB_X1Y118_O = CLBLM_L_X10Y131_SLICE_X12Y131_AQ;
  assign RIOB33_X105Y117_IOB_X1Y117_O = CLBLM_L_X12Y132_SLICE_X16Y132_AQ;
  assign LIOI3_X0Y155_ILOGIC_X0Y156_D = LIOB33_X0Y155_IOB_X0Y156_I;
  assign LIOI3_X0Y155_ILOGIC_X0Y155_D = LIOB33_X0Y155_IOB_X0Y155_I;
  assign RIOI3_X105Y201_ILOGIC_X1Y202_D = RIOB33_X105Y201_IOB_X1Y202_I;
  assign RIOI3_X105Y201_ILOGIC_X1Y201_D = RIOB33_X105Y201_IOB_X1Y201_I;
  assign RIOI3_X105Y205_ILOGIC_X1Y205_D = RIOB33_X105Y205_IOB_X1Y205_I;
  assign RIOI3_TBYTESRC_X105Y181_ILOGIC_X1Y182_D = RIOB33_X105Y181_IOB_X1Y182_I;
  assign RIOI3_TBYTESRC_X105Y181_ILOGIC_X1Y181_D = RIOB33_X105Y181_IOB_X1Y181_I;
  assign LIOI3_SING_X0Y199_ILOGIC_X0Y199_D = LIOB33_SING_X0Y199_IOB_X0Y199_I;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A1 = CLBLL_L_X4Y131_SLICE_X4Y131_DQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A2 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO2;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A3 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A4 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A5 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A6 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_AX = CLBLM_R_X5Y130_SLICE_X6Y130_DO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B1 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B2 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B3 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B4 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B5 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B6 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_BX = CLBLM_R_X3Y130_SLICE_X3Y130_CO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C1 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C2 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C3 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C4 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C5 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C6 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_CX = CLBLM_R_X5Y129_SLICE_X7Y129_DO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D1 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D2 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D3 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D4 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D5 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D6 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A1 = LIOB33_X0Y143_IOB_X0Y143_I;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A2 = BRAM_L_X6Y130_RAMB18_X0Y52_DO19;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A3 = CLBLM_R_X5Y130_SLICE_X6Y130_AQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A5 = CLBLM_R_X3Y131_SLICE_X2Y131_B5Q;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A6 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B1 = CLBLM_R_X5Y130_SLICE_X6Y130_AQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B2 = BRAM_L_X6Y130_RAMB18_X0Y52_DO19;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B3 = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B5 = LIOB33_X0Y91_IOB_X0Y91_I;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B6 = CLBLM_R_X3Y131_SLICE_X2Y131_B5Q;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1 = CLBLM_R_X7Y134_SLICE_X9Y134_AQ;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_D1 = CLBLL_L_X54Y119_SLICE_X82Y119_AQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_BX = CLBLL_L_X4Y130_SLICE_X5Y130_CO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C1 = LIOB33_X0Y15_IOB_X0Y15_I;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C2 = CLBLM_R_X5Y130_SLICE_X6Y130_CQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C3 = CLBLM_R_X5Y131_SLICE_X6Y131_BO5;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C4 = CLBLM_R_X5Y131_SLICE_X6Y131_CQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C5 = BRAM_L_X6Y130_RAMB18_X0Y52_DO0;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C6 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D1 = BRAM_L_X6Y125_RAMB18_X0Y50_DO20;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D2 = CLBLM_R_X5Y130_SLICE_X7Y130_A5Q;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D3 = LIOB33_X0Y11_IOB_X0Y11_I;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D4 = CLBLL_L_X4Y131_SLICE_X4Y131_AO5;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D5 = CLBLL_L_X4Y131_SLICE_X5Y131_BQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D6 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_DX = CLBLL_L_X4Y130_SLICE_X4Y130_CO6;
  assign RIOB33_X105Y119_IOB_X1Y120_O = CLBLM_L_X10Y133_SLICE_X13Y133_BQ;
  assign RIOB33_X105Y119_IOB_X1Y119_O = CLBLM_R_X11Y133_SLICE_X14Y133_AQ;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_T1 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A1 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A2 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A3 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A4 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A5 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A6 = CLBLM_R_X5Y127_SLICE_X7Y127_CQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_AX = CLBLM_R_X5Y131_SLICE_X6Y131_BO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B1 = CLBLM_L_X8Y136_SLICE_X10Y136_A5Q;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B2 = CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B3 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B5 = BRAM_L_X6Y130_RAMB18_X0Y52_DO4;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B6 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C1 = BRAM_L_X6Y130_RAMB18_X0Y52_DO4;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C2 = CLBLM_R_X5Y131_SLICE_X7Y131_CQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C3 = CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C4 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C5 = CLBLM_L_X8Y136_SLICE_X10Y136_A5Q;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C6 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign LIOI3_SING_X0Y200_ILOGIC_X0Y200_D = LIOB33_SING_X0Y200_IOB_X0Y200_I;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D1 = BRAM_L_X6Y135_RAMB18_X0Y54_DO23;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D2 = BRAM_R_X17Y135_RAMB18_X1Y54_DO22;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D3 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO7;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D4 = CLBLL_L_X4Y128_SLICE_X5Y128_AQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D5 = BRAM_R_X17Y135_RAMB18_X1Y54_DO23;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D6 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A1 = CLBLM_R_X5Y129_SLICE_X6Y129_AQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A2 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A3 = BRAM_L_X6Y140_RAMB18_X0Y56_DO3;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A4 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A5 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A6 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_AX = CLBLM_R_X5Y131_SLICE_X6Y131_DO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B1 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B2 = CLBLM_L_X8Y132_SLICE_X11Y132_A5Q;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B3 = CLBLM_R_X5Y131_SLICE_X7Y131_A5Q;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B5 = BRAM_L_X6Y130_RAMB18_X0Y52_DO0;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_ADDRARDADDR0 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_ADDRARDADDR1 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_ADDRARDADDR2 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_ADDRARDADDR3 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_ADDRARDADDR4 = CLBLM_R_X7Y136_SLICE_X8Y136_DO6;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_ADDRARDADDR5 = CLBLM_R_X7Y136_SLICE_X8Y136_CO6;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_ADDRARDADDR6 = CLBLM_R_X7Y134_SLICE_X8Y134_DO6;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_ADDRARDADDR7 = CLBLM_R_X7Y134_SLICE_X8Y134_CO6;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_ADDRARDADDR8 = CLBLM_L_X10Y134_SLICE_X13Y134_BO6;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_ADDRARDADDR9 = CLBLM_L_X10Y137_SLICE_X12Y137_DO6;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_ADDRARDADDR10 = CLBLM_L_X8Y136_SLICE_X11Y136_DO6;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_ADDRARDADDR11 = CLBLM_L_X8Y137_SLICE_X11Y137_DO6;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_ADDRARDADDR12 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_ADDRARDADDR13 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_ADDRATIEHIGH0 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_ADDRATIEHIGH1 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_ADDRBTIEHIGH0 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_ADDRBTIEHIGH1 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_ADDRBWRADDR0 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_ADDRBWRADDR1 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_ADDRBWRADDR2 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_ADDRBWRADDR3 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_ADDRBWRADDR4 = CLBLM_R_X7Y132_SLICE_X8Y132_DO6;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_ADDRBWRADDR5 = CLBLM_R_X7Y131_SLICE_X8Y131_DO6;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_ADDRBWRADDR6 = CLBLM_R_X7Y130_SLICE_X8Y130_DO6;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_ADDRBWRADDR7 = CLBLM_R_X7Y131_SLICE_X8Y131_CO6;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_ADDRBWRADDR8 = CLBLM_R_X7Y132_SLICE_X8Y132_CO6;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_ADDRBWRADDR9 = CLBLM_R_X7Y133_SLICE_X8Y133_DO6;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_ADDRBWRADDR10 = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_ADDRBWRADDR11 = CLBLL_L_X4Y131_SLICE_X5Y131_DO6;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_ADDRBWRADDR12 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_ADDRBWRADDR13 = 1'b0;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D2 = CLBLM_R_X5Y131_SLICE_X6Y131_A5Q;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D3 = CLBLM_R_X5Y131_SLICE_X7Y131_BO5;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_CLKARDCLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_CLKBWRCLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_DIADI0 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_DIADI1 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_DIADI2 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_DIADI3 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_DIADI4 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_DIADI5 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_DIADI6 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_DIADI7 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_DIADI8 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_DIADI9 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_DIADI10 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_DIADI11 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_DIADI12 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_DIADI13 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_DIADI14 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_DIADI15 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_DIBDI0 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_DIBDI1 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_DIBDI2 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_DIBDI3 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_DIBDI4 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_DIBDI5 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_DIBDI6 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_DIBDI7 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_DIBDI8 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_DIBDI9 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_DIBDI10 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_DIBDI11 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_DIBDI12 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_DIBDI13 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_DIBDI14 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_DIBDI15 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_DIPADIP0 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_DIPADIP1 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_DIPBDIP0 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_DIPBDIP1 = 1'b1;
  assign RIOI3_X105Y79_OLOGIC_X1Y80_D1 = CLBLM_L_X8Y131_SLICE_X11Y131_BQ;
  assign RIOI3_X105Y79_OLOGIC_X1Y80_T1 = 1'b1;
  assign RIOI3_X105Y79_OLOGIC_X1Y79_D1 = CLBLL_L_X54Y105_SLICE_X82Y105_AQ;
  assign RIOI3_X105Y79_OLOGIC_X1Y79_T1 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_ENARDEN = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_ENBWREN = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_REGCEAREGCE = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_REGCEB = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_REGCLKARDRCLK = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_REGCLKB = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_RSTRAMARSTRAM = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_RSTRAMB = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_RSTREGARSTREG = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_RSTREGB = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_WEA0 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_WEA1 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_WEA2 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_WEA3 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_WEBWE0 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_WEBWE1 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_WEBWE2 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_WEBWE3 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_WEBWE4 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_WEBWE5 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_WEBWE6 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y51_WEBWE7 = 1'b0;
  assign LIOI3_X0Y159_ILOGIC_X0Y160_D = LIOB33_X0Y159_IOB_X0Y160_I;
  assign LIOI3_X0Y159_ILOGIC_X0Y159_D = LIOB33_X0Y159_IOB_X0Y159_I;
  assign RIOI3_X105Y203_ILOGIC_X1Y204_D = RIOB33_X105Y203_IOB_X1Y204_I;
  assign RIOI3_X105Y203_ILOGIC_X1Y203_D = RIOB33_X105Y203_IOB_X1Y203_I;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A1 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A2 = CLBLM_R_X5Y132_SLICE_X6Y132_B5Q;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A3 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A4 = BRAM_L_X6Y140_RAMB18_X0Y56_DO17;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A5 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A6 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_AX = CLBLL_L_X4Y132_SLICE_X4Y132_DO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B1 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B2 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B3 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B4 = CLBLM_R_X5Y132_SLICE_X6Y132_BQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B5 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B6 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO3;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_BX = CLBLL_L_X4Y132_SLICE_X5Y132_CO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C1 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO5;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C2 = BRAM_R_X17Y135_RAMB18_X1Y54_DO22;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C3 = CLBLM_R_X5Y127_SLICE_X6Y127_B5Q;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C4 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C5 = BRAM_L_X6Y135_RAMB18_X0Y54_DO22;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C6 = BRAM_R_X17Y135_RAMB18_X1Y54_DO21;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D1 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D2 = CLBLM_R_X3Y157_SLICE_X3Y157_CQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D3 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D4 = CLBLM_R_X5Y132_SLICE_X7Y132_CO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D5 = CLBLM_R_X5Y127_SLICE_X6Y127_B5Q;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D6 = 1'b1;
  assign RIOB33_X105Y123_IOB_X1Y124_O = CLBLM_R_X7Y130_SLICE_X9Y130_BQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A1 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A2 = BRAM_L_X6Y130_RAMB18_X0Y52_DO5;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A3 = CLBLM_R_X5Y132_SLICE_X6Y132_AQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A4 = CLBLM_L_X10Y135_SLICE_X12Y135_A5Q;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A5 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A6 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_A1 = CLBLL_L_X2Y142_SLICE_X0Y142_DQ;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_A2 = CLBLL_L_X2Y142_SLICE_X0Y142_BQ;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_A3 = CLBLL_L_X2Y142_SLICE_X0Y142_AQ;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_A4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B1 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B2 = CLBLM_R_X5Y132_SLICE_X6Y132_BQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B4 = CLBLM_R_X5Y133_SLICE_X6Y133_AQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B5 = CLBLM_R_X7Y134_SLICE_X9Y134_B5Q;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B6 = BRAM_L_X6Y130_RAMB18_X0Y52_DO3;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_B1 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_B2 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_BX = CLBLL_L_X4Y132_SLICE_X5Y132_DO6;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_B3 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C1 = BRAM_L_X6Y130_RAMB18_X0Y52_DO5;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C2 = CLBLM_R_X7Y132_SLICE_X8Y132_CQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C4 = CLBLM_R_X5Y132_SLICE_X6Y132_AO5;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C5 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C6 = CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_C1 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_C2 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_C3 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_C4 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_C5 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_C6 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_D1 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_D2 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_D3 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_D4 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_D5 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_D6 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D1 = CLBLM_R_X5Y132_SLICE_X6Y132_BQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D2 = CLBLM_R_X7Y132_SLICE_X8Y132_BQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D3 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D4 = BRAM_L_X6Y130_RAMB18_X0Y52_DO3;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D5 = CLBLM_R_X5Y133_SLICE_X6Y133_AO5;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D2 = CLBLL_L_X4Y130_SLICE_X5Y130_A5Q;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D3 = LIOB33_X0Y11_IOB_X0Y12_I;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_A1 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_A2 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_A3 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_A4 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_A5 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_A6 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_B1 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_B2 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_B3 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_B4 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_B5 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_B6 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_C1 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_C2 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_C3 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_C4 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_C5 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_C6 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_D1 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_D2 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_D3 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_D4 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_D5 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_D6 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A3 = CLBLL_L_X4Y130_SLICE_X5Y130_AQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A5 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A6 = CLBLM_R_X3Y131_SLICE_X3Y131_AO5;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_AX = CLBLL_L_X4Y130_SLICE_X4Y130_DO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A1 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A2 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A3 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A4 = BRAM_L_X6Y140_RAMB18_X0Y56_DO19;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A5 = CLBLM_R_X5Y129_SLICE_X7Y129_AQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A6 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B1 = CLBLL_L_X4Y130_SLICE_X4Y130_AO5;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B2 = BRAM_L_X6Y130_RAMB18_X0Y52_DO1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B1 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B2 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO2;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B3 = CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B4 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B5 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B6 = 1'b1;
  assign RIOB33_X105Y125_IOB_X1Y126_O = CLBLM_R_X7Y130_SLICE_X9Y130_CQ;
  assign RIOB33_X105Y125_IOB_X1Y125_O = CLBLM_R_X5Y132_SLICE_X7Y132_AQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C1 = CLBLM_R_X3Y130_SLICE_X2Y130_AQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C2 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C3 = BRAM_L_X6Y140_RAMB18_X0Y56_DO0;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C4 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C5 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C6 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D1 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D2 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D3 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO0;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D4 = BRAM_L_X6Y140_RAMB18_X0Y56_DO17;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D5 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO0;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D6 = CLBLM_R_X7Y130_SLICE_X8Y130_B5Q;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_A1 = CLBLL_L_X2Y142_SLICE_X0Y142_CQ;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_A2 = CLBLL_L_X2Y142_SLICE_X0Y142_BQ;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_A3 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_A4 = CLBLL_L_X2Y142_SLICE_X0Y142_AQ;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_A5 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_A6 = CLBLL_L_X2Y142_SLICE_X0Y142_DQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A4 = CLBLM_R_X7Y134_SLICE_X9Y134_B5Q;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A5 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A1 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_B1 = CLBLL_L_X2Y142_SLICE_X0Y142_CQ;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_B2 = CLBLL_L_X2Y142_SLICE_X0Y142_BQ;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_B3 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_B4 = CLBLL_L_X2Y142_SLICE_X0Y142_AQ;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_B5 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_B6 = CLBLL_L_X2Y142_SLICE_X0Y142_DQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A6 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B1 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO7;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_C1 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_C2 = CLBLL_L_X2Y142_SLICE_X0Y142_AQ;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_C3 = CLBLL_L_X2Y142_SLICE_X0Y142_DQ;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_C4 = CLBLL_L_X2Y142_SLICE_X0Y142_BQ;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_C5 = CLBLL_L_X2Y142_SLICE_X0Y142_CQ;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_C6 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B4 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO7;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B5 = CLBLL_L_X4Y145_SLICE_X4Y145_BQ;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_BX = CLBLL_L_X4Y133_SLICE_X5Y133_DO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C1 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO1;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C2 = BRAM_L_X6Y140_RAMB18_X0Y56_DO18;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C3 = CLBLM_R_X5Y130_SLICE_X6Y130_DQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C4 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_D1 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_D2 = CLBLL_L_X2Y142_SLICE_X0Y142_AQ;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_D3 = CLBLL_L_X2Y142_SLICE_X0Y142_DQ;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_D4 = CLBLL_L_X2Y142_SLICE_X0Y142_BQ;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_D5 = CLBLL_L_X2Y142_SLICE_X0Y142_CQ;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_D6 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D1 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D2 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D3 = CLBLM_R_X5Y130_SLICE_X6Y130_DQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D4 = CLBLM_R_X5Y133_SLICE_X6Y133_CO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D5 = CLBLM_R_X3Y147_SLICE_X3Y147_DQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D6 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_A1 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_A2 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_A3 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_A4 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_A5 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_A6 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_B1 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_B2 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_B3 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_B4 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_B5 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_B6 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_C1 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_C2 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_C3 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_C4 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_C5 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_C6 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_D1 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_D2 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_D3 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_D4 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_D5 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_D6 = 1'b1;
  assign RIOI3_X105Y83_OLOGIC_X1Y84_D1 = CLBLM_L_X10Y132_SLICE_X12Y132_BQ;
  assign RIOI3_X105Y83_OLOGIC_X1Y84_T1 = 1'b1;
  assign RIOI3_X105Y83_OLOGIC_X1Y83_D1 = CLBLM_L_X8Y131_SLICE_X10Y131_BQ;
  assign RIOI3_X105Y83_OLOGIC_X1Y83_T1 = 1'b1;
  assign RIOB33_X105Y127_IOB_X1Y128_O = CLBLM_L_X8Y134_SLICE_X10Y134_AQ;
  assign RIOB33_X105Y127_IOB_X1Y127_O = CLBLM_R_X5Y133_SLICE_X7Y133_AQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A1 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A2 = CLBLM_R_X5Y134_SLICE_X7Y134_A5Q;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A3 = BRAM_L_X6Y125_RAMB18_X0Y50_DO23;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A5 = BRAM_L_X6Y135_RAMB18_X0Y54_DO7;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A6 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B1 = BRAM_L_X6Y140_RAMB18_X0Y56_DO23;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B2 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B3 = CLBLL_L_X4Y132_SLICE_X5Y132_BQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B4 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B5 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B6 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C1 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO4;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C2 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C3 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C4 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C5 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C6 = CLBLM_R_X5Y131_SLICE_X7Y131_CQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D1 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D2 = CLBLM_R_X7Y132_SLICE_X8Y132_CQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D3 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D4 = CLBLM_R_X3Y147_SLICE_X2Y147_BQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D5 = CLBLM_R_X7Y134_SLICE_X8Y134_AO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D6 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A1 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_ADDRARDADDR0 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_ADDRARDADDR1 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_ADDRARDADDR2 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_ADDRARDADDR3 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_ADDRARDADDR4 = CLBLM_R_X5Y129_SLICE_X7Y129_DO6;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_ADDRARDADDR5 = CLBLM_R_X5Y129_SLICE_X7Y129_CO6;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_ADDRARDADDR6 = CLBLL_L_X4Y129_SLICE_X5Y129_DO6;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_ADDRARDADDR7 = CLBLM_R_X5Y129_SLICE_X6Y129_CO6;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_ADDRARDADDR8 = CLBLM_R_X5Y130_SLICE_X6Y130_DO6;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_ADDRARDADDR9 = CLBLL_L_X4Y130_SLICE_X4Y130_DO6;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_ADDRARDADDR10 = CLBLL_L_X4Y130_SLICE_X5Y130_CO6;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_ADDRARDADDR11 = CLBLM_R_X3Y134_SLICE_X3Y134_AO6;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_ADDRARDADDR12 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_ADDRARDADDR13 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_ADDRATIEHIGH0 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_ADDRATIEHIGH1 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_ADDRBTIEHIGH0 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_ADDRBTIEHIGH1 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_ADDRBWRADDR0 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_ADDRBWRADDR1 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_ADDRBWRADDR2 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_ADDRBWRADDR3 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_ADDRBWRADDR4 = CLBLM_R_X5Y130_SLICE_X6Y130_CO6;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_ADDRBWRADDR5 = CLBLL_L_X4Y130_SLICE_X5Y130_BO6;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_ADDRBWRADDR6 = CLBLL_L_X4Y130_SLICE_X4Y130_CO6;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_ADDRBWRADDR7 = CLBLM_R_X5Y132_SLICE_X6Y132_DO6;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_ADDRBWRADDR8 = CLBLM_R_X5Y131_SLICE_X6Y131_DO6;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_ADDRBWRADDR9 = CLBLM_R_X5Y132_SLICE_X6Y132_CO6;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_ADDRBWRADDR10 = CLBLL_L_X4Y132_SLICE_X4Y132_DO6;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_ADDRBWRADDR11 = CLBLL_L_X4Y133_SLICE_X5Y133_CO6;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_ADDRBWRADDR12 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_ADDRBWRADDR13 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_DIADI5 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C4 = CLBLL_L_X4Y132_SLICE_X5Y132_A5Q;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_RDCLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_WRCLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_DIADI0 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D2 = CLBLL_L_X2Y155_SLICE_X0Y155_CQ;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_DIADI1 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_DIADI2 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_DIADI3 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_DIADI4 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_DIADI5 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_DIADI6 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_DIADI7 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_DIADI8 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_DIADI9 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_DIADI10 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_DIADI11 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_DIADI12 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_DIADI13 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_DIADI14 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_DIADI15 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_DIBDI0 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_DIBDI1 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_DIBDI2 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_DIBDI3 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_DIBDI4 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_DIBDI5 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_DIBDI6 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_DIBDI7 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_DIBDI8 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_DIBDI9 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_DIBDI10 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_DIBDI11 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_DIBDI12 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_DIBDI13 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_DIBDI14 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_DIBDI15 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_DIPADIP0 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_DIPADIP1 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_DIPBDIP0 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_DIPBDIP1 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_DIADI13 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_DIADI15 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_DIBDI0 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y8_D = LIOB33_X0Y7_IOB_X0Y8_I;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_RDEN = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_WREN = 1'b1;
  assign LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y7_D = LIOB33_X0Y7_IOB_X0Y7_I;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_DIBDI6 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_REGCE = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_REGCEB = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_RDRCLK = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_REGCLKB = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_RST = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_RSTRAMB = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_RSTREG = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_RSTREGB = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_WEA0 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_WEA1 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_WEA2 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_WEA3 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_WEBWE0 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_WEBWE1 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_WEBWE2 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_WEBWE3 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_WEBWE4 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_WEBWE5 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_WEBWE6 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y52_WEBWE7 = 1'b0;
  assign RIOB33_X105Y129_IOB_X1Y130_O = CLBLM_L_X8Y132_SLICE_X11Y132_BQ;
  assign RIOB33_X105Y129_IOB_X1Y129_O = CLBLM_R_X7Y133_SLICE_X9Y133_AQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D1 = BRAM_L_X6Y140_RAMB18_X0Y56_DO19;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D2 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO3;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D3 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO3;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D4 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO2;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D5 = CLBLM_R_X5Y129_SLICE_X6Y129_A5Q;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D6 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO2;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A1 = BRAM_L_X6Y140_RAMB18_X0Y56_DO5;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A2 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO5;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A3 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO4;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A4 = CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A5 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO4;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A6 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO5;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B1 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B2 = BRAM_L_X6Y140_RAMB18_X0Y56_DO22;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B3 = CLBLM_R_X5Y132_SLICE_X7Y132_A5Q;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B4 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO5;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B5 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO5;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B6 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C1 = CLBLM_R_X3Y134_SLICE_X2Y134_AQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C2 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO7;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C3 = BRAM_R_X17Y135_RAMB18_X1Y54_DO23;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C4 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO7;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C5 = BRAM_L_X6Y135_RAMB18_X0Y54_DO22;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C6 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D1 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO5;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D2 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D3 = BRAM_L_X6Y140_RAMB18_X0Y56_DO22;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D4 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D5 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO5;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D6 = CLBLM_R_X5Y130_SLICE_X6Y130_B5Q;
  assign RIOB33_X105Y131_IOB_X1Y132_O = CLBLL_L_X54Y133_SLICE_X82Y133_AQ;
  assign RIOB33_X105Y131_IOB_X1Y131_O = CLBLM_R_X5Y134_SLICE_X7Y134_BQ;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A1 = CLBLM_R_X3Y142_SLICE_X2Y142_DQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A2 = CLBLM_R_X5Y129_SLICE_X7Y129_B5Q;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A3 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO7;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A4 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A5 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO7;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A6 = CLBLM_R_X5Y136_SLICE_X7Y136_CO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B1 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B2 = CLBLL_L_X4Y131_SLICE_X5Y131_CQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B3 = BRAM_L_X6Y140_RAMB18_X0Y56_DO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B4 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO5;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B5 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO5;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B6 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO6;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1 = CLBLM_L_X8Y135_SLICE_X10Y135_AQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C1 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO1;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C2 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO0;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C3 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO0;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C4 = BRAM_L_X6Y140_RAMB18_X0Y56_DO17;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C5 = CLBLM_R_X5Y129_SLICE_X7Y129_B5Q;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C6 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO1;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D1 = CLBLM_R_X3Y155_SLICE_X3Y155_AQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D2 = CLBLL_L_X4Y131_SLICE_X5Y131_CQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D3 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D4 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D5 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D6 = CLBLM_R_X5Y136_SLICE_X7Y136_BO6;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A1 = BRAM_L_X6Y140_RAMB18_X0Y56_DO3;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A2 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO2;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A3 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO2;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A4 = CLBLM_R_X5Y132_SLICE_X6Y132_BQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A5 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO3;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A6 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO3;
  assign RIOI3_X105Y85_OLOGIC_X1Y86_D1 = CLBLM_L_X8Y132_SLICE_X11Y132_CQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B1 = CLBLL_L_X4Y155_SLICE_X4Y155_BQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B2 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B3 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO7;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B4 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO7;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B5 = CLBLM_R_X5Y136_SLICE_X6Y136_AO6;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B6 = CLBLM_R_X5Y132_SLICE_X6Y132_BQ;
  assign RIOI3_X105Y85_OLOGIC_X1Y86_T1 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C1 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C2 = BRAM_L_X6Y140_RAMB18_X0Y56_DO18;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C3 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO2;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C4 = CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C5 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C6 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO2;
  assign RIOI3_X105Y85_OLOGIC_X1Y85_D1 = CLBLM_L_X10Y132_SLICE_X12Y132_CQ;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1 = 1'b1;
  assign RIOI3_X105Y85_OLOGIC_X1Y85_T1 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D1 = CLBLM_R_X5Y137_SLICE_X7Y137_BO6;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D2 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO7;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D3 = CLBLM_R_X3Y153_SLICE_X2Y153_BQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D4 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D5 = CLBLM_R_X5Y129_SLICE_X6Y129_BQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D6 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO7;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A2 = BRAM_L_X6Y130_RAMB18_X0Y52_DO3;
  assign LIOI3_X0Y165_ILOGIC_X0Y166_D = LIOB33_X0Y165_IOB_X0Y166_I;
  assign RIOB33_X105Y133_IOB_X1Y134_O = CLBLM_R_X5Y133_SLICE_X7Y133_BQ;
  assign RIOB33_X105Y133_IOB_X1Y133_O = CLBLM_R_X7Y133_SLICE_X9Y133_BQ;
  assign LIOI3_X0Y165_ILOGIC_X0Y165_D = LIOB33_X0Y165_IOB_X0Y165_I;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A3 = CLBLM_R_X5Y133_SLICE_X6Y133_AQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B2 = CLBLM_R_X5Y133_SLICE_X7Y133_DO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B3 = CLBLM_R_X7Y130_SLICE_X8Y130_B5Q;
  assign LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y20_D = LIOB33_X0Y19_IOB_X0Y20_I;
  assign LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y19_D = LIOB33_X0Y19_IOB_X0Y19_I;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B6 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_A1 = 1'b1;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_A2 = 1'b1;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_A3 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO5;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_A4 = CLBLM_R_X5Y127_SLICE_X7Y127_BQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_A5 = 1'b1;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_A6 = 1'b1;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_B1 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO1;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_B2 = BRAM_L_X6Y140_RAMB18_X0Y56_DO1;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_B3 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO0;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_B4 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO1;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_B5 = CLBLM_R_X5Y129_SLICE_X6Y129_BQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_B6 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO0;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C5 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO2;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_C1 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO4;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C6 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO2;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_C2 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO3;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_C3 = CLBLM_R_X5Y126_SLICE_X7Y126_BQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_C4 = BRAM_L_X6Y140_RAMB18_X0Y56_DO4;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_C5 = BRAM_L_X6Y140_RAMB18_X0Y56_DO3;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_C6 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO4;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_D1 = BRAM_L_X6Y140_RAMB18_X0Y56_DO7;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_D2 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_D3 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO7;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_D4 = CLBLM_R_X5Y137_SLICE_X7Y137_CO6;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_D5 = CLBLM_R_X5Y126_SLICE_X7Y126_BQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_D6 = CLBLM_R_X3Y153_SLICE_X3Y153_BQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_A1 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO4;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_A2 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO5;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_A3 = CLBLM_R_X3Y130_SLICE_X3Y130_BQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_A4 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO4;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_A5 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO5;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_A6 = BRAM_L_X6Y140_RAMB18_X0Y56_DO5;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_B1 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_B2 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO7;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_B3 = CLBLL_L_X4Y134_SLICE_X4Y134_AQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_B4 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_B5 = BRAM_L_X6Y140_RAMB18_X0Y56_DO23;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_B6 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO7;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_C1 = CLBLM_R_X3Y130_SLICE_X3Y130_BQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_C2 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_C3 = 1'b1;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_C4 = CLBLM_R_X5Y137_SLICE_X6Y137_AO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_C5 = 1'b1;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_C6 = CLBLL_L_X2Y155_SLICE_X1Y155_AQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_D1 = CLBLL_L_X4Y134_SLICE_X4Y134_AQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_D2 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_D3 = 1'b1;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_D4 = CLBLM_R_X3Y145_SLICE_X3Y145_AQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_D5 = 1'b1;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_D6 = CLBLM_R_X5Y137_SLICE_X6Y137_BO6;
  assign RIOB33_X105Y135_IOB_X1Y136_O = CLBLM_R_X5Y135_SLICE_X7Y135_AQ;
  assign RIOB33_X105Y135_IOB_X1Y135_O = CLBLM_R_X7Y137_SLICE_X9Y137_AQ;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A1 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A2 = CLBLL_L_X4Y131_SLICE_X5Y131_CQ;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A3 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A4 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A5 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A6 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B1 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO3;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B2 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO3;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B3 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO2;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B4 = BRAM_L_X6Y140_RAMB18_X0Y56_DO18;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B5 = CLBLM_R_X5Y129_SLICE_X7Y129_AQ;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B6 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO3;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C1 = BRAM_L_X6Y140_RAMB18_X0Y56_DO23;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C2 = CLBLM_R_X5Y126_SLICE_X7Y126_B5Q;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C3 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO7;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C4 = CLBLM_R_X3Y142_SLICE_X2Y142_CQ;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C5 = CLBLM_R_X5Y138_SLICE_X7Y138_DO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C6 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D1 = BRAM_L_X6Y140_RAMB18_X0Y56_DO18;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D2 = CLBLM_R_X5Y126_SLICE_X7Y126_B5Q;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D3 = BRAM_L_X6Y140_RAMB18_X0Y56_DO19;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D4 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO3;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D5 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO3;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D6 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO2;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A1 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO4;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A2 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A3 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A4 = CLBLL_L_X4Y131_SLICE_X5Y131_BQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A5 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A6 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B1 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B2 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B3 = CLBLM_R_X3Y130_SLICE_X3Y130_BQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B4 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO5;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B5 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B6 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C1 = CLBLL_L_X4Y127_SLICE_X5Y127_AQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C2 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C3 = BRAM_L_X6Y140_RAMB18_X0Y56_DO5;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C4 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO5;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C5 = BRAM_L_X6Y140_RAMB18_X0Y56_DO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C6 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D1 = CLBLL_L_X4Y127_SLICE_X5Y127_AQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D2 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D3 = CLBLM_R_X3Y153_SLICE_X3Y153_CQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D4 = CLBLM_R_X5Y138_SLICE_X6Y138_CO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D5 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D6 = 1'b1;
  assign RIOI3_X105Y111_OLOGIC_X1Y112_D1 = CLBLM_R_X7Y131_SLICE_X9Y131_BQ;
  assign RIOB33_X105Y137_IOB_X1Y138_O = CLBLM_R_X7Y137_SLICE_X8Y137_BQ;
  assign RIOB33_X105Y137_IOB_X1Y137_O = CLBLM_R_X5Y137_SLICE_X7Y137_AQ;
  assign RIOI3_X105Y89_OLOGIC_X1Y90_D1 = CLBLM_L_X10Y130_SLICE_X12Y130_BQ;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_ADDRARDADDR0 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_ADDRARDADDR1 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_ADDRARDADDR2 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_ADDRARDADDR3 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_ADDRARDADDR4 = CLBLL_L_X4Y137_SLICE_X4Y137_CO6;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_ADDRARDADDR5 = CLBLL_L_X4Y138_SLICE_X4Y138_BO6;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_ADDRARDADDR6 = CLBLM_R_X3Y137_SLICE_X2Y137_CO6;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_ADDRARDADDR7 = CLBLM_R_X5Y136_SLICE_X6Y136_BO6;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_ADDRARDADDR8 = CLBLL_L_X4Y135_SLICE_X4Y135_CO6;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_ADDRARDADDR9 = CLBLM_R_X5Y134_SLICE_X6Y134_DO6;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_ADDRARDADDR10 = CLBLL_L_X4Y135_SLICE_X4Y135_DO6;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_ADDRARDADDR11 = CLBLM_R_X3Y137_SLICE_X3Y137_DO6;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_ADDRARDADDR12 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_ADDRARDADDR13 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_ADDRATIEHIGH0 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_ADDRATIEHIGH1 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_ADDRBTIEHIGH0 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_ADDRBTIEHIGH1 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_ADDRBWRADDR0 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_ADDRBWRADDR1 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_ADDRBWRADDR2 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_ADDRBWRADDR3 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_ADDRBWRADDR4 = CLBLL_L_X4Y134_SLICE_X5Y134_CO6;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_ADDRBWRADDR5 = CLBLM_R_X5Y133_SLICE_X6Y133_BO6;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_ADDRBWRADDR6 = CLBLM_R_X5Y133_SLICE_X6Y133_DO6;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_ADDRBWRADDR7 = CLBLM_R_X7Y133_SLICE_X8Y133_AO6;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_ADDRBWRADDR8 = CLBLM_R_X7Y135_SLICE_X8Y135_AO6;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_ADDRBWRADDR9 = CLBLM_R_X5Y134_SLICE_X7Y134_DO6;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_ADDRBWRADDR10 = CLBLM_R_X3Y135_SLICE_X3Y135_AO6;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_ADDRBWRADDR11 = CLBLL_L_X4Y134_SLICE_X5Y134_DO6;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_ADDRBWRADDR12 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_ADDRBWRADDR13 = 1'b0;
  assign RIOI3_X105Y89_OLOGIC_X1Y89_T1 = 1'b1;
  assign RIOI3_X105Y111_OLOGIC_X1Y112_T1 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_CLKARDCLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_CLKBWRCLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_DIADI0 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_DIADI1 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_DIADI2 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_DIADI3 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_DIADI4 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_DIADI5 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_DIADI6 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_DIADI7 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_DIADI8 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_DIADI9 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_DIADI10 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_DIADI11 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_DIADI12 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_DIADI13 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_DIADI14 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_DIADI15 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_DIBDI0 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_DIBDI1 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_DIBDI2 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_DIBDI3 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_DIBDI4 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_DIBDI5 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_DIBDI6 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_DIBDI7 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_DIBDI8 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_DIBDI9 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_DIBDI10 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_DIBDI11 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_DIBDI12 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_DIBDI13 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_DIBDI14 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_DIBDI15 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_DIPADIP0 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_DIPADIP1 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_DIPBDIP0 = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_DIPBDIP1 = 1'b1;
  assign RIOI3_X105Y111_OLOGIC_X1Y111_D1 = CLBLM_R_X7Y130_SLICE_X9Y130_AQ;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_ENARDEN = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_ENBWREN = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_REGCEAREGCE = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_REGCEB = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_REGCLKARDRCLK = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_REGCLKB = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_RSTRAMARSTRAM = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_RSTRAMB = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_RSTREGARSTREG = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_RSTREGB = 1'b1;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_WEA0 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_WEA1 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_WEA2 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_WEA3 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_WEBWE0 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_WEBWE1 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_WEBWE2 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_WEBWE3 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_WEBWE4 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_WEBWE5 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_WEBWE6 = 1'b0;
  assign BRAM_L_X6Y130_RAMB18_X0Y53_WEBWE7 = 1'b0;
  assign RIOI3_X105Y111_OLOGIC_X1Y111_T1 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A1 = CLBLM_R_X3Y149_SLICE_X2Y149_CQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A2 = CLBLM_R_X5Y138_SLICE_X7Y138_BO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A3 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO7;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A4 = BRAM_L_X6Y140_RAMB18_X0Y56_DO23;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A5 = CLBLM_R_X5Y129_SLICE_X7Y129_AQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A6 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign LIOI3_X0Y167_ILOGIC_X0Y168_D = LIOB33_X0Y167_IOB_X0Y168_I;
  assign LIOI3_X0Y167_ILOGIC_X0Y167_D = LIOB33_X0Y167_IOB_X0Y167_I;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B1 = BRAM_L_X6Y140_RAMB18_X0Y56_DO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B2 = CLBLM_R_X3Y132_SLICE_X3Y132_CQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B3 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO7;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B4 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO7;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B5 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO7;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B6 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C1 = BRAM_L_X6Y140_RAMB18_X0Y56_DO21;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C2 = CLBLM_R_X5Y127_SLICE_X7Y127_CQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C3 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C4 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO5;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C5 = BRAM_L_X6Y140_RAMB18_X0Y56_DO22;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C6 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D1 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D2 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D3 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D4 = CLBLM_R_X5Y139_SLICE_X7Y139_CO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D5 = CLBLM_R_X3Y145_SLICE_X2Y145_CQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D6 = CLBLM_R_X5Y127_SLICE_X7Y127_CQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A1 = CLBLL_L_X4Y132_SLICE_X5Y132_BQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A2 = BRAM_L_X6Y140_RAMB18_X0Y56_DO22;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A3 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO7;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A4 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO7;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A5 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO7;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A6 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B1 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B2 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO2;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B3 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO2;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B4 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO1;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B5 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO2;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B6 = BRAM_L_X6Y140_RAMB18_X0Y56_DO17;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C1 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO1;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C2 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO1;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C3 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO0;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C4 = CLBLM_R_X5Y132_SLICE_X6Y132_B5Q;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C5 = BRAM_L_X6Y140_RAMB18_X0Y56_DO16;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C6 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO1;
  assign LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y31_D = LIOB33_X0Y31_IOB_X0Y31_I;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D1 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO7;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D2 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D3 = BRAM_L_X6Y140_RAMB18_X0Y56_DO22;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D4 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO7;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D5 = CLBLM_R_X5Y127_SLICE_X7Y127_DQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D6 = BRAM_L_X6Y140_RAMB18_X0Y56_DO23;
  assign RIOB33_X105Y139_IOB_X1Y140_O = CLBLM_R_X7Y138_SLICE_X9Y138_AQ;
  assign RIOB33_X105Y139_IOB_X1Y139_O = CLBLL_L_X54Y138_SLICE_X82Y138_AQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A1 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A2 = CLBLM_R_X5Y139_SLICE_X7Y139_BO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A3 = CLBLM_R_X3Y132_SLICE_X3Y132_CQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A4 = CLBLL_L_X2Y155_SLICE_X0Y155_DQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A5 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A6 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B1 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B2 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B3 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B4 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B5 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B6 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C1 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C2 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C3 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C4 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C5 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C6 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D1 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D2 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D3 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D4 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D5 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D6 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A1 = CLBLM_R_X5Y132_SLICE_X6Y132_B5Q;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A2 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO7;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A3 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A4 = CLBLM_R_X5Y139_SLICE_X6Y139_CO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A5 = BRAM_L_X6Y140_RAMB18_X0Y56_DO23;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A6 = CLBLM_R_X3Y149_SLICE_X2Y149_AQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B1 = CLBLM_R_X5Y139_SLICE_X6Y139_BO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B2 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B3 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B4 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B5 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B6 = CLBLM_R_X3Y149_SLICE_X2Y149_BQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C1 = CLBLM_R_X5Y139_SLICE_X6Y139_AO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C2 = CLBLL_L_X4Y132_SLICE_X5Y132_BQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C3 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C4 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C5 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C6 = CLBLM_R_X3Y151_SLICE_X2Y151_AQ;
  assign RIOB33_X105Y141_IOB_X1Y142_O = CLBLM_R_X7Y138_SLICE_X9Y138_CQ;
  assign RIOB33_X105Y141_IOB_X1Y141_O = CLBLM_R_X7Y138_SLICE_X9Y138_BQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D1 = CLBLM_R_X5Y127_SLICE_X7Y127_DQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D2 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D3 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D4 = CLBLM_R_X5Y139_SLICE_X6Y139_DO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D5 = CLBLM_R_X3Y145_SLICE_X2Y145_DQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D6 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_A1 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_A2 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_A3 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_A4 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_A5 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_A6 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_B1 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_B2 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_B3 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_B4 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_B5 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_B6 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_C1 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_C2 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_C3 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_C4 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_C5 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_C6 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D4 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_D1 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_D2 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_D3 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_D4 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_D5 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_D6 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_A1 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_A2 = BRAM_R_X17Y135_RAMB18_X1Y54_DO3;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_A3 = CLBLM_R_X5Y130_SLICE_X6Y130_AQ;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_A4 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_A5 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_A6 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D5 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_B1 = CLBLM_R_X3Y132_SLICE_X3Y132_AQ;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_B2 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_B3 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_B4 = BRAM_R_X17Y135_RAMB18_X1Y54_DO4;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_B5 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_B6 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_C1 = CLBLM_L_X10Y135_SLICE_X13Y135_AO6;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_C2 = BRAM_R_X17Y135_RAMB18_X1Y54_DO7;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_C3 = CLBLM_R_X3Y132_SLICE_X3Y132_AQ;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_C4 = CLBLM_R_X25Y157_SLICE_X36Y157_BQ;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_C5 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_C6 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO7;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D6 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_D1 = CLBLM_R_X5Y130_SLICE_X6Y130_AQ;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_D2 = BRAM_R_X17Y135_RAMB18_X1Y54_DO7;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_D3 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_D4 = CLBLM_L_X10Y135_SLICE_X12Y135_CO6;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_D5 = CLBLM_L_X16Y157_SLICE_X22Y157_AQ;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_D6 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO7;
  assign RIOI3_X105Y91_OLOGIC_X1Y92_D1 = CLBLM_R_X11Y131_SLICE_X14Y131_AQ;
  assign RIOI3_X105Y91_OLOGIC_X1Y92_T1 = 1'b1;
  assign RIOI3_X105Y91_OLOGIC_X1Y91_D1 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign RIOI3_X105Y91_OLOGIC_X1Y91_T1 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A2 = CLBLM_R_X7Y132_SLICE_X8Y132_A5Q;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A3 = BRAM_L_X6Y135_RAMB18_X0Y54_DO4;
  assign RIOB33_X105Y143_IOB_X1Y144_O = CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  assign RIOB33_X105Y143_IOB_X1Y143_O = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A1 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO3;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_A1 = 1'b1;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_A2 = 1'b1;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_A3 = 1'b1;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_A4 = 1'b1;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_A5 = 1'b1;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_A6 = 1'b1;
  assign RIOB33_X105Y145_IOB_X1Y146_O = CLBLM_R_X5Y138_SLICE_X7Y138_AQ;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_B1 = 1'b1;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_B2 = 1'b1;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_B3 = 1'b1;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_B4 = 1'b1;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_B5 = 1'b1;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_B6 = 1'b1;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_C1 = 1'b1;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_C2 = 1'b1;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_C3 = 1'b1;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_C4 = 1'b1;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_C5 = 1'b1;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_C6 = 1'b1;
  assign LIOI3_X0Y171_ILOGIC_X0Y172_D = LIOB33_X0Y171_IOB_X0Y172_I;
  assign LIOI3_X0Y171_ILOGIC_X0Y171_D = LIOB33_X0Y171_IOB_X0Y171_I;
  assign RIOB33_X105Y145_IOB_X1Y145_O = CLBLM_R_X5Y138_SLICE_X6Y138_BQ;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_D1 = 1'b1;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_D2 = 1'b1;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_D3 = 1'b1;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_D4 = 1'b1;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_D5 = 1'b1;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_D6 = 1'b1;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_A1 = CLBLM_R_X3Y131_SLICE_X3Y131_B5Q;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_A2 = 1'b1;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_A3 = 1'b1;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_A4 = BRAM_R_X17Y135_RAMB18_X1Y54_DO2;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_A5 = 1'b1;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_A6 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_ADDRARDADDR0 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_ADDRARDADDR1 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_ADDRARDADDR2 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_ADDRARDADDR3 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_ADDRARDADDR4 = CLBLL_L_X4Y137_SLICE_X5Y137_DO6;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_ADDRARDADDR5 = CLBLM_R_X5Y136_SLICE_X6Y136_DO6;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_ADDRARDADDR6 = CLBLL_L_X4Y136_SLICE_X5Y136_DO6;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_ADDRARDADDR7 = CLBLL_L_X4Y136_SLICE_X4Y136_CO6;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_ADDRARDADDR8 = CLBLL_L_X4Y137_SLICE_X5Y137_CO6;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_ADDRARDADDR9 = CLBLM_R_X5Y137_SLICE_X6Y137_CO6;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_ADDRARDADDR10 = CLBLM_R_X5Y136_SLICE_X7Y136_DO6;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_ADDRARDADDR11 = CLBLM_R_X3Y137_SLICE_X2Y137_DO6;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_ADDRARDADDR12 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_ADDRARDADDR13 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_ADDRATIEHIGH0 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_ADDRATIEHIGH1 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_ADDRBTIEHIGH0 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_ADDRBTIEHIGH1 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_ADDRBWRADDR0 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_ADDRBWRADDR1 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_ADDRBWRADDR2 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_ADDRBWRADDR3 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_ADDRBWRADDR4 = CLBLL_L_X4Y135_SLICE_X5Y135_DO6;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_ADDRBWRADDR5 = CLBLM_R_X5Y136_SLICE_X7Y136_AO6;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_ADDRBWRADDR6 = CLBLL_L_X4Y136_SLICE_X5Y136_CO6;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_ADDRBWRADDR7 = CLBLM_R_X5Y135_SLICE_X7Y135_CO6;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_ADDRBWRADDR8 = CLBLM_R_X7Y138_SLICE_X8Y138_AO6;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_ADDRBWRADDR9 = CLBLM_R_X7Y137_SLICE_X8Y137_DO6;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_ADDRBWRADDR10 = CLBLM_R_X3Y135_SLICE_X3Y135_DO6;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_ADDRBWRADDR11 = CLBLM_R_X5Y137_SLICE_X6Y137_DO6;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_ADDRBWRADDR12 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_ADDRBWRADDR13 = 1'b0;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_D1 = CLBLM_L_X16Y155_SLICE_X22Y155_AQ;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_RDCLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_WRCLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_DIADI0 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_DIADI1 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_DIADI2 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_DIADI3 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_DIADI4 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_DIADI5 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_DIADI6 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_DIADI7 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_DIADI8 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_DIADI9 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_DIADI10 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_DIADI11 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_DIADI12 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_DIADI13 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_DIADI14 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_DIADI15 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_DIBDI0 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_DIBDI1 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_DIBDI2 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_DIBDI3 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_DIBDI4 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_DIBDI5 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_DIBDI6 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_DIBDI7 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_DIBDI8 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_DIBDI9 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_DIBDI10 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_DIBDI11 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_DIBDI12 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_DIBDI13 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_DIBDI14 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_DIBDI15 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_DIPADIP0 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_DIPADIP1 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_DIPBDIP0 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_DIPBDIP1 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A3 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A4 = CLBLL_L_X4Y134_SLICE_X4Y134_AQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A5 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO7;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A6 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_RDEN = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_WREN = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B1 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B2 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B3 = CLBLM_R_X5Y127_SLICE_X7Y127_DQ;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_REGCE = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_REGCEB = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_RDRCLK = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_REGCLKB = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_RST = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_RSTRAMB = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_RSTREG = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_RSTREGB = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_WEA0 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_WEA1 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_WEA2 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_WEA3 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_WEBWE0 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_WEBWE1 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_WEBWE2 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_WEBWE3 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_WEBWE4 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_WEBWE5 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_WEBWE6 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y54_WEBWE7 = 1'b0;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B6 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B3 = CLBLM_L_X16Y153_SLICE_X22Y153_AQ;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_A1 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_A2 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_A3 = BRAM_R_X17Y135_RAMB18_X1Y54_DO6;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_A4 = CLBLM_R_X3Y132_SLICE_X2Y132_AQ;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_A5 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_A6 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_B1 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_B2 = BRAM_R_X17Y135_RAMB18_X1Y54_DO7;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_B3 = CLBLM_R_X3Y132_SLICE_X2Y132_BQ;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_B4 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_B5 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_B6 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_C1 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_C2 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_C3 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_C4 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_C5 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_C6 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_D1 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_D2 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_D3 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_D4 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_D5 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_D6 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign RIOB33_X105Y147_IOB_X1Y148_O = CLBLM_R_X7Y137_SLICE_X9Y137_BQ;
  assign RIOB33_X105Y147_IOB_X1Y147_O = CLBLL_L_X54Y141_SLICE_X82Y141_AQ;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_A1 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_A2 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_A3 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_A4 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_A5 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_C2 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_C3 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_C4 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_C6 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_D1 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_D2 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_D3 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_D4 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_D5 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_D6 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_A1 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_A2 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_A3 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_A4 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_A5 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_A6 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_AX = LIOB33_X0Y205_IOB_X0Y205_I;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_B1 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_B2 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_B3 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_B4 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_B5 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_B6 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_B1 = 1'b1;
  assign RIOI3_X105Y95_OLOGIC_X1Y96_D1 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_C1 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_C2 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_C3 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_C4 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_C5 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_C6 = 1'b1;
  assign RIOI3_X105Y95_OLOGIC_X1Y96_T1 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_D1 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_D2 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_D3 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_D4 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_D5 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_D6 = 1'b1;
  assign RIOI3_X105Y95_OLOGIC_X1Y95_D1 = CLBLM_R_X11Y131_SLICE_X14Y131_BQ;
  assign RIOI3_X105Y95_OLOGIC_X1Y95_T1 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_C4 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_C5 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_C6 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign LIOI3_X0Y173_ILOGIC_X0Y174_D = LIOB33_X0Y173_IOB_X0Y174_I;
  assign LIOI3_X0Y173_ILOGIC_X0Y173_D = LIOB33_X0Y173_IOB_X0Y173_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_D = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_D = LIOB33_X0Y51_IOB_X0Y51_I;
  assign RIOB33_X105Y151_IOB_X1Y152_O = CLBLM_R_X7Y129_SLICE_X9Y129_BQ;
  assign RIOB33_X105Y151_IOB_X1Y151_O = CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D = LIOB33_X0Y57_IOB_X0Y57_I;
  assign RIOB33_X105Y153_IOB_X1Y154_O = CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  assign RIOB33_X105Y153_IOB_X1Y153_O = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign RIOB33_X105Y91_IOB_X1Y92_O = CLBLM_R_X11Y131_SLICE_X14Y131_AQ;
  assign RIOI3_X105Y97_OLOGIC_X1Y98_D1 = CLBLM_R_X7Y125_SLICE_X8Y125_CQ;
  assign RIOI3_X105Y97_OLOGIC_X1Y98_T1 = 1'b1;
  assign RIOB33_X105Y155_IOB_X1Y156_O = CLBLM_R_X7Y129_SLICE_X8Y129_BQ;
  assign RIOB33_X105Y155_IOB_X1Y155_O = CLBLM_R_X7Y136_SLICE_X8Y136_AQ;
  assign RIOI3_X105Y97_OLOGIC_X1Y97_D1 = CLBLM_R_X7Y125_SLICE_X8Y125_BQ;
  assign RIOI3_X105Y97_OLOGIC_X1Y97_T1 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B5 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B6 = CLBLM_R_X3Y132_SLICE_X2Y132_DQ;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_ADDRARDADDR0 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_ADDRARDADDR1 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_ADDRARDADDR2 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_ADDRARDADDR3 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_ADDRARDADDR4 = CLBLM_L_X10Y136_SLICE_X12Y136_DO6;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_ADDRARDADDR5 = CLBLM_L_X8Y137_SLICE_X10Y137_DO6;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_ADDRARDADDR6 = CLBLM_R_X7Y136_SLICE_X9Y136_DO6;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_ADDRARDADDR7 = CLBLM_L_X8Y136_SLICE_X10Y136_CO6;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_ADDRARDADDR8 = CLBLM_L_X8Y136_SLICE_X11Y136_BO6;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_ADDRARDADDR9 = CLBLM_L_X10Y137_SLICE_X13Y137_BO6;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_ADDRARDADDR10 = CLBLM_L_X10Y137_SLICE_X12Y137_CO6;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_ADDRARDADDR11 = CLBLM_L_X8Y137_SLICE_X11Y137_CO6;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_ADDRARDADDR12 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_ADDRARDADDR13 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_ADDRATIEHIGH0 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_ADDRATIEHIGH1 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_ADDRBTIEHIGH0 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_ADDRBTIEHIGH1 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_ADDRBWRADDR0 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_ADDRBWRADDR1 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_ADDRBWRADDR2 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_ADDRBWRADDR3 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_ADDRBWRADDR4 = CLBLM_R_X7Y131_SLICE_X8Y131_AO6;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_ADDRBWRADDR5 = CLBLM_R_X7Y132_SLICE_X8Y132_BO6;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_ADDRBWRADDR6 = CLBLM_R_X7Y135_SLICE_X8Y135_DO6;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_A1 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_A2 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_ADDRBWRADDR7 = CLBLM_R_X7Y133_SLICE_X8Y133_CO6;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_ADDRBWRADDR8 = CLBLM_R_X7Y135_SLICE_X8Y135_BO6;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_A5 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_A3 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_A4 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_ADDRBWRADDR9 = CLBLM_R_X7Y135_SLICE_X8Y135_CO6;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_A6 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_ADDRBWRADDR10 = CLBLM_R_X3Y135_SLICE_X3Y135_BO6;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_ADDRBWRADDR11 = CLBLM_R_X3Y135_SLICE_X3Y135_CO6;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_B2 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_B3 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_B4 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_B5 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_B6 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_AX = LIOB33_SING_X0Y199_IOB_X0Y199_I;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_B1 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_CLKARDCLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_CLKBWRCLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_C1 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_C2 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_C3 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_DIADI3 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_BX = LIOB33_SING_X0Y200_IOB_X0Y200_I;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_C6 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_DIADI7 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_C4 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_C5 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_DIADI11 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_DIADI12 = 1'b0;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_CX = LIOB33_X0Y203_IOB_X0Y203_I;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_DIADI14 = 1'b0;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_D1 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_D2 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_D3 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_D4 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_D5 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_D6 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_DIBDI5 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_DIBDI6 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_DX = LIOB33_X0Y213_IOB_X0Y213_I;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_DIBDI8 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_DIBDI9 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_DIBDI10 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_DIBDI11 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_DIBDI12 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_DIBDI13 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_DIBDI14 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_DIBDI15 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_DIPADIP0 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_DIPADIP1 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_DIPBDIP0 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_DIPBDIP1 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B1 = BRAM_L_X6Y135_RAMB18_X0Y54_DO21;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B2 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B3 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO5;
  assign LIOI3_X0Y175_ILOGIC_X0Y176_D = LIOB33_X0Y175_IOB_X0Y176_I;
  assign LIOI3_X0Y175_ILOGIC_X0Y175_D = LIOB33_X0Y175_IOB_X0Y175_I;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B4 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B5 = BRAM_R_X17Y135_RAMB18_X1Y54_DO22;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_A1 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_A2 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_A3 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_A4 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_A5 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_A6 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B6 = CLBLL_L_X4Y131_SLICE_X5Y131_B5Q;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_AX = LIOB33_X0Y195_IOB_X0Y195_I;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_B1 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_B2 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_B3 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_B4 = 1'b1;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_D = LIOB33_X0Y53_IOB_X0Y54_I;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_ENARDEN = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_ENBWREN = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_B5 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_B6 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_BX = LIOB33_X0Y197_IOB_X0Y197_I;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_C1 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_C2 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_C3 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_C4 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_C5 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_C6 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_D = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A6 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO7;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_REGCEAREGCE = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_REGCEB = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_REGCLKARDRCLK = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_REGCLKB = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_D1 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_D2 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_D3 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_D4 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_D5 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_D6 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_RSTRAMARSTRAM = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_RSTRAMB = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_RSTREGARSTREG = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_RSTREGB = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_WEA0 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_WEA1 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_WEA2 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_WEA3 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_WEBWE0 = 1'b0;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_D = LIOB33_X0Y69_IOB_X0Y69_I;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_WEBWE1 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_WEBWE2 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_WEBWE3 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_WEBWE4 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_WEBWE5 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_WEBWE6 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_WEBWE7 = 1'b0;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C5 = CLBLM_R_X5Y135_SLICE_X7Y135_DO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C6 = CLBLM_R_X3Y142_SLICE_X2Y142_AQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B3 = BRAM_L_X6Y140_RAMB18_X0Y56_DO19;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOB33_X105Y157_IOB_X1Y158_O = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign RIOB33_X105Y157_IOB_X1Y157_O = CLBLM_L_X8Y130_SLICE_X10Y130_BQ;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_A6 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_AX = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_B1 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_B2 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_B3 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_B4 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_B5 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_B6 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_C1 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_C5 = 1'b1;
  assign RIOB33_X105Y159_IOB_X1Y160_O = CLBLM_R_X7Y137_SLICE_X8Y137_AQ;
  assign RIOB33_X105Y159_IOB_X1Y159_O = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign RIOI3_X105Y89_OLOGIC_X1Y90_T1 = 1'b1;
  assign RIOI3_X105Y89_OLOGIC_X1Y89_D1 = CLBLM_R_X11Y130_SLICE_X14Y130_AQ;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_A1 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_A2 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_A3 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_A4 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_A5 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_A6 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B4 = CLBLM_L_X8Y137_SLICE_X10Y137_B5Q;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_AX = LIOB33_X0Y209_IOB_X0Y210_I;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_B1 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_B2 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_B3 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_B4 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_B5 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_B6 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_BX = LIOB33_X0Y211_IOB_X0Y211_I;
  assign RIOI3_X105Y101_OLOGIC_X1Y102_D1 = CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_C1 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_C2 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_C3 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_C4 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_C5 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_C6 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign RIOI3_X105Y101_OLOGIC_X1Y102_T1 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_CX = LIOB33_X0Y211_IOB_X0Y212_I;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_D1 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_D2 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_D3 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_D4 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_D5 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_D6 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_DX = LIOB33_X0Y219_IOB_X0Y219_I;
  assign RIOI3_X105Y101_OLOGIC_X1Y101_D1 = CLBLM_R_X7Y126_SLICE_X8Y126_AQ;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_D1 = CLBLL_L_X54Y96_SLICE_X82Y96_AQ;
  assign RIOI3_X105Y101_OLOGIC_X1Y101_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_T1 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_A1 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_A2 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_A3 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_A4 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_A5 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_A6 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_D1 = CLBLM_R_X7Y137_SLICE_X9Y137_DQ;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_AX = LIOB33_X0Y203_IOB_X0Y204_I;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_B1 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_B2 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_B3 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_B4 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_B5 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_B6 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_T1 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_BX = LIOB33_X0Y209_IOB_X0Y209_I;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_C1 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_C2 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_C3 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_C4 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_C5 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_C6 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_D1 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_D2 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_D3 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_D4 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_D5 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_D6 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D3 = CLBLM_R_X3Y131_SLICE_X3Y131_DQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D5 = CLBLM_R_X3Y133_SLICE_X3Y133_BQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D6 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign RIOB33_X105Y161_IOB_X1Y162_O = CLBLM_L_X8Y132_SLICE_X11Y132_AQ;
  assign RIOB33_X105Y161_IOB_X1Y161_O = CLBLM_R_X5Y134_SLICE_X7Y134_AQ;
  assign LIOI3_X0Y177_ILOGIC_X0Y178_D = LIOB33_X0Y177_IOB_X0Y178_I;
  assign LIOI3_X0Y177_ILOGIC_X0Y177_D = LIOB33_X0Y177_IOB_X0Y177_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_D = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_D = LIOB33_X0Y55_IOB_X0Y55_I;
  assign LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y82_D = LIOB33_X0Y81_IOB_X0Y82_I;
  assign LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y81_D = LIOB33_X0Y81_IOB_X0Y81_I;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_ADDRARDADDR0 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_ADDRARDADDR1 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_ADDRARDADDR2 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_ADDRARDADDR3 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_ADDRARDADDR4 = CLBLM_R_X3Y139_SLICE_X2Y139_AO6;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_ADDRARDADDR5 = CLBLL_L_X4Y139_SLICE_X4Y139_BO6;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_ADDRARDADDR6 = CLBLL_L_X4Y139_SLICE_X5Y139_CO6;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_ADDRARDADDR7 = CLBLL_L_X4Y139_SLICE_X4Y139_AO6;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_ADDRARDADDR8 = CLBLM_R_X3Y138_SLICE_X3Y138_AO6;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_ADDRARDADDR9 = CLBLL_L_X4Y140_SLICE_X5Y140_BO6;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_ADDRARDADDR10 = CLBLM_R_X3Y138_SLICE_X2Y138_AO6;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_ADDRARDADDR11 = CLBLM_R_X5Y140_SLICE_X7Y140_AO6;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_ADDRARDADDR12 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_ADDRARDADDR13 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_ADDRATIEHIGH0 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_ADDRATIEHIGH1 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_ADDRBTIEHIGH0 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_ADDRBTIEHIGH1 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_ADDRBWRADDR0 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_ADDRBWRADDR1 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_ADDRBWRADDR2 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_ADDRBWRADDR3 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_ADDRBWRADDR4 = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_ADDRBWRADDR5 = CLBLM_R_X5Y140_SLICE_X6Y140_AO6;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_ADDRBWRADDR6 = CLBLM_R_X5Y140_SLICE_X6Y140_BO6;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_ADDRBWRADDR7 = CLBLM_R_X5Y139_SLICE_X7Y139_AO6;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_ADDRBWRADDR8 = CLBLM_R_X7Y140_SLICE_X8Y140_AO6;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_ADDRBWRADDR9 = CLBLM_R_X7Y140_SLICE_X8Y140_CO6;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_ADDRBWRADDR10 = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_ADDRBWRADDR11 = CLBLM_R_X5Y140_SLICE_X6Y140_CO6;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_ADDRBWRADDR12 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_ADDRBWRADDR13 = 1'b0;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_A1 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_A2 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_RDCLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_WRCLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_DIADI0 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_DIADI1 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_DIADI2 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_DIADI3 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_DIADI4 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_DIADI5 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_DIADI6 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_DIADI7 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_DIADI8 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_DIADI9 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_DIADI10 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_DIADI11 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_DIADI12 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_DIADI13 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_DIADI14 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_DIADI15 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_DIBDI0 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_DIBDI1 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_DIBDI2 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_DIBDI3 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_DIBDI4 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_DIBDI5 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_DIBDI6 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_DIBDI7 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_DIBDI8 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_DIBDI9 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_DIBDI10 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_DIBDI11 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_DIBDI12 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_DIBDI13 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_DIBDI14 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_DIBDI15 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_DIPADIP0 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_DIPADIP1 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_DIPBDIP0 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_DIPBDIP1 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_D4 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_D5 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_D6 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_DX = LIOB33_X0Y235_IOB_X0Y235_I;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_A1 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_A2 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_A3 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_A4 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_A5 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_A6 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_B1 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_B2 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_B3 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_B4 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_RDEN = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_WREN = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_B5 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_B6 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_C1 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_C2 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_C3 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_C4 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_C5 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_C6 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_REGCE = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_REGCEB = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_RDRCLK = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_REGCLKB = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_RST = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_D1 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_RSTRAMB = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_RSTREG = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_RSTREGB = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_WEA0 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_WEA1 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_WEA2 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_WEA3 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_WEBWE0 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_WEBWE1 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_WEBWE2 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_WEBWE3 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_WEBWE4 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_WEBWE5 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_WEBWE6 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y56_WEBWE7 = 1'b0;
  assign RIOB33_X105Y163_IOB_X1Y164_O = CLBLM_R_X7Y134_SLICE_X9Y134_AQ;
  assign RIOB33_X105Y163_IOB_X1Y163_O = CLBLM_L_X8Y135_SLICE_X10Y135_AQ;
  assign RIOB33_X105Y165_IOB_X1Y166_O = CLBLM_L_X8Y136_SLICE_X10Y136_AQ;
  assign RIOB33_X105Y165_IOB_X1Y165_O = CLBLM_R_X7Y134_SLICE_X9Y134_BQ;
  assign RIOI3_X105Y103_OLOGIC_X1Y103_D1 = CLBLM_R_X7Y126_SLICE_X8Y126_CQ;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_D1 = CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  assign RIOI3_X105Y103_OLOGIC_X1Y103_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_D1 = CLBLM_L_X10Y132_SLICE_X12Y132_DQ;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_T1 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X37Y149_A1 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X37Y149_A2 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X37Y149_A3 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X37Y149_A4 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X37Y149_A5 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X37Y149_A6 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X37Y149_AX = RIOB33_X105Y181_IOB_X1Y182_I;
  assign CLBLM_R_X25Y149_SLICE_X37Y149_B1 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X37Y149_B2 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X37Y149_B3 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X37Y149_B4 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X37Y149_B5 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X37Y149_B6 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X37Y149_C1 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X37Y149_C2 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X37Y149_C3 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X37Y149_C4 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X37Y149_C5 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X37Y149_C6 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X37Y149_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X25Y149_SLICE_X37Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X25Y149_SLICE_X37Y149_D1 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X37Y149_D2 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X37Y149_D3 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X37Y149_D4 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X37Y149_D5 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X37Y149_D6 = 1'b1;
  assign LIOI3_X0Y179_ILOGIC_X0Y180_D = LIOB33_X0Y179_IOB_X0Y180_I;
  assign RIOI3_TBYTETERM_X105Y187_ILOGIC_X1Y188_D = RIOB33_X105Y187_IOB_X1Y188_I;
  assign LIOI3_X0Y179_ILOGIC_X0Y179_D = LIOB33_X0Y179_IOB_X0Y179_I;
  assign CLBLM_R_X25Y149_SLICE_X36Y149_A1 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X36Y149_A2 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X36Y149_A3 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X36Y149_A4 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X36Y149_A5 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X36Y149_A6 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X36Y149_AX = RIOB33_X105Y179_IOB_X1Y179_I;
  assign RIOI3_TBYTETERM_X105Y187_ILOGIC_X1Y187_D = RIOB33_X105Y187_IOB_X1Y187_I;
  assign CLBLM_R_X25Y149_SLICE_X36Y149_B1 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X36Y149_B2 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X36Y149_B3 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X36Y149_B4 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X36Y149_B5 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X36Y149_B6 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X36Y149_BX = RIOB33_X105Y179_IOB_X1Y180_I;
  assign CLBLM_R_X25Y149_SLICE_X36Y149_C1 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X36Y149_C2 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X36Y149_C3 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X36Y149_C4 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X36Y149_C5 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X36Y149_C6 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X36Y149_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_D = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_D = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLM_R_X25Y149_SLICE_X36Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X25Y149_SLICE_X36Y149_D1 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X36Y149_D2 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X36Y149_D3 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X36Y149_D4 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X36Y149_D5 = 1'b1;
  assign CLBLM_R_X25Y149_SLICE_X36Y149_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y93_ILOGIC_X0Y94_D = LIOB33_X0Y93_IOB_X0Y94_I;
  assign LIOI3_TBYTESRC_X0Y93_ILOGIC_X0Y93_D = LIOB33_X0Y93_IOB_X0Y93_I;
  assign RIOB33_X105Y167_IOB_X1Y168_O = CLBLM_L_X8Y137_SLICE_X10Y137_AQ;
  assign RIOB33_X105Y167_IOB_X1Y167_O = CLBLM_L_X10Y135_SLICE_X12Y135_AQ;
  assign RIOB33_X105Y169_IOB_X1Y170_O = CLBLM_L_X56Y151_SLICE_X84Y151_AQ;
  assign RIOB33_X105Y169_IOB_X1Y169_O = CLBLM_L_X8Y137_SLICE_X10Y137_BQ;
  assign RIOI3_X105Y105_OLOGIC_X1Y106_D1 = CLBLM_R_X5Y131_SLICE_X7Y131_AQ;
  assign CLBLM_R_X25Y151_SLICE_X37Y151_A1 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X37Y151_A2 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X37Y151_A3 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X37Y151_A4 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X37Y151_A5 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X37Y151_A6 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X37Y151_B1 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X37Y151_B2 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X37Y151_B3 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X37Y151_B4 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X37Y151_B5 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X37Y151_B6 = 1'b1;
  assign RIOI3_X105Y105_OLOGIC_X1Y106_T1 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X37Y151_C1 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X37Y151_C2 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X37Y151_C3 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X37Y151_C4 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X37Y151_C5 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X37Y151_C6 = 1'b1;
  assign RIOI3_X105Y105_OLOGIC_X1Y105_D1 = CLBLM_R_X7Y129_SLICE_X9Y129_CQ;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_D1 = CLBLM_R_X7Y131_SLICE_X9Y131_DQ;
  assign RIOI3_X105Y105_OLOGIC_X1Y105_T1 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X37Y151_D1 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X37Y151_D2 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X37Y151_D3 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X37Y151_D4 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X37Y151_D5 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X37Y151_D6 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_T1 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X36Y151_A1 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X36Y151_A2 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X36Y151_A3 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X36Y151_A4 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X36Y151_A5 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X36Y151_A6 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_D1 = CLBLM_R_X7Y131_SLICE_X9Y131_CQ;
  assign CLBLM_R_X25Y151_SLICE_X36Y151_AX = RIOB33_X105Y183_IOB_X1Y184_I;
  assign CLBLM_R_X25Y151_SLICE_X36Y151_B1 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X36Y151_B2 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X36Y151_B3 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X36Y151_B4 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X36Y151_B5 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X36Y151_B6 = 1'b1;
  assign RIOB33_X105Y171_IOB_X1Y171_O = CLBLM_R_X15Y135_SLICE_X21Y135_AQ;
  assign RIOB33_X105Y171_IOB_X1Y172_O = CLBLM_L_X16Y136_SLICE_X22Y136_AQ;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_T1 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X36Y151_BX = RIOB33_X105Y187_IOB_X1Y188_I;
  assign CLBLM_R_X25Y151_SLICE_X36Y151_C1 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X36Y151_C2 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X36Y151_C3 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X36Y151_C4 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X36Y151_C5 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X36Y151_C6 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X36Y151_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X25Y151_SLICE_X36Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X25Y151_SLICE_X36Y151_CX = RIOB33_X105Y189_IOB_X1Y189_I;
  assign CLBLM_R_X25Y151_SLICE_X36Y151_D1 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X36Y151_D2 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X36Y151_D3 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X36Y151_D4 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X36Y151_D5 = 1'b1;
  assign CLBLM_R_X25Y151_SLICE_X36Y151_D6 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_ADDRARDADDR0 = 1'b0;
  assign LIOI3_X0Y183_ILOGIC_X0Y184_D = LIOB33_X0Y183_IOB_X0Y184_I;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_ADDRARDADDR1 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_ADDRARDADDR2 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_ADDRARDADDR3 = 1'b0;
  assign LIOI3_X0Y183_ILOGIC_X0Y183_D = LIOB33_X0Y183_IOB_X0Y183_I;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_ADDRARDADDR4 = CLBLL_L_X4Y140_SLICE_X4Y140_BO6;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_ADDRARDADDR5 = CLBLM_R_X3Y138_SLICE_X3Y138_CO6;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_ADDRARDADDR6 = CLBLL_L_X4Y140_SLICE_X4Y140_AO6;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_ADDRARDADDR7 = CLBLM_R_X3Y138_SLICE_X3Y138_BO6;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_ADDRARDADDR8 = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_ADDRARDADDR9 = CLBLL_L_X4Y139_SLICE_X5Y139_DO6;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_ADDRARDADDR10 = CLBLM_R_X5Y138_SLICE_X6Y138_DO6;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_ADDRARDADDR11 = CLBLM_R_X3Y138_SLICE_X3Y138_DO6;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_ADDRARDADDR12 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_ADDRARDADDR13 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_ADDRATIEHIGH0 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_ADDRATIEHIGH1 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_ADDRBTIEHIGH0 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_ADDRBTIEHIGH1 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_ADDRBWRADDR0 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_ADDRBWRADDR1 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_ADDRBWRADDR2 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_ADDRBWRADDR3 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_ADDRBWRADDR4 = CLBLL_L_X4Y139_SLICE_X4Y139_DO6;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_ADDRBWRADDR5 = CLBLM_R_X7Y139_SLICE_X8Y139_AO6;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_ADDRBWRADDR6 = CLBLM_R_X7Y140_SLICE_X8Y140_DO6;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_ADDRBWRADDR8 = CLBLM_R_X7Y140_SLICE_X8Y140_BO6;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_ADDRBWRADDR9 = CLBLM_R_X7Y138_SLICE_X8Y138_DO6;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_ADDRBWRADDR10 = CLBLM_R_X5Y139_SLICE_X7Y139_DO6;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_ADDRBWRADDR11 = CLBLM_R_X5Y140_SLICE_X6Y140_DO6;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_ADDRBWRADDR12 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_ADDRBWRADDR13 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_ADDRBWRADDR7 = CLBLM_R_X5Y138_SLICE_X7Y138_CO6;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_D = LIOB33_X0Y61_IOB_X0Y62_I;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_CLKARDCLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_CLKBWRCLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_D = LIOB33_X0Y61_IOB_X0Y61_I;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_DIADI0 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_DIADI1 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_DIADI2 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_DIADI3 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_DIADI4 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_DIADI5 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_DIADI6 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_DIADI7 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_DIADI8 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_DIADI9 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_DIADI10 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_DIADI11 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_DIADI12 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_DIADI13 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_DIADI14 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_DIADI15 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_DIBDI0 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_DIBDI1 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_DIBDI2 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_DIBDI3 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_DIBDI4 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_DIBDI5 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_DIBDI6 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_DIBDI7 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_DIBDI8 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_DIBDI9 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_DIBDI10 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_DIBDI11 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_DIBDI12 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_DIBDI13 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_DIBDI14 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_DIBDI15 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_DIPADIP0 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_DIPADIP1 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_DIPBDIP0 = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_DIPBDIP1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D = LIOB33_X0Y107_IOB_X0Y107_I;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_ENARDEN = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_ENBWREN = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_REGCEAREGCE = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_REGCEB = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_REGCLKARDRCLK = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_REGCLKB = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_RSTRAMARSTRAM = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_RSTRAMB = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_RSTREGARSTREG = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_RSTREGB = 1'b1;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_WEA0 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_WEA1 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_WEA2 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_WEA3 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_WEBWE0 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_WEBWE1 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_WEBWE2 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_WEBWE3 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_WEBWE4 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_WEBWE5 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_WEBWE6 = 1'b0;
  assign BRAM_L_X6Y140_RAMB18_X0Y57_WEBWE7 = 1'b0;
  assign RIOB33_X105Y173_IOB_X1Y174_O = CLBLM_L_X16Y135_SLICE_X22Y135_BQ;
  assign RIOB33_X105Y173_IOB_X1Y173_O = CLBLM_L_X16Y135_SLICE_X22Y135_AQ;
  assign CLBLM_L_X16Y149_SLICE_X23Y149_A1 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X23Y149_A2 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X23Y149_A3 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X23Y149_A4 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X23Y149_A5 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X23Y149_A6 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X23Y149_B1 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X23Y149_B2 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X23Y149_B3 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X23Y149_B4 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X23Y149_B5 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X23Y149_B6 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X23Y149_C1 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X23Y149_C2 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X23Y149_C3 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X23Y149_C4 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X23Y149_C5 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X23Y149_C6 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X23Y149_D1 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X23Y149_D2 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X23Y149_D3 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X23Y149_D4 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X23Y149_D5 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X23Y149_D6 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X22Y149_A1 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X22Y149_A2 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X22Y149_A3 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X22Y149_A4 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X22Y149_A5 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X22Y149_A6 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X22Y149_AX = RIOB33_X105Y177_IOB_X1Y178_I;
  assign CLBLM_L_X16Y149_SLICE_X22Y149_B1 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X22Y149_B2 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X22Y149_B3 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X22Y149_B4 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X22Y149_B5 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X22Y149_B6 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X22Y149_BX = RIOB33_X105Y181_IOB_X1Y181_I;
  assign CLBLM_L_X16Y149_SLICE_X22Y149_C1 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X22Y149_C2 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X22Y149_C3 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X22Y149_C4 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X22Y149_C5 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X22Y149_C6 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X22Y149_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_L_X16Y149_SLICE_X22Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y149_SLICE_X22Y149_D1 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X22Y149_D2 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X22Y149_D3 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X22Y149_D4 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X22Y149_D5 = 1'b1;
  assign CLBLM_L_X16Y149_SLICE_X22Y149_D6 = 1'b1;
  assign RIOB33_X105Y175_IOB_X1Y176_O = CLBLM_L_X16Y137_SLICE_X22Y137_AQ;
  assign RIOB33_X105Y175_IOB_X1Y175_O = CLBLM_R_X13Y136_SLICE_X18Y136_AQ;
  assign CLBLM_R_X25Y153_SLICE_X37Y153_A1 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X37Y153_A2 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X37Y153_A3 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X37Y153_A4 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X37Y153_A5 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X37Y153_A6 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X37Y153_B1 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X37Y153_B2 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X37Y153_B3 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X37Y153_B4 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X37Y153_B5 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X37Y153_B6 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X37Y153_C1 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X37Y153_C2 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X37Y153_C3 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X37Y153_C4 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X37Y153_C5 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X37Y153_C6 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X37Y153_D1 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X37Y153_D2 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X37Y153_D3 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X37Y153_D4 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X37Y153_D5 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X37Y153_D6 = 1'b1;
  assign CLK_HROW_BOT_R_X139Y78_BUFHCE_X0Y20_CE = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X36Y153_A1 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X36Y153_A2 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X36Y153_A3 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X36Y153_A4 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X36Y153_A5 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X36Y153_A6 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X36Y153_AX = RIOB33_X105Y195_IOB_X1Y195_I;
  assign CLBLM_R_X25Y153_SLICE_X36Y153_B1 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X36Y153_B2 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X36Y153_B3 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X36Y153_B4 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X36Y153_B5 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X36Y153_B6 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X36Y153_BX = RIOB33_X105Y195_IOB_X1Y196_I;
  assign CLBLM_R_X25Y153_SLICE_X36Y153_C1 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X36Y153_C2 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X36Y153_C3 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X36Y153_C4 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X36Y153_C5 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X36Y153_C6 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X36Y153_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X25Y153_SLICE_X36Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X25Y153_SLICE_X36Y153_D1 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X36Y153_D2 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X36Y153_D3 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X36Y153_D4 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X36Y153_D5 = 1'b1;
  assign CLBLM_R_X25Y153_SLICE_X36Y153_D6 = 1'b1;
  assign RIOI3_X105Y109_OLOGIC_X1Y110_D1 = CLBLM_R_X7Y129_SLICE_X8Y129_DQ;
  assign RIOI3_X105Y109_OLOGIC_X1Y110_T1 = 1'b1;
  assign RIOI3_X105Y109_OLOGIC_X1Y109_D1 = CLBLM_R_X7Y129_SLICE_X8Y129_CQ;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_D1 = CLBLM_R_X7Y137_SLICE_X8Y137_BQ;
  assign RIOI3_X105Y109_OLOGIC_X1Y109_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_D1 = CLBLM_R_X5Y137_SLICE_X7Y137_AQ;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_T1 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A1 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A2 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A3 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A4 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A5 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A6 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B1 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B2 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B3 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B4 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B5 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B6 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C1 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C2 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C3 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C4 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C5 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C6 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D1 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D2 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D3 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D4 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D5 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D6 = 1'b1;
  assign LIOI3_X0Y185_ILOGIC_X0Y186_D = LIOB33_X0Y185_IOB_X0Y186_I;
  assign LIOI3_X0Y185_ILOGIC_X0Y185_D = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A1 = BRAM_R_X17Y135_RAMB18_X1Y54_DO16;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A2 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A3 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A4 = CLBLM_R_X3Y131_SLICE_X3Y131_BQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A5 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A6 = 1'b1;
  assign RIOB33_X105Y177_IOB_X1Y177_O = CLBLM_L_X16Y137_SLICE_X22Y137_BQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B1 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B2 = CLBLM_R_X3Y131_SLICE_X3Y131_CQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B3 = BRAM_R_X17Y135_RAMB18_X1Y54_DO18;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B4 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B5 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B6 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C1 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C2 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C3 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C4 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C5 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C6 = 1'b1;
  assign LIOI3_X0Y65_ILOGIC_X0Y66_D = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y65_D = LIOB33_X0Y65_IOB_X0Y65_I;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D1 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D2 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D3 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D4 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D5 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D6 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X37Y154_A1 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X37Y154_A2 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X37Y154_A3 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X37Y154_A4 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X37Y154_A5 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X37Y154_A6 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X37Y154_B1 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X37Y154_B2 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X37Y154_B3 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X37Y154_B4 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X37Y154_B5 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X37Y154_B6 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X37Y154_C1 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X37Y154_C2 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X37Y154_C3 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X37Y154_C4 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X37Y154_C5 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X37Y154_C6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_D = LIOB33_X0Y119_IOB_X0Y120_I;
  assign LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y119_D = LIOB33_X0Y119_IOB_X0Y119_I;
  assign CLBLM_R_X25Y154_SLICE_X37Y154_D1 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X37Y154_D2 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X37Y154_D3 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X37Y154_D4 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X37Y154_D5 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X37Y154_D6 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X36Y154_A1 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X36Y154_A2 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X36Y154_A3 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X36Y154_A4 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X36Y154_A5 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X36Y154_A6 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X36Y154_AX = RIOB33_SING_X105Y200_IOB_X1Y200_I;
  assign CLBLM_R_X25Y154_SLICE_X36Y154_B1 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X36Y154_B2 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X36Y154_B3 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X36Y154_B4 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X36Y154_B5 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X36Y154_B6 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B5 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B6 = CLBLM_R_X7Y132_SLICE_X8Y132_CQ;
  assign CLBLM_R_X25Y154_SLICE_X36Y154_BX = RIOB33_X105Y197_IOB_X1Y198_I;
  assign CLBLM_R_X25Y154_SLICE_X36Y154_C1 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X36Y154_C2 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X36Y154_C3 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X36Y154_C4 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X36Y154_C5 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X36Y154_C6 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X36Y154_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X25Y154_SLICE_X36Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X25Y154_SLICE_X36Y154_CX = RIOB33_SING_X105Y199_IOB_X1Y199_I;
  assign CLBLM_R_X25Y154_SLICE_X36Y154_D1 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X36Y154_D2 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X36Y154_D3 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X36Y154_D4 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X36Y154_D5 = 1'b1;
  assign CLBLM_R_X25Y154_SLICE_X36Y154_D6 = 1'b1;
  assign CLK_HROW_BOT_R_X139Y78_BUFHCE_X0Y20_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C2 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C3 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C5 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_A1 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_A2 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_A3 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_A4 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_A5 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_A6 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D4 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_AX = RIOB33_X105Y183_IOB_X1Y183_I;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D5 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_B1 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_B2 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_B3 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_B4 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_B5 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_B6 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D6 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_C1 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A1 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A2 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A3 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_C5 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_C6 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A4 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A5 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A6 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_C2 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_C3 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B1 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B2 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_D1 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_D2 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_D3 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_D4 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_D5 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_D6 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B3 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B4 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B5 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B6 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A1 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_A1 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_A2 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_A3 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_A4 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_A5 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_A6 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C5 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C6 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_AX = RIOB33_X105Y185_IOB_X1Y185_I;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B1 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_B1 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_B2 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_B3 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D1 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_B6 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D2 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D3 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D4 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D5 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D6 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_C1 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_C2 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C5 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_C5 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_BX = RIOB33_X105Y185_IOB_X1Y186_I;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D1 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D2 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D3 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D4 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D5 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D6 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_D1 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_D2 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_D3 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_D4 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_D5 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_D6 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_CX = RIOB33_X105Y187_IOB_X1Y187_I;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A1 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A2 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_DX = RIOB33_X105Y191_IOB_X1Y191_I;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A3 = CLBLM_R_X5Y130_SLICE_X6Y130_DQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A1 = CLBLL_L_X4Y127_SLICE_X5Y127_AQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A2 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A3 = CLBLM_R_X7Y129_SLICE_X9Y129_B5Q;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A4 = BRAM_L_X6Y125_RAMB18_X0Y50_DO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A5 = LIOB33_X0Y19_IOB_X0Y20_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A6 = CLBLM_R_X5Y127_SLICE_X6Y127_B5Q;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B1 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B1 = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B2 = CLBLL_L_X4Y128_SLICE_X5Y128_BQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B3 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B4 = BRAM_L_X6Y125_RAMB18_X0Y50_DO7;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B5 = CLBLM_R_X5Y127_SLICE_X7Y127_DQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B6 = CLBLL_L_X4Y128_SLICE_X5Y128_AO5;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C1 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C1 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C2 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C3 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C4 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C5 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C6 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C4 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C5 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C6 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D1 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D2 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D3 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D4 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D5 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D6 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D5 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D1 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D2 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D3 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D4 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D6 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_B2 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_B5 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_A1 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_A2 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_A3 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_A4 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_A5 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_A6 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_B1 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_B2 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_B3 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_B4 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_C1 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_B5 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_B6 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_C2 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_C1 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_C2 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_C3 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_C4 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_C5 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_C6 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_C5 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_D1 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_D2 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_D3 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_D4 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_D5 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_D6 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_A1 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_A2 = CLBLM_R_X25Y157_SLICE_X37Y157_AQ;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_A3 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_A4 = CLBLM_R_X3Y133_SLICE_X3Y133_AQ;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_A5 = CLBLM_L_X10Y135_SLICE_X12Y135_BO6;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_A6 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_B1 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_B2 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_B3 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_B4 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_B5 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_B6 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_C1 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_C2 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_C3 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_C4 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_C5 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_C6 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_D1 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_D2 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_D3 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_D4 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_D5 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_D6 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_D6 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_A1 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_A2 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_A3 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_A4 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_A5 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_A6 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_B1 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_B2 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_B3 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_B4 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_B5 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_B6 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_A1 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_A2 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_A3 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_A4 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_C1 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_C2 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_C3 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_C4 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_A5 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_C6 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_A6 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_B1 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_B2 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_B3 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_B4 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_B5 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_B6 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_D1 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_D2 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_D3 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_D4 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_D5 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_D6 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_C1 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_C2 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_C3 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_C4 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A1 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_A1 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_A2 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_A3 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_A4 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_A5 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_A6 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A6 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_AX = RIOB33_X105Y189_IOB_X1Y190_I;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B1 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_B1 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_B2 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_B3 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_B4 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_B5 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_B6 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_D6 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C1 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C2 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C3 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C4 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C5 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C6 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_BX = RIOB33_X105Y191_IOB_X1Y192_I;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_C1 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_C2 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_C3 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D1 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D2 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D3 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D4 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D5 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_D1 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_D2 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_D3 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A2 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_D4 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_D5 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_D6 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_A1 = BRAM_L_X6Y125_RAMB18_X0Y50_DO7;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_A2 = CLBLM_L_X8Y130_SLICE_X10Y130_A5Q;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_A3 = CLBLL_L_X4Y128_SLICE_X5Y128_AQ;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_A4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A3 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A4 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A5 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A6 = BRAM_L_X6Y135_RAMB18_X0Y54_DO20;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B1 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B2 = CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B3 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO4;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B4 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B5 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B6 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_C4 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C1 = CLBLM_R_X5Y132_SLICE_X6Y132_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C2 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C3 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C4 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C5 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C6 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO5;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_C5 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_C6 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_D1 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_D2 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_D3 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_D4 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_D5 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_D6 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D1 = CLBLL_L_X4Y133_SLICE_X5Y133_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D2 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D3 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO7;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D4 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D5 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D6 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_A1 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_A2 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_A3 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_A4 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_A5 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_A6 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_B1 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_B2 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_B3 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_B4 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_B5 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_B6 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_C1 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_C2 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_C3 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_C4 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_C5 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_C6 = 1'b1;
  assign LIOI3_X0Y189_ILOGIC_X0Y190_D = LIOB33_X0Y189_IOB_X0Y190_I;
  assign LIOI3_X0Y189_ILOGIC_X0Y189_D = LIOB33_X0Y189_IOB_X0Y189_I;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_D1 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_D2 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_D3 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_D4 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_D5 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_D6 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_D4 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_A1 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_A2 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_A3 = BRAM_R_X17Y135_RAMB18_X1Y54_DO5;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_D5 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_A4 = CLBLM_R_X3Y133_SLICE_X3Y133_AQ;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_A5 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_A6 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_D6 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_A1 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_A2 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_A3 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_A4 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_A5 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_A6 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_B5 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_B1 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_B2 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_B3 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_B4 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_B5 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_B6 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_B6 = CLBLM_R_X11Y136_SLICE_X14Y136_CO6;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_C5 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_C1 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_C2 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_C3 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_C4 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_C5 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_C6 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_C6 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_D1 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_D2 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_D3 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_D4 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_D5 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y132_D = LIOB33_X0Y131_IOB_X0Y132_I;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_D1 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_D2 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_D3 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_D4 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_D5 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_D6 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y131_D = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_A1 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_A2 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_A3 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_A4 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_A5 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_A6 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_AX = LIOB33_X0Y229_IOB_X0Y230_I;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_B1 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_B2 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_B3 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_B4 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_B5 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_B6 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_BX = LIOB33_X0Y233_IOB_X0Y233_I;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_C1 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_C2 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_C3 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_C4 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_C5 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_C6 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_CX = LIOB33_X0Y239_IOB_X0Y239_I;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_D1 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_D2 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_D3 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_D4 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_D5 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_D6 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_A1 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_A2 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_A3 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_A4 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_A5 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_A6 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_DX = LIOB33_X0Y241_IOB_X0Y241_I;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_B1 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A1 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A2 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_B4 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_B5 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_B6 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A3 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A4 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A5 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A6 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_B2 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_AX = CLBLL_L_X4Y129_SLICE_X5Y129_BO6;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_C3 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_C4 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_C5 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_C6 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B1 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B2 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B3 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B4 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B5 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B6 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C1 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C2 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C3 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_D2 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_D3 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_D4 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_D5 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_D6 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C4 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C5 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C6 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A1 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO0;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A2 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_A1 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_A2 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_A3 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_A4 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_A5 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_A6 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A6 = CLBLM_R_X5Y130_SLICE_X6Y130_CQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D1 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D2 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_AX = RIOB33_X105Y193_IOB_X1Y193_I;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D4 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D5 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_B2 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B4 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO4;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B5 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_B6 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C1 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C2 = CLBLM_R_X5Y132_SLICE_X7Y132_A5Q;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C3 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C5 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_C1 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_C2 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_C3 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_C4 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_C5 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_C6 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D1 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D2 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D3 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D4 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D5 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_D1 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_D2 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_D3 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_D4 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_D5 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_D6 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A3 = CLBLL_L_X4Y129_SLICE_X5Y129_AQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A6 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A5 = CLBLM_R_X7Y129_SLICE_X8Y129_B5Q;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A1 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A2 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B1 = CLBLM_R_X7Y136_SLICE_X8Y136_A5Q;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B2 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B3 = LIOB33_X0Y73_IOB_X0Y73_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B4 = BRAM_L_X6Y125_RAMB18_X0Y50_DO17;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B5 = CLBLL_L_X4Y129_SLICE_X4Y129_AQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B6 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B1 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C1 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C2 = BRAM_L_X6Y125_RAMB18_X0Y50_DO18;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B5 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C3 = LIOB33_X0Y23_IOB_X0Y24_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C4 = CLBLL_L_X4Y129_SLICE_X5Y129_AQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C5 = CLBLL_L_X4Y129_SLICE_X5Y129_CQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C6 = CLBLM_R_X7Y129_SLICE_X8Y129_B5Q;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C1 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C2 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C3 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C4 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D1 = CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D2 = BRAM_L_X6Y125_RAMB18_X0Y50_DO18;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D3 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D4 = CLBLL_L_X4Y129_SLICE_X5Y129_AO5;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D5 = CLBLL_L_X4Y129_SLICE_X5Y129_CQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D6 = LIOB33_X0Y9_IOB_X0Y9_I;
  assign CLBLM_R_X25Y157_SLICE_X37Y157_A5 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X37Y157_A6 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D1 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D2 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D3 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D4 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D5 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D6 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X37Y157_B2 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X37Y157_B3 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X37Y157_B4 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X37Y157_B5 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X37Y157_B6 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X37Y157_B1 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X37Y157_C1 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X37Y157_C2 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X37Y157_C3 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X37Y157_C4 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X37Y157_C5 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X37Y157_C6 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X37Y157_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X25Y157_SLICE_X37Y157_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X25Y157_SLICE_X37Y157_D1 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X37Y157_D2 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X37Y157_D3 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X37Y157_D4 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X37Y157_D5 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X37Y157_D6 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X36Y157_A1 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X36Y157_A2 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X36Y157_A3 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X36Y157_A4 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X36Y157_A5 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X36Y157_A6 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X36Y157_AX = RIOB33_X105Y201_IOB_X1Y201_I;
  assign CLBLM_R_X25Y157_SLICE_X36Y157_B1 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X36Y157_B2 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X36Y157_B3 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X36Y157_B4 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X36Y157_B5 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X36Y157_B6 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X36Y157_BX = RIOB33_X105Y203_IOB_X1Y204_I;
  assign CLBLM_R_X25Y157_SLICE_X36Y157_C1 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X36Y157_C2 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X36Y157_C3 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X36Y157_C4 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X36Y157_C5 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X36Y157_C6 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X36Y157_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X25Y157_SLICE_X36Y157_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X25Y157_SLICE_X36Y157_D1 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X36Y157_D2 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X36Y157_D3 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X36Y157_D4 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X36Y157_D5 = 1'b1;
  assign CLBLM_R_X25Y157_SLICE_X36Y157_D6 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_A1 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_A2 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_A3 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_A4 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_A5 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_A6 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A1 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A2 = CLBLM_L_X8Y135_SLICE_X10Y135_A5Q;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A3 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A4 = BRAM_L_X6Y130_RAMB18_X0Y52_DO1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A5 = CLBLL_L_X4Y131_SLICE_X4Y131_AQ;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_B2 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_B3 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A6 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_B6 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_B1 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B1 = CLBLM_L_X8Y135_SLICE_X10Y135_A5Q;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B2 = CLBLL_L_X4Y130_SLICE_X4Y130_BQ;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_C1 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_C2 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_C3 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B3 = CLBLL_L_X4Y131_SLICE_X4Y131_AQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B4 = BRAM_L_X6Y130_RAMB18_X0Y52_DO1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_C6 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B5 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B6 = LIOB33_X0Y31_IOB_X0Y31_I;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C2 = BRAM_L_X6Y130_RAMB18_X0Y52_DO2;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C3 = CLBLL_L_X4Y131_SLICE_X4Y131_BO5;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C4 = CLBLM_R_X5Y130_SLICE_X6Y130_DQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C5 = CLBLL_L_X4Y131_SLICE_X4Y131_DQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C6 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_D1 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_D4 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_D5 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_D6 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_D2 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_D3 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A4 = BRAM_L_X6Y135_RAMB18_X0Y54_DO4;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A5 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO4;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A6 = CLBLM_R_X7Y129_SLICE_X9Y129_A5Q;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A1 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO3;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_A2 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D1 = CLBLM_R_X3Y130_SLICE_X3Y130_BQ;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_A4 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_A5 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_A6 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D5 = CLBLM_R_X3Y130_SLICE_X3Y130_AO5;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D6 = BRAM_L_X6Y125_RAMB18_X0Y50_DO21;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B1 = CLBLM_L_X16Y149_SLICE_X22Y149_AQ;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B2 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B3 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO7;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B4 = BRAM_R_X17Y135_RAMB18_X1Y54_DO7;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B5 = CLBLM_L_X10Y134_SLICE_X13Y134_AO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B6 = CLBLM_R_X7Y129_SLICE_X9Y129_A5Q;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_B6 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C1 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C2 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C3 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C4 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C5 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_C1 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_C2 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_C3 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_C4 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_C5 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_C6 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D2 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D3 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D1 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A1 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A2 = CLBLM_R_X3Y131_SLICE_X3Y131_CQ;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_D1 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_D2 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_D3 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A2 = BRAM_L_X6Y135_RAMB18_X0Y54_DO3;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A3 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO2;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A4 = BRAM_R_X17Y135_RAMB18_X1Y54_DO3;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A5 = BRAM_L_X6Y135_RAMB18_X0Y54_DO2;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_D4 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_D5 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_D6 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B3 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B4 = CLBLL_L_X4Y130_SLICE_X4Y130_BQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B5 = CLBLM_R_X7Y130_SLICE_X8Y130_B5Q;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B6 = LIOB33_X0Y15_IOB_X0Y16_I;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A6 = CLBLM_R_X7Y134_SLICE_X9Y134_B5Q;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_BX = CLBLL_L_X4Y130_SLICE_X5Y130_DO6;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_DIADI1 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B6 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C1 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C2 = CLBLL_L_X4Y131_SLICE_X5Y131_CQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C3 = CLBLL_L_X4Y131_SLICE_X5Y131_AO5;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C5 = LIOB33_X0Y13_IOB_X0Y13_I;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C6 = CLBLM_R_X5Y130_SLICE_X6Y130_B5Q;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B5 = CLBLM_L_X10Y134_SLICE_X12Y134_AO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C1 = CLBLM_R_X3Y131_SLICE_X3Y131_CQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D1 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D2 = CLBLM_R_X3Y131_SLICE_X3Y131_AO5;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D5 = CLBLL_L_X4Y130_SLICE_X5Y130_AQ;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_DIADI2 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D6 = CLBLM_R_X3Y131_SLICE_X3Y131_CQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C6 = CLBLM_L_X8Y134_SLICE_X10Y134_BO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D1 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D2 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D3 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D4 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D5 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D6 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_DIADI3 = 1'b1;
  assign RIOI3_X105Y115_OLOGIC_X1Y116_D1 = CLBLM_L_X10Y133_SLICE_X13Y133_AQ;
  assign RIOI3_X105Y115_OLOGIC_X1Y116_T1 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_DIADI4 = 1'b1;
  assign RIOI3_X105Y115_OLOGIC_X1Y115_D1 = CLBLL_L_X54Y123_SLICE_X82Y123_AQ;
  assign RIOI3_X105Y115_OLOGIC_X1Y115_T1 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_DIADI7 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_DIADI8 = 1'b0;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_DIADI9 = 1'b0;
  assign LIOI3_X0Y191_ILOGIC_X0Y192_D = LIOB33_X0Y191_IOB_X0Y192_I;
  assign LIOI3_X0Y191_ILOGIC_X0Y191_D = LIOB33_X0Y191_IOB_X0Y191_I;
  assign CLBLM_L_X16Y155_SLICE_X23Y155_A1 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A1 = LIOB33_X0Y75_IOB_X0Y76_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A2 = BRAM_L_X6Y125_RAMB18_X0Y50_DO20;
  assign CLBLM_L_X16Y155_SLICE_X23Y155_A4 = 1'b1;
  assign CLBLM_L_X16Y155_SLICE_X23Y155_A5 = 1'b1;
  assign CLBLM_L_X16Y155_SLICE_X23Y155_A6 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A3 = CLBLM_R_X7Y132_SLICE_X8Y132_A5Q;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A5 = CLBLL_L_X4Y131_SLICE_X5Y131_AQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A6 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_DIADI10 = 1'b0;
  assign CLBLM_L_X16Y155_SLICE_X23Y155_B2 = 1'b1;
  assign CLBLM_L_X16Y155_SLICE_X23Y155_B3 = 1'b1;
  assign CLBLM_L_X16Y155_SLICE_X23Y155_B4 = 1'b1;
  assign CLBLM_L_X16Y155_SLICE_X23Y155_B5 = 1'b1;
  assign CLBLM_L_X16Y155_SLICE_X23Y155_B6 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_AX = CLBLL_L_X4Y130_SLICE_X4Y130_AO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B1 = CLBLM_R_X7Y134_SLICE_X9Y134_A5Q;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B2 = CLBLL_L_X4Y131_SLICE_X4Y131_BQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B3 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B4 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B5 = BRAM_L_X6Y130_RAMB18_X0Y52_DO2;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B6 = 1'b1;
  assign LIOI3_X0Y71_ILOGIC_X0Y72_D = LIOB33_X0Y71_IOB_X0Y72_I;
  assign CLBLM_L_X16Y155_SLICE_X23Y155_C1 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C1 = CLBLL_L_X4Y132_SLICE_X4Y132_AQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C2 = CLBLL_L_X4Y131_SLICE_X4Y131_CQ;
  assign LIOI3_X0Y71_ILOGIC_X0Y71_D = LIOB33_X0Y71_IOB_X0Y71_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C3 = LIOB33_X0Y89_IOB_X0Y89_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C4 = BRAM_L_X6Y130_RAMB18_X0Y52_DO17;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C5 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C6 = CLBLM_R_X3Y131_SLICE_X2Y131_AQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y155_SLICE_X23Y155_D1 = 1'b1;
  assign CLBLM_L_X16Y155_SLICE_X23Y155_D2 = 1'b1;
  assign CLBLM_L_X16Y155_SLICE_X23Y155_D3 = 1'b1;
  assign CLBLM_L_X16Y155_SLICE_X23Y155_D4 = 1'b1;
  assign CLBLM_L_X16Y155_SLICE_X23Y155_D5 = 1'b1;
  assign CLBLM_L_X16Y155_SLICE_X23Y155_D6 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D1 = BRAM_L_X6Y130_RAMB18_X0Y52_DO2;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D2 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D3 = CLBLL_L_X4Y131_SLICE_X4Y131_DQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D5 = CLBLM_R_X7Y134_SLICE_X9Y134_A5Q;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D6 = CLBLL_L_X4Y131_SLICE_X4Y131_BQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A4 = BRAM_L_X6Y135_RAMB18_X0Y54_DO4;
  assign CLBLM_L_X16Y155_SLICE_X22Y155_A4 = 1'b1;
  assign CLBLM_L_X16Y155_SLICE_X22Y155_A5 = 1'b1;
  assign CLBLM_L_X16Y155_SLICE_X22Y155_A6 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_DIADI12 = 1'b0;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B1 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B2 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO0;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B3 = CLBLL_L_X4Y132_SLICE_X4Y132_AQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B4 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B5 = BRAM_R_X17Y135_RAMB18_X1Y54_DO0;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B6 = BRAM_L_X6Y135_RAMB18_X0Y54_DO1;
  assign CLBLM_L_X16Y155_SLICE_X22Y155_B5 = 1'b1;
  assign CLBLM_L_X16Y155_SLICE_X22Y155_B6 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C1 = BRAM_L_X6Y135_RAMB18_X0Y54_DO2;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C2 = BRAM_L_X6Y135_RAMB18_X0Y54_DO1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C3 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C4 = BRAM_R_X17Y135_RAMB18_X1Y54_DO2;
  assign CLBLM_L_X16Y155_SLICE_X22Y155_C1 = 1'b1;
  assign CLBLM_L_X16Y155_SLICE_X22Y155_C2 = 1'b1;
  assign CLBLM_L_X16Y155_SLICE_X22Y155_C3 = 1'b1;
  assign CLBLM_L_X16Y155_SLICE_X22Y155_C4 = 1'b1;
  assign CLBLM_L_X16Y155_SLICE_X22Y155_C5 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A1 = CLBLL_L_X4Y131_SLICE_X5Y131_B5Q;
  assign CLBLM_L_X16Y155_SLICE_X22Y155_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D3 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A2 = CLBLM_R_X7Y137_SLICE_X8Y137_A5Q;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_D = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D6 = BRAM_L_X6Y135_RAMB18_X0Y54_DO0;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A3 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A4 = BRAM_L_X6Y125_RAMB18_X0Y50_DO22;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A5 = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A6 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_AX = CLBLL_L_X4Y131_SLICE_X4Y131_AO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B1 = LIOB33_X0Y25_IOB_X0Y26_I;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B2 = CLBLL_L_X4Y131_SLICE_X5Y131_BQ;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B3 = CLBLL_L_X4Y131_SLICE_X5Y131_AQ;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B4 = BRAM_L_X6Y125_RAMB18_X0Y50_DO20;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A3 = BRAM_L_X6Y130_RAMB18_X0Y52_DO5;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B5 = CLBLM_R_X7Y132_SLICE_X8Y132_A5Q;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B6 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_BX = CLBLL_L_X4Y131_SLICE_X5Y131_AO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C1 = LIOB33_X0Y27_IOB_X0Y28_I;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C2 = CLBLL_L_X4Y131_SLICE_X5Y131_CQ;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C3 = BRAM_L_X6Y125_RAMB18_X0Y50_DO22;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C5 = CLBLL_L_X4Y131_SLICE_X5Y131_B5Q;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C6 = CLBLM_R_X7Y137_SLICE_X8Y137_A5Q;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B2 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO5;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B3 = CLBLM_R_X3Y133_SLICE_X3Y133_AQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B4 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO4;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B1 = BRAM_R_X17Y135_RAMB18_X1Y54_DO4;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D1 = CLBLL_L_X4Y128_SLICE_X5Y128_AQ;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D2 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D3 = CLBLM_R_X3Y157_SLICE_X3Y157_DQ;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D4 = CLBLM_R_X5Y131_SLICE_X7Y131_DO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D5 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D6 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B6 = BRAM_L_X6Y135_RAMB18_X0Y54_DO5;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C1 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO2;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C2 = CLBLM_R_X5Y130_SLICE_X6Y130_AQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C3 = BRAM_R_X17Y135_RAMB18_X1Y54_DO2;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C4 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO3;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C5 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO3;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C6 = BRAM_L_X6Y135_RAMB18_X0Y54_DO3;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D1 = BRAM_L_X6Y135_RAMB18_X0Y54_DO4;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D2 = BRAM_L_X6Y135_RAMB18_X0Y54_DO5;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D3 = BRAM_R_X17Y135_RAMB18_X1Y54_DO5;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D4 = CLBLM_L_X10Y135_SLICE_X12Y135_A5Q;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D5 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO5;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D6 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO4;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A1 = LIOB33_X0Y141_IOB_X0Y141_I;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A2 = BRAM_L_X6Y130_RAMB18_X0Y52_DO17;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A3 = CLBLL_L_X4Y132_SLICE_X4Y132_AQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A4 = CLBLM_R_X3Y131_SLICE_X2Y131_AQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A5 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A6 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B1 = BRAM_L_X6Y130_RAMB18_X0Y52_DO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B2 = CLBLL_L_X4Y132_SLICE_X4Y132_BQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B3 = LIOB33_X0Y85_IOB_X0Y86_I;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B4 = CLBLM_L_X8Y137_SLICE_X10Y137_A5Q;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B5 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B6 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C1 = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C2 = CLBLL_L_X4Y132_SLICE_X4Y132_CQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C3 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C4 = CLBLL_L_X4Y132_SLICE_X4Y132_AO5;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C5 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C6 = CLBLL_L_X4Y131_SLICE_X4Y131_CQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D2 = CLBLL_L_X4Y132_SLICE_X4Y132_BO5;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D3 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D4 = CLBLL_L_X4Y133_SLICE_X4Y133_AQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D5 = BRAM_L_X6Y130_RAMB18_X0Y52_DO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D6 = CLBLM_R_X5Y132_SLICE_X7Y132_A5Q;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A1 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO7;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A2 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A3 = BRAM_L_X6Y135_RAMB18_X0Y54_DO7;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A4 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO7;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A5 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A6 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B1 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO0;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B2 = BRAM_R_X17Y135_RAMB18_X1Y54_DO0;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B3 = CLBLM_R_X3Y131_SLICE_X3Y131_AQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B4 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B5 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B6 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C1 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO2;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C2 = BRAM_R_X17Y135_RAMB18_X1Y54_DO1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C3 = CLBLM_R_X3Y131_SLICE_X3Y131_B5Q;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C4 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C5 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO2;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C6 = BRAM_L_X6Y135_RAMB18_X0Y54_DO2;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A1 = BRAM_L_X6Y130_RAMB18_X0Y52_DO5;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A2 = CLBLM_R_X5Y132_SLICE_X6Y132_AQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A3 = CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A4 = CLBLM_L_X10Y135_SLICE_X12Y135_A5Q;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A6 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_AX = CLBLL_L_X4Y133_SLICE_X5Y133_CO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D1 = CLBLM_L_X10Y136_SLICE_X13Y136_AO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B1 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D3 = BRAM_L_X6Y135_RAMB18_X0Y54_DO0;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B2 = CLBLL_L_X4Y132_SLICE_X5Y132_BQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B4 = CLBLM_R_X3Y132_SLICE_X2Y132_DQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D6 = CLBLM_L_X16Y152_SLICE_X22Y152_AQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B5 = CLBLM_R_X3Y132_SLICE_X3Y132_CQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B6 = CLBLM_R_X3Y132_SLICE_X2Y132_BO5;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D5 = CLBLM_L_X10Y136_SLICE_X13Y136_BO5;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C1 = CLBLL_L_X2Y132_SLICE_X1Y132_AQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C2 = CLBLM_R_X5Y132_SLICE_X7Y132_B5Q;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A1 = BRAM_L_X6Y135_RAMB18_X0Y54_DO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A2 = CLBLM_L_X8Y137_SLICE_X10Y137_A5Q;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A3 = BRAM_R_X17Y135_RAMB18_X1Y54_DO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A4 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO5;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C6 = CLBLM_R_X3Y132_SLICE_X2Y132_AO5;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A5 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A6 = BRAM_L_X6Y135_RAMB18_X0Y54_DO5;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C3 = CLBLM_R_X3Y132_SLICE_X2Y132_CQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B1 = BRAM_R_X17Y135_RAMB18_X1Y54_DO4;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D1 = CLBLL_L_X4Y131_SLICE_X4Y131_CQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D2 = CLBLL_L_X4Y132_SLICE_X4Y132_AO5;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D3 = CLBLM_R_X5Y132_SLICE_X6Y132_B5Q;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D4 = CLBLL_L_X4Y132_SLICE_X4Y132_CQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D6 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B2 = BRAM_L_X6Y135_RAMB18_X0Y54_DO3;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B3 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO3;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B4 = BRAM_L_X6Y135_RAMB18_X0Y54_DO4;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B5 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO4;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B6 = CLBLM_L_X8Y136_SLICE_X10Y136_A5Q;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C1 = BRAM_L_X6Y135_RAMB18_X0Y54_DO7;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C2 = CLBLM_L_X8Y136_SLICE_X10Y136_A5Q;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C3 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO7;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C4 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C5 = CLBLM_L_X16Y154_SLICE_X22Y154_AQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C6 = CLBLM_L_X10Y136_SLICE_X12Y136_BO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D1 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D2 = CLBLM_L_X10Y136_SLICE_X13Y136_AO5;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D3 = CLBLM_L_X10Y136_SLICE_X13Y136_BO5;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D4 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO0;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D5 = CLBLM_R_X25Y149_SLICE_X37Y149_AQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D6 = CLBLM_R_X7Y129_SLICE_X8Y129_A5Q;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE = 1'b1;
  assign RIOI3_X105Y117_OLOGIC_X1Y118_D1 = CLBLM_L_X10Y131_SLICE_X12Y131_AQ;
  assign RIOI3_X105Y117_OLOGIC_X1Y118_T1 = 1'b1;
  assign RIOI3_X105Y117_OLOGIC_X1Y117_D1 = CLBLM_L_X12Y132_SLICE_X16Y132_AQ;
  assign RIOI3_X105Y117_OLOGIC_X1Y117_T1 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A1 = CLBLM_L_X8Y137_SLICE_X10Y137_A5Q;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A2 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A3 = CLBLL_L_X4Y133_SLICE_X4Y133_AQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A4 = CLBLL_L_X4Y132_SLICE_X4Y132_BQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A5 = BRAM_L_X6Y130_RAMB18_X0Y52_DO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A6 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_AX = CLBLL_L_X4Y133_SLICE_X4Y133_CO6;
  assign CLBLM_L_X16Y157_SLICE_X23Y157_A1 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B1 = CLBLM_R_X3Y133_SLICE_X3Y133_AO5;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B2 = CLBLL_L_X4Y133_SLICE_X4Y133_BQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B3 = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B5 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B6 = CLBLM_R_X3Y132_SLICE_X3Y132_BQ;
  assign CLBLM_L_X16Y157_SLICE_X23Y157_A2 = 1'b1;
  assign CLBLM_L_X16Y157_SLICE_X23Y157_A3 = 1'b1;
  assign CLBLM_L_X16Y157_SLICE_X23Y157_A4 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C1 = CLBLL_L_X4Y133_SLICE_X4Y133_BQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C2 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C3 = CLBLM_R_X3Y132_SLICE_X3Y132_BQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C4 = CLBLL_L_X4Y133_SLICE_X4Y133_A5Q;
  assign CLBLM_L_X16Y157_SLICE_X23Y157_B6 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C5 = CLBLM_R_X3Y133_SLICE_X3Y133_AO5;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_L_X16Y157_SLICE_X23Y157_B1 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y157_SLICE_X23Y157_B2 = 1'b1;
  assign CLBLM_L_X16Y157_SLICE_X23Y157_B3 = 1'b1;
  assign CLBLM_L_X16Y157_SLICE_X23Y157_B4 = 1'b1;
  assign CLBLM_L_X16Y157_SLICE_X23Y157_B5 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D1 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D2 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D3 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D4 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D5 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D6 = 1'b1;
  assign CLBLM_L_X16Y157_SLICE_X23Y157_C4 = 1'b1;
  assign CLBLM_L_X16Y157_SLICE_X23Y157_D1 = 1'b1;
  assign CLBLM_L_X16Y157_SLICE_X23Y157_D2 = 1'b1;
  assign CLBLM_L_X16Y157_SLICE_X23Y157_D3 = 1'b1;
  assign CLBLM_L_X16Y157_SLICE_X23Y157_D4 = 1'b1;
  assign CLBLM_L_X16Y157_SLICE_X23Y157_D5 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A1 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO4;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A2 = CLBLM_R_X7Y131_SLICE_X9Y131_A5Q;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A3 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO5;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A4 = BRAM_L_X6Y135_RAMB18_X0Y54_DO4;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A5 = BRAM_R_X17Y135_RAMB18_X1Y54_DO5;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A6 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO5;
  assign CLBLM_L_X16Y157_SLICE_X23Y157_D6 = 1'b1;
  assign CLBLM_L_X16Y157_SLICE_X22Y157_A1 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B1 = CLBLM_L_X16Y151_SLICE_X22Y151_CQ;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B2 = CLBLM_R_X7Y131_SLICE_X9Y131_A5Q;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B3 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B4 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B5 = CLBLM_L_X10Y137_SLICE_X13Y137_AO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B6 = 1'b1;
  assign CLBLM_L_X16Y157_SLICE_X22Y157_A2 = 1'b1;
  assign CLBLM_L_X16Y157_SLICE_X22Y157_A3 = 1'b1;
  assign CLBLM_L_X16Y157_SLICE_X22Y157_A4 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C1 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C2 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C3 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C4 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C5 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C6 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A1 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A2 = CLBLM_L_X8Y137_SLICE_X10Y137_B5Q;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A3 = CLBLL_L_X4Y133_SLICE_X5Y133_AQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A4 = BRAM_L_X6Y130_RAMB18_X0Y52_DO7;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A5 = LIOB33_X0Y87_IOB_X0Y87_I;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A6 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B1 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D1 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D2 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D3 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D4 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D5 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D6 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B2 = CLBLL_L_X4Y133_SLICE_X5Y133_BQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B3 = CLBLL_L_X4Y133_SLICE_X5Y133_AQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B5 = BRAM_L_X6Y130_RAMB18_X0Y52_DO7;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B6 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C1 = BRAM_L_X6Y130_RAMB18_X0Y52_DO7;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A1 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A2 = CLBLM_R_X7Y137_SLICE_X8Y137_A5Q;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A3 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO5;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C2 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C3 = CLBLL_L_X4Y133_SLICE_X5Y133_BQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C4 = CLBLL_L_X4Y133_SLICE_X5Y133_AO5;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C6 = CLBLL_L_X4Y132_SLICE_X5Y132_A5Q;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A4 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A5 = BRAM_R_X17Y135_RAMB18_X1Y54_DO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A6 = BRAM_L_X6Y135_RAMB18_X0Y54_DO5;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D1 = CLBLM_R_X5Y133_SLICE_X6Y133_BQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D2 = CLBLM_R_X3Y132_SLICE_X3Y132_AO5;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B1 = CLBLM_R_X7Y128_SLICE_X8Y128_A5Q;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B2 = BRAM_R_X17Y135_RAMB18_X1Y54_DO5;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B3 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO4;
  assign LIOI3_X0Y195_ILOGIC_X0Y196_D = LIOB33_X0Y195_IOB_X0Y196_I;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B4 = BRAM_R_X17Y135_RAMB18_X1Y54_DO4;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C1 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign LIOI3_X0Y195_ILOGIC_X0Y195_D = LIOB33_X0Y195_IOB_X0Y195_I;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B5 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO5;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B6 = BRAM_L_X6Y135_RAMB18_X0Y54_DO5;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C2 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C3 = CLBLM_R_X25Y151_SLICE_X36Y151_BQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C4 = CLBLM_L_X10Y137_SLICE_X12Y137_AO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C5 = CLBLM_R_X7Y137_SLICE_X8Y137_A5Q;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C6 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D1 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D2 = CLBLM_R_X7Y128_SLICE_X8Y128_A5Q;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D3 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D4 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D5 = CLBLM_R_X25Y149_SLICE_X36Y149_AQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D6 = CLBLM_L_X10Y137_SLICE_X12Y137_BO6;
  assign LIOI3_X0Y73_ILOGIC_X0Y74_D = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y73_D = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y158_D = LIOB33_X0Y157_IOB_X0Y158_I;
  assign LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y157_D = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A1 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A2 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A3 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A4 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A5 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A6 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_AX = CLBLM_R_X3Y134_SLICE_X3Y134_AO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B1 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B2 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B3 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B4 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B5 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B6 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C1 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C2 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C3 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C4 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C5 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C6 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D1 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D2 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D3 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D4 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D5 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D6 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A1 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A2 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A3 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A4 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A5 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A6 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B1 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B2 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B3 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B4 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B5 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B6 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A1 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A2 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A3 = CLBLL_L_X4Y133_SLICE_X5Y133_BQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A4 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO7;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A5 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A6 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C3 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C1 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C6 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C2 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B1 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B2 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B3 = CLBLL_L_X2Y132_SLICE_X1Y132_AQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B4 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B5 = BRAM_L_X6Y140_RAMB18_X0Y56_DO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B6 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C1 = CLBLL_L_X4Y145_SLICE_X4Y145_AQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C2 = CLBLL_L_X4Y135_SLICE_X5Y135_AO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C3 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO0;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C4 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D6 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C5 = CLBLM_R_X5Y130_SLICE_X6Y130_CQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C6 = CLBLM_R_X5Y134_SLICE_X6Y134_AO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D1 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D2 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D4 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D5 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A1 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A2 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A5 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A6 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D1 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D2 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D3 = CLBLM_R_X3Y147_SLICE_X2Y147_DQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D4 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D5 = CLBLM_R_X5Y134_SLICE_X6Y134_CO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D6 = CLBLL_L_X4Y132_SLICE_X5Y132_A5Q;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A4 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B1 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B2 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B3 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B4 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B5 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B6 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C1 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C2 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C3 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C4 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C5 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C6 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D1 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D2 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D3 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D4 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D5 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D6 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C4 = BRAM_L_X6Y125_RAMB18_X0Y50_DO22;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_A1 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO0;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_A2 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_A3 = BRAM_L_X6Y140_RAMB18_X0Y56_DO0;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_A4 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_A5 = CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_A6 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_B1 = BRAM_L_X6Y140_RAMB18_X0Y56_DO6;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_B2 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO5;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_B3 = CLBLL_L_X4Y133_SLICE_X4Y133_AQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_B4 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO5;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_B5 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO6;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_B6 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO6;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_C1 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO7;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_C2 = CLBLL_L_X4Y135_SLICE_X5Y135_CO6;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_C3 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_C4 = CLBLM_R_X5Y131_SLICE_X7Y131_CQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_C5 = CLBLM_R_X3Y155_SLICE_X3Y155_CQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_C6 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO7;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_D1 = CLBLL_L_X4Y133_SLICE_X4Y133_AQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_D2 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_D3 = CLBLL_L_X2Y157_SLICE_X1Y157_AQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_D4 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_D5 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_D6 = CLBLL_L_X4Y135_SLICE_X4Y135_BO6;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_A1 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO0;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_A2 = BRAM_L_X6Y140_RAMB18_X0Y56_DO16;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_A3 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_A4 = CLBLM_R_X5Y127_SLICE_X6Y127_CQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_A5 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_A6 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_B1 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_B2 = CLBLL_L_X4Y133_SLICE_X4Y133_BQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_B3 = BRAM_L_X6Y140_RAMB18_X0Y56_DO5;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_B4 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_B5 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_B6 = 1'b1;
  assign RIOI3_X105Y121_OLOGIC_X1Y122_D1 = CLBLM_L_X10Y133_SLICE_X13Y133_CQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_C1 = CLBLM_R_X5Y131_SLICE_X7Y131_CQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_C2 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO3;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_C3 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO4;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_C4 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO3;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_C5 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO4;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_C6 = BRAM_L_X6Y140_RAMB18_X0Y56_DO4;
  assign RIOI3_X105Y121_OLOGIC_X1Y122_T1 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_D1 = CLBLL_L_X4Y135_SLICE_X5Y135_AO6;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_D2 = CLBLM_R_X5Y130_SLICE_X7Y130_CQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_D3 = CLBLM_R_X3Y141_SLICE_X2Y141_CQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_D4 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_D5 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO0;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_D6 = CLBLM_R_X5Y134_SLICE_X6Y134_BO6;
  assign RIOI3_X105Y121_OLOGIC_X1Y121_D1 = CLBLM_R_X11Y133_SLICE_X14Y133_BQ;
  assign RIOI3_X105Y121_OLOGIC_X1Y121_T1 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X82Y96_A1 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X82Y96_A2 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X82Y96_A3 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X82Y96_A4 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X82Y96_A5 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X82Y96_A6 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X82Y96_AX = CLBLM_L_X8Y130_SLICE_X11Y130_AO5;
  assign CLBLL_L_X54Y96_SLICE_X82Y96_B1 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X82Y96_B2 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X82Y96_B3 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X82Y96_B4 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X82Y96_B5 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X82Y96_B6 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X82Y96_C1 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X82Y96_C2 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X82Y96_C3 = 1'b1;
  assign CLBLL_L_X54Y123_SLICE_X83Y123_C1 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X82Y96_C4 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X82Y96_C5 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X82Y96_C6 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X82Y96_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X0Y20_O;
  assign CLBLL_L_X54Y96_SLICE_X82Y96_D1 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X82Y96_D2 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X82Y96_D3 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X82Y96_D4 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X82Y96_D5 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X82Y96_D6 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X83Y96_A1 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X83Y96_A2 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X83Y96_A3 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X83Y96_A4 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X83Y96_A5 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X83Y96_A6 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X83Y96_B1 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X83Y96_B2 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X83Y96_B3 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X83Y96_B4 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X83Y96_B5 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X83Y96_B6 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X83Y96_C1 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X83Y96_C2 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X83Y96_C3 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X83Y96_C4 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X83Y96_C5 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X83Y96_C6 = 1'b1;
  assign LIOI3_X0Y197_ILOGIC_X0Y198_D = LIOB33_X0Y197_IOB_X0Y198_I;
  assign LIOI3_X0Y197_ILOGIC_X0Y197_D = LIOB33_X0Y197_IOB_X0Y197_I;
  assign CLBLL_L_X54Y96_SLICE_X83Y96_D1 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X83Y96_D2 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X83Y96_D3 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X83Y96_D4 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X83Y96_D5 = 1'b1;
  assign CLBLL_L_X54Y96_SLICE_X83Y96_D6 = 1'b1;
  assign LIOI3_X0Y75_ILOGIC_X0Y76_D = LIOB33_X0Y75_IOB_X0Y76_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y75_D = LIOB33_X0Y75_IOB_X0Y75_I;
  assign LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y170_D = LIOB33_X0Y169_IOB_X0Y170_I;
  assign LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y169_D = LIOB33_X0Y169_IOB_X0Y169_I;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_A1 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO6;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_A2 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO6;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_A3 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO5;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_A4 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO6;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_A5 = CLBLL_L_X2Y132_SLICE_X1Y132_AQ;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_A6 = BRAM_L_X6Y140_RAMB18_X0Y56_DO5;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_B1 = BRAM_L_X6Y140_RAMB18_X0Y56_DO3;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_B2 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO3;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_B3 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO2;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_B4 = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_B5 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO3;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_B6 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO2;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_C1 = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_C2 = CLBLL_L_X4Y136_SLICE_X4Y136_BO6;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_C3 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO7;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_C4 = CLBLM_R_X3Y153_SLICE_X2Y153_DQ;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_C5 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO7;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_C6 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_D1 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_D2 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_D3 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_D4 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_D5 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_D6 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_A1 = CLBLM_R_X5Y129_SLICE_X6Y129_AQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_A2 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO2;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_A3 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO3;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_A4 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO3;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_A5 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO3;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_A6 = BRAM_L_X6Y140_RAMB18_X0Y56_DO2;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_B1 = BRAM_L_X6Y140_RAMB18_X0Y56_DO2;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_B2 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO2;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_B3 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO1;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_B4 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO1;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_B5 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO2;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_B6 = CLBLL_L_X4Y129_SLICE_X5Y129_CQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_C1 = CLBLM_R_X5Y136_SLICE_X6Y136_CO6;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_C2 = CLBLM_R_X3Y141_SLICE_X2Y141_BQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_C3 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_C4 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_C5 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_C6 = CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_D1 = CLBLM_R_X3Y153_SLICE_X2Y153_CQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_D2 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_D3 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_D4 = CLBLL_L_X4Y129_SLICE_X5Y129_CQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_D5 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_D6 = CLBLL_L_X4Y136_SLICE_X5Y136_BO6;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_A1 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO1;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_A2 = BRAM_L_X6Y140_RAMB18_X0Y56_DO0;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_A3 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO0;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_A4 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO1;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_A5 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO1;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_A6 = CLBLL_L_X4Y132_SLICE_X4Y132_CQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_B1 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO1;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_B2 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO2;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_B3 = CLBLL_L_X4Y131_SLICE_X4Y131_DQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_B4 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO1;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_B5 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO2;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_B6 = BRAM_L_X6Y140_RAMB18_X0Y56_DO2;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_C1 = CLBLL_L_X4Y135_SLICE_X4Y135_AO6;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_C2 = CLBLM_R_X3Y155_SLICE_X3Y155_BQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_C3 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_C4 = CLBLM_R_X5Y131_SLICE_X6Y131_CQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_C5 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO0;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_C6 = CLBLM_R_X3Y137_SLICE_X3Y137_AO6;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_D1 = BRAM_L_X6Y140_RAMB18_X0Y56_DO0;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_D2 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO0;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_D3 = BRAM_L_X6Y140_RAMB18_X0Y56_DO1;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_D4 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO1;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_D5 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO1;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_D6 = CLBLM_R_X5Y125_SLICE_X7Y125_CQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_A1 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO7;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_A2 = 1'b1;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_A3 = CLBLL_L_X4Y128_SLICE_X5Y128_BQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_A4 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO7;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_A5 = 1'b1;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_A6 = 1'b1;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_B1 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO3;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_B2 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO3;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_B3 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO4;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_B4 = BRAM_L_X6Y140_RAMB18_X0Y56_DO4;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_B5 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO4;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_B6 = CLBLL_L_X4Y131_SLICE_X5Y131_BQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_C1 = CLBLL_L_X4Y155_SLICE_X4Y155_AQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_C2 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO7;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_C3 = CLBLL_L_X4Y131_SLICE_X5Y131_BQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_C4 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO7;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_C5 = CLBLL_L_X4Y137_SLICE_X5Y137_BO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_C6 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_D1 = CLBLL_L_X4Y137_SLICE_X5Y137_AO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_D2 = CLBLM_R_X5Y129_SLICE_X7Y129_BQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_D3 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO0;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_D4 = CLBLM_R_X3Y153_SLICE_X2Y153_AQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_D5 = CLBLL_L_X4Y135_SLICE_X4Y135_AO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_D6 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign RIOI3_X105Y123_OLOGIC_X1Y124_D1 = CLBLM_R_X7Y130_SLICE_X9Y130_BQ;
  assign RIOI3_X105Y123_OLOGIC_X1Y124_T1 = 1'b1;
  assign RIOI3_X105Y123_OLOGIC_X1Y123_D1 = CLBLM_L_X12Y132_SLICE_X16Y132_BQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A2 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A3 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A4 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A5 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A6 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_AX = CLBLM_R_X7Y125_SLICE_X8Y125_DO6;
  assign RIOI3_X105Y123_OLOGIC_X1Y123_T1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B2 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B3 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B4 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B5 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B6 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_BX = CLBLM_R_X5Y125_SLICE_X7Y125_DO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C2 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C3 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C4 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C5 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C6 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D2 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D3 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D4 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D5 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D6 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A2 = CLBLM_R_X5Y125_SLICE_X7Y125_BQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A3 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A4 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO2;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A5 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A6 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B1 = CLBLM_R_X7Y125_SLICE_X8Y125_B5Q;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B2 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B3 = BRAM_L_X6Y125_RAMB18_X0Y50_DO1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B4 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B5 = LIOB33_X0Y97_IOB_X0Y97_I;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B6 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C1 = CLBLM_R_X7Y125_SLICE_X8Y125_C5Q;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C2 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C3 = LIOB33_X0Y97_IOB_X0Y98_I;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C4 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO2;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C5 = BRAM_L_X6Y125_RAMB18_X0Y50_DO2;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A1 = BRAM_L_X6Y140_RAMB18_X0Y56_DO1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A2 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A3 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A4 = CLBLL_L_X4Y130_SLICE_X4Y130_BQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A5 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO0;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A6 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO0;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C6 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B1 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO7;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D1 = BRAM_L_X6Y125_RAMB18_X0Y50_DO1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D2 = CLBLM_R_X5Y125_SLICE_X7Y125_CQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D3 = CLBLM_R_X7Y125_SLICE_X9Y125_AQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D4 = CLBLM_R_X5Y125_SLICE_X7Y125_AO5;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D5 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D6 = LIOB33_X0Y1_IOB_X0Y1_I;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B2 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO7;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B3 = CLBLL_L_X2Y155_SLICE_X0Y155_AQ;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B4 = CLBLL_L_X4Y130_SLICE_X4Y130_BQ;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B5 = CLBLL_L_X4Y138_SLICE_X4Y138_AO6;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B6 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C1 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO2;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C2 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO3;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C3 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO3;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C5 = BRAM_L_X6Y140_RAMB18_X0Y56_DO3;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C6 = CLBLM_R_X5Y126_SLICE_X6Y126_BQ;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C4 = BRAM_L_X6Y140_RAMB18_X0Y56_DO2;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D1 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D2 = BRAM_L_X6Y140_RAMB18_X0Y56_DO2;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D3 = CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D4 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO2;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D5 = BRAM_L_X6Y140_RAMB18_X0Y56_DO1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D6 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO2;
  assign LIOI3_X0Y201_ILOGIC_X0Y202_D = LIOB33_X0Y201_IOB_X0Y202_I;
  assign LIOI3_X0Y201_ILOGIC_X0Y201_D = LIOB33_X0Y201_IOB_X0Y201_I;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A1 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO5;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A2 = CLBLL_L_X4Y133_SLICE_X4Y133_BQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A3 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO4;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A4 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO5;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A5 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO5;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A6 = BRAM_L_X6Y140_RAMB18_X0Y56_DO4;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B1 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO4;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B2 = BRAM_L_X6Y140_RAMB18_X0Y56_DO3;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B3 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO4;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B4 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO3;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B5 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO4;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B6 = CLBLM_R_X3Y133_SLICE_X3Y133_BQ;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_D = LIOB33_X0Y77_IOB_X0Y78_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y77_D = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C1 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO2;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C2 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO2;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C3 = BRAM_L_X6Y140_RAMB18_X0Y56_DO1;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C4 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO1;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C5 = CLBLL_L_X4Y130_SLICE_X5Y130_AQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C6 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO2;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D1 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO5;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D2 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO4;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D3 = CLBLM_R_X5Y127_SLICE_X7Y127_BQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D4 = BRAM_L_X6Y140_RAMB18_X0Y56_DO4;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D5 = BRAM_L_X6Y140_RAMB18_X0Y56_DO5;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D6 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO5;
  assign LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y182_D = LIOB33_X0Y181_IOB_X0Y182_I;
  assign LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y181_D = LIOB33_X0Y181_IOB_X0Y181_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A1 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A2 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A3 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A4 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A5 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A6 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_AX = CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B1 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B2 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B3 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B4 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B5 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B6 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C1 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C2 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C3 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C4 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C5 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C6 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D1 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D2 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D3 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D4 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D5 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D6 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A1 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A2 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A3 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A4 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A5 = CLBLM_R_X7Y125_SLICE_X9Y125_AQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A6 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B1 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B2 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO2;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B3 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B4 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B5 = CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B6 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C1 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C2 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C3 = CLBLM_R_X5Y126_SLICE_X7Y126_B5Q;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C4 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C5 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C6 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO3;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_A1 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_A2 = CLBLL_L_X4Y136_SLICE_X5Y136_AO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_A3 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO7;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_A4 = CLBLL_L_X2Y157_SLICE_X1Y157_BQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_A5 = BRAM_L_X6Y140_RAMB18_X0Y56_DO7;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_A6 = CLBLM_R_X5Y129_SLICE_X6Y129_AQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_B1 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D1 = LIOB33_SING_X0Y99_IOB_X0Y99_I;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D2 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D3 = BRAM_L_X6Y125_RAMB18_X0Y50_DO3;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D4 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO3;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D5 = CLBLM_R_X7Y126_SLICE_X8Y126_D5Q;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D6 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_B4 = CLBLL_L_X4Y156_SLICE_X4Y156_AQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_B5 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO7;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_B6 = BRAM_L_X6Y140_RAMB18_X0Y56_DO7;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_C1 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO7;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_C2 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO0;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_C3 = BRAM_L_X6Y140_RAMB18_X0Y56_DO7;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_C4 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO0;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_C5 = BRAM_L_X6Y140_RAMB18_X0Y56_DO0;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_C6 = CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_D1 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_D2 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_D3 = CLBLM_R_X5Y127_SLICE_X6Y127_CQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_D4 = CLBLL_L_X4Y139_SLICE_X5Y139_BO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_D5 = CLBLM_R_X3Y141_SLICE_X2Y141_AQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_D6 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_A1 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO0;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_A2 = CLBLM_R_X5Y130_SLICE_X7Y130_BQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_A3 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO0;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_A4 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO7;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_A5 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO0;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_A6 = BRAM_L_X6Y140_RAMB18_X0Y56_DO23;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_B1 = CLBLM_R_X5Y127_SLICE_X6Y127_CQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_B2 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO7;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_B3 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO0;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_B4 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO0;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_B5 = BRAM_L_X6Y140_RAMB18_X0Y56_DO16;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_B6 = BRAM_L_X6Y140_RAMB18_X0Y56_DO23;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_C1 = CLBLL_L_X2Y158_SLICE_X0Y158_AQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_C2 = CLBLL_L_X4Y138_SLICE_X5Y138_CO6;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_C3 = CLBLL_L_X4Y130_SLICE_X5Y130_AQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_C4 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_C5 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_C6 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_D1 = CLBLM_R_X5Y127_SLICE_X7Y127_BQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_D2 = CLBLL_L_X4Y138_SLICE_X5Y138_DO6;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_D3 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_D4 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_D5 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_D6 = CLBLL_L_X2Y152_SLICE_X0Y152_AQ;
  assign CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_CE = 1'b1;
  assign CLK_HROW_TOP_R_X139Y182_BUFHCE_X1Y44_CE = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A1 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A2 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A3 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A4 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A5 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A6 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B1 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B2 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B3 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B4 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B5 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B6 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C1 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C2 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C3 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C4 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C5 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C6 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D1 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D2 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D3 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D4 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D5 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D6 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A1 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO0;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A2 = CLBLM_R_X7Y127_SLICE_X8Y127_A5Q;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A3 = BRAM_L_X6Y125_RAMB18_X0Y50_DO0;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A5 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A6 = 1'b1;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_D = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B1 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B2 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B3 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B4 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B5 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A1 = CLBLL_L_X4Y138_SLICE_X4Y138_DO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A2 = CLBLM_R_X3Y151_SLICE_X2Y151_DQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A3 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A4 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A5 = CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A6 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C2 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B6 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C5 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B2 = CLBLL_L_X4Y139_SLICE_X4Y139_CO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B3 = CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B4 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B5 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B6 = CLBLM_R_X3Y151_SLICE_X2Y151_BQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C2 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C3 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C4 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C5 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C6 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D6 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D1 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D2 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D3 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D4 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D5 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D2 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D3 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D4 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D5 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D6 = 1'b1;
  assign RIOI3_X105Y125_OLOGIC_X1Y126_T1 = 1'b1;
  assign RIOI3_X105Y125_OLOGIC_X1Y125_D1 = CLBLM_R_X5Y132_SLICE_X7Y132_AQ;
  assign RIOI3_X105Y125_OLOGIC_X1Y125_T1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A2 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A3 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A4 = CLBLM_R_X3Y149_SLICE_X3Y149_AQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A5 = CLBLL_L_X4Y139_SLICE_X5Y139_AO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A6 = CLBLM_R_X5Y130_SLICE_X7Y130_BQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B2 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B3 = CLBLL_L_X4Y138_SLICE_X5Y138_AO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B4 = CLBLL_L_X4Y133_SLICE_X4Y133_BQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B5 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B6 = CLBLL_L_X2Y157_SLICE_X0Y157_BQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C2 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C3 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C4 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C5 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C6 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D2 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D3 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D4 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D5 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D6 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_A1 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_A2 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_A3 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_A4 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_A5 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_A6 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_AX = CLBLM_R_X7Y130_SLICE_X8Y130_AO5;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_B1 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_B2 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_B3 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_B4 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_B5 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_B6 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_C1 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_C2 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_C3 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_C4 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_C5 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_C6 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_D1 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_D2 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_D3 = 1'b1;
  assign LIOI3_X0Y203_ILOGIC_X0Y204_D = LIOB33_X0Y203_IOB_X0Y204_I;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_D4 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_D5 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_D6 = 1'b1;
  assign LIOI3_X0Y203_ILOGIC_X0Y203_D = LIOB33_X0Y203_IOB_X0Y203_I;
  assign CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLK_HROW_TOP_R_X139Y182_BUFHCE_X1Y44_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_A1 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_A2 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_A3 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_A4 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_A5 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_A6 = 1'b1;
  assign LIOI3_X0Y79_ILOGIC_X0Y80_D = LIOB33_X0Y79_IOB_X0Y80_I;
  assign LIOI3_X0Y79_ILOGIC_X0Y79_D = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_B1 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_B2 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_B3 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_B4 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_B5 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_B6 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_C1 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_C2 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_C3 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_C4 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_C5 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_C6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y194_D = LIOB33_X0Y193_IOB_X0Y194_I;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_D1 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_D2 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_D3 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_D4 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_D5 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_D6 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A1 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A2 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A3 = CLBLM_R_X5Y128_SLICE_X7Y128_AQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A4 = BRAM_L_X6Y135_RAMB18_X0Y54_DO16;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A5 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A6 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B1 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B2 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B3 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B4 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B5 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B6 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C1 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C2 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C3 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C4 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C5 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C6 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D1 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D2 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D3 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D4 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D5 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D6 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A1 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A2 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A3 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO5;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A4 = BRAM_L_X6Y125_RAMB18_X0Y50_DO5;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A5 = CLBLM_R_X7Y128_SLICE_X8Y128_A5Q;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A6 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B1 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B2 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B3 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO4;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B4 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B5 = CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B6 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C1 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C2 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C3 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C4 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C5 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C6 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D1 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D2 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D3 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D4 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D5 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D6 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A1 = LIOB33_X0Y119_IOB_X0Y119_I;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A2 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A3 = CLBLM_R_X7Y129_SLICE_X9Y129_A5Q;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A4 = BRAM_L_X6Y125_RAMB18_X0Y50_DO4;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A5 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO4;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A6 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B3 = CLBLM_R_X3Y132_SLICE_X2Y132_AQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B4 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B1 = CLBLM_R_X7Y129_SLICE_X9Y129_B5Q;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B2 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B3 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B4 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B5 = BRAM_L_X6Y125_RAMB18_X0Y50_DO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B6 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C2 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C3 = CLBLM_R_X5Y127_SLICE_X7Y127_B5Q;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C4 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C5 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C6 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO5;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D2 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D3 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D4 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D5 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D6 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C1 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO7;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A1 = BRAM_L_X6Y135_RAMB18_X0Y54_DO0;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A2 = BRAM_L_X6Y125_RAMB18_X0Y50_DO16;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A3 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A5 = CLBLM_R_X7Y129_SLICE_X8Y129_A5Q;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A6 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C2 = BRAM_L_X6Y135_RAMB18_X0Y54_DO7;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C3 = BRAM_R_X17Y135_RAMB18_X1Y54_DO7;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B1 = BRAM_L_X6Y125_RAMB18_X0Y50_DO18;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B2 = CLBLM_R_X7Y129_SLICE_X8Y129_B5Q;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B3 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B5 = BRAM_L_X6Y135_RAMB18_X0Y54_DO2;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B6 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C4 = BRAM_L_X6Y135_RAMB18_X0Y54_DO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C1 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C2 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C3 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C4 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C5 = CLBLM_R_X5Y129_SLICE_X7Y129_B5Q;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C6 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C6 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D1 = CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D2 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D3 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D4 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D5 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D6 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO2;
  assign RIOI3_X105Y127_OLOGIC_X1Y128_D1 = CLBLM_L_X8Y134_SLICE_X10Y134_AQ;
  assign RIOI3_X105Y127_OLOGIC_X1Y128_T1 = 1'b1;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_D1 = CLBLM_R_X5Y133_SLICE_X7Y133_AQ;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_T1 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_ADDRBWRADDR12 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_ADDRBWRADDR13 = 1'b0;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_DIADI0 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_DIADI1 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_DIADI2 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_DIADI4 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A1 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_DIADI5 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A2 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A3 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A4 = CLBLM_R_X5Y129_SLICE_X6Y129_A5Q;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A5 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO3;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_DIADI6 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A6 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B1 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B2 = BRAM_L_X6Y140_RAMB18_X0Y56_DO16;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B3 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B4 = CLBLM_R_X5Y130_SLICE_X7Y130_BQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B5 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B6 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_DIADI8 = 1'b0;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C1 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_DIADI9 = 1'b0;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C2 = BRAM_L_X6Y140_RAMB18_X0Y56_DO18;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C3 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C4 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C5 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_DIADI10 = 1'b0;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C6 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D1 = CLBLL_L_X4Y129_SLICE_X5Y129_AQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D2 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D3 = BRAM_L_X6Y135_RAMB18_X0Y54_DO18;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D4 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D5 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D6 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_DIADI13 = 1'b0;
  assign LIOI3_X0Y205_ILOGIC_X0Y206_D = LIOB33_X0Y205_IOB_X0Y206_I;
  assign LIOI3_X0Y205_ILOGIC_X0Y205_D = LIOB33_X0Y205_IOB_X0Y205_I;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A1 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A2 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A3 = CLBLL_L_X4Y128_SLICE_X5Y128_AQ;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_DIADI15 = 1'b0;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A4 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO7;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A5 = BRAM_L_X6Y135_RAMB18_X0Y54_DO23;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A6 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_DIBDI0 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_AX = CLBLL_L_X4Y129_SLICE_X5Y129_DO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B1 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO0;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B2 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_DIBDI1 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B3 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B4 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B5 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B6 = CLBLM_R_X5Y130_SLICE_X7Y130_CQ;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_DIBDI2 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_BX = CLBLL_L_X4Y130_SLICE_X5Y130_BO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C1 = CLBLM_R_X5Y125_SLICE_X7Y125_BQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C2 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO2;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_DIBDI3 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C3 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C4 = BRAM_R_X17Y135_RAMB18_X1Y54_DO17;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C5 = BRAM_L_X6Y135_RAMB18_X0Y54_DO18;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C6 = BRAM_R_X17Y135_RAMB18_X1Y54_DO18;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_DIBDI4 = 1'b1;
  assign LIOI3_X0Y83_ILOGIC_X0Y84_D = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y83_ILOGIC_X0Y83_D = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D1 = CLBLM_R_X5Y125_SLICE_X7Y125_BQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D2 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D3 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D4 = CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D5 = CLBLL_L_X4Y156_SLICE_X4Y156_CQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D6 = 1'b1;
  assign BRAM_L_X6Y135_RAMB18_X0Y55_DIBDI7 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y207_ILOGIC_X0Y208_D = LIOB33_X0Y207_IOB_X0Y208_I;
  assign LIOI3_TBYTESRC_X0Y207_ILOGIC_X0Y207_D = LIOB33_X0Y207_IOB_X0Y207_I;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A1 = BRAM_L_X6Y135_RAMB18_X0Y54_DO5;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A2 = BRAM_L_X6Y125_RAMB18_X0Y50_DO21;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A3 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A5 = CLBLM_R_X7Y131_SLICE_X9Y131_A5Q;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A6 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B1 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B2 = CLBLM_R_X5Y130_SLICE_X7Y130_A5Q;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B3 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B4 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B5 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO4;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B6 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C1 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C2 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO5;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C3 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C4 = CLBLL_L_X4Y130_SLICE_X5Y130_A5Q;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C5 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C6 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D1 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D2 = CLBLM_R_X5Y130_SLICE_X6Y130_B5Q;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D3 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D4 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D5 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D6 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A1 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A2 = CLBLM_R_X7Y130_SLICE_X8Y130_AO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A3 = CLBLM_R_X5Y128_SLICE_X7Y128_AQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A4 = CLBLM_R_X3Y155_SLICE_X2Y155_AQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A5 = CLBLM_L_X8Y130_SLICE_X11Y130_AO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A6 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO0;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B1 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B2 = CLBLL_L_X4Y129_SLICE_X4Y129_AQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B3 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B4 = BRAM_L_X6Y135_RAMB18_X0Y54_DO16;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B5 = BRAM_R_X17Y135_RAMB18_X1Y54_DO17;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B6 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO0;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C1 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO7;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C2 = BRAM_R_X17Y135_RAMB18_X1Y54_DO23;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C3 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C4 = CLBLM_R_X5Y126_SLICE_X6Y126_AQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C5 = CLBLL_L_X4Y156_SLICE_X4Y156_DQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C6 = CLBLM_L_X8Y131_SLICE_X10Y131_CO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D1 = CLBLL_L_X4Y156_SLICE_X4Y156_BQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D2 = BRAM_R_X17Y135_RAMB18_X1Y54_DO23;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D3 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D4 = CLBLM_L_X8Y131_SLICE_X10Y131_DO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D5 = CLBLM_R_X5Y125_SLICE_X7Y125_AQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D6 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO7;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_A1 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_A2 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_A3 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_A4 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_A5 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_A6 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_AX = CLBLM_L_X8Y133_SLICE_X11Y133_AO5;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_B1 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_B2 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_B3 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_B4 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_B5 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_B6 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_C1 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_C2 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_C3 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_C4 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_C5 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_C6 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_D1 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_D2 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_D3 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_D4 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_D5 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_D6 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_A1 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_A2 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_A3 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_A4 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_A5 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_A6 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_B1 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_B2 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_B3 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_B4 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_B5 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_B6 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_C1 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_C2 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_C3 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_C4 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_C5 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_C6 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_D1 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_D2 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_D3 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_D4 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_D5 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_D6 = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_D1 = CLBLM_L_X8Y132_SLICE_X11Y132_BQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A1 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A2 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A3 = CLBLL_L_X4Y133_SLICE_X4Y133_AQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A4 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A5 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A6 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B1 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO2;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B2 = BRAM_R_X17Y135_RAMB18_X1Y54_DO18;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B3 = CLBLL_L_X4Y129_SLICE_X5Y129_AQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B4 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO2;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B5 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B6 = BRAM_L_X6Y135_RAMB18_X0Y54_DO17;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_T1 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C1 = BRAM_R_X17Y135_RAMB18_X1Y54_DO20;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C2 = BRAM_L_X6Y135_RAMB18_X0Y54_DO20;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C3 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO3;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C4 = BRAM_R_X17Y135_RAMB18_X1Y54_DO19;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C5 = CLBLM_R_X5Y126_SLICE_X7Y126_AQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C6 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO4;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_D1 = CLBLM_R_X7Y133_SLICE_X9Y133_AQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D1 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO7;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D2 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO0;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D3 = CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D4 = BRAM_L_X6Y135_RAMB18_X0Y54_DO16;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D5 = BRAM_R_X17Y135_RAMB18_X1Y54_DO23;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A1 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A2 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A3 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A4 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A5 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A6 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D6 = BRAM_R_X17Y135_RAMB18_X1Y54_DO16;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_AX = LIOB33_X0Y165_IOB_X0Y166_I;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A1 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B1 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A4 = BRAM_L_X6Y125_RAMB18_X0Y50_DO20;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A5 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A6 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B2 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B3 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B4 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B5 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B1 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B2 = CLBLL_L_X4Y129_SLICE_X4Y129_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B3 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO7;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B4 = CLBLM_R_X3Y158_SLICE_X3Y158_CQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B5 = CLBLM_R_X7Y131_SLICE_X8Y131_BO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B6 = BRAM_L_X6Y135_RAMB18_X0Y54_DO23;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_BX = LIOB33_X0Y167_IOB_X0Y167_I;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C1 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C2 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_BX = CLBLM_R_X5Y132_SLICE_X6Y132_DO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C3 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C4 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C5 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C6 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C5 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C1 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO7;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C2 = CLBLM_R_X7Y132_SLICE_X9Y132_CO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C3 = CLBLM_R_X5Y126_SLICE_X7Y126_AQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D1 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D2 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D3 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D4 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D5 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D6 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_CX = CLBLM_R_X5Y132_SLICE_X6Y132_CO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D1 = CLBLM_R_X3Y158_SLICE_X3Y158_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D2 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D3 = CLBLM_R_X7Y132_SLICE_X9Y132_DO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D4 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D5 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D6 = CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A1 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A2 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A3 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A4 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A5 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A6 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B1 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B2 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B3 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B4 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B5 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B6 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C1 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C2 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C3 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C4 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C5 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C6 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D1 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D2 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D3 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D4 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D5 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D6 = 1'b1;
  assign LIOI3_X0Y209_ILOGIC_X0Y210_D = LIOB33_X0Y209_IOB_X0Y210_I;
  assign LIOI3_X0Y209_ILOGIC_X0Y209_D = LIOB33_X0Y209_IOB_X0Y209_I;
  assign LIOI3_X0Y85_ILOGIC_X0Y86_D = LIOB33_X0Y85_IOB_X0Y86_I;
  assign LIOI3_X0Y85_ILOGIC_X0Y85_D = LIOB33_X0Y85_IOB_X0Y85_I;
  assign LIOI3_TBYTESRC_X0Y219_ILOGIC_X0Y220_D = LIOB33_X0Y219_IOB_X0Y220_I;
  assign LIOI3_TBYTESRC_X0Y219_ILOGIC_X0Y219_D = LIOB33_X0Y219_IOB_X0Y219_I;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A1 = CLBLL_L_X4Y133_SLICE_X4Y133_A5Q;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A2 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A3 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A4 = BRAM_L_X6Y140_RAMB18_X0Y56_DO21;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A5 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A6 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B1 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B2 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B3 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B4 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B5 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B6 = CLBLM_R_X5Y125_SLICE_X7Y125_CQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C1 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO2;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C2 = BRAM_R_X17Y135_RAMB18_X1Y54_DO19;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C3 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO3;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C4 = BRAM_L_X6Y135_RAMB18_X0Y54_DO18;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C5 = CLBLM_R_X5Y128_SLICE_X6Y128_AQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C6 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO3;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A1 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A2 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A3 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D4 = BRAM_R_X17Y135_RAMB18_X1Y54_DO20;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D5 = BRAM_L_X6Y135_RAMB18_X0Y54_DO21;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D6 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A4 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A5 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A6 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D1 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO4;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D2 = BRAM_R_X17Y135_RAMB18_X1Y54_DO21;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_AX = LIOB33_X0Y169_IOB_X0Y169_I;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B1 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B2 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B3 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B4 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B5 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B6 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A1 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO7;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A2 = CLBLM_R_X7Y132_SLICE_X8Y132_BQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A3 = CLBLL_L_X4Y146_SLICE_X4Y146_AQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C1 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C2 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C3 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C4 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C5 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B4 = CLBLM_R_X7Y132_SLICE_X8Y132_BQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B5 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO2;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B6 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO3;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C6 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B2 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO2;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C1 = BRAM_L_X6Y135_RAMB18_X0Y54_DO23;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D1 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D2 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D3 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D5 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D6 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D4 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C2 = CLBLM_R_X7Y133_SLICE_X9Y133_CO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C3 = CLBLM_R_X5Y128_SLICE_X6Y128_AQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C4 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C5 = CLBLM_R_X3Y155_SLICE_X2Y155_BQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C6 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO7;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D1 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D2 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D3 = CLBLM_R_X7Y133_SLICE_X9Y133_DO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D4 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D5 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D6 = CLBLL_L_X2Y157_SLICE_X0Y157_DQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A1 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A2 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A3 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A4 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A5 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A6 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B1 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B2 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B3 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B4 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B5 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B6 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C1 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C2 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C3 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C4 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C5 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C6 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D1 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D2 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D3 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D4 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D5 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y193_D = LIOB33_X0Y193_IOB_X0Y193_I;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A2 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A3 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A4 = BRAM_R_X17Y135_RAMB18_X1Y54_DO22;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A5 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A6 = CLBLM_R_X3Y132_SLICE_X2Y132_CQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B2 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B3 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B4 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B5 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B6 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A1 = BRAM_L_X6Y130_RAMB18_X0Y52_DO2;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A2 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO2;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A3 = LIOB33_X0Y133_IOB_X0Y134_I;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A5 = CLBLM_R_X7Y134_SLICE_X9Y134_A5Q;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A6 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B1 = CLBLM_R_X7Y134_SLICE_X9Y134_B5Q;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B2 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B3 = BRAM_L_X6Y130_RAMB18_X0Y52_DO3;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B4 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO3;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B5 = LIOB33_X0Y135_IOB_X0Y135_I;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B6 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C1 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C1 = CLBLL_L_X4Y131_SLICE_X5Y131_AQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C2 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO3;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C3 = BRAM_L_X6Y135_RAMB18_X0Y54_DO19;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C4 = BRAM_R_X17Y135_RAMB18_X1Y54_DO20;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C2 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C5 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO4;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C6 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO4;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C3 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C4 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D1 = BRAM_L_X6Y135_RAMB18_X0Y54_DO3;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D2 = CLBLM_R_X7Y126_SLICE_X8Y126_D5Q;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D3 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO2;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D4 = BRAM_R_X17Y135_RAMB18_X1Y54_DO2;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D5 = BRAM_R_X17Y135_RAMB18_X1Y54_DO3;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D6 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO3;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C6 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A1 = BRAM_L_X6Y140_RAMB18_X0Y56_DO21;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A2 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO5;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A3 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO4;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A4 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO5;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A5 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO4;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A6 = CLBLM_R_X7Y132_SLICE_X8Y132_CQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B1 = BRAM_L_X6Y135_RAMB18_X0Y54_DO20;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B2 = BRAM_R_X17Y135_RAMB18_X1Y54_DO21;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B3 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO5;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B4 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO5;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B5 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO4;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B6 = CLBLM_R_X3Y130_SLICE_X3Y130_AQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C1 = BRAM_R_X17Y135_RAMB18_X1Y54_DO7;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C2 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO7;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C3 = CLBLM_R_X7Y134_SLICE_X9Y134_DO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C4 = CLBLM_R_X7Y126_SLICE_X8Y126_D5Q;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C5 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C6 = CLBLM_R_X3Y157_SLICE_X2Y157_DQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D1 = CLBLM_R_X7Y125_SLICE_X8Y125_C5Q;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D2 = CLBLM_L_X8Y134_SLICE_X10Y134_DO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D3 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D4 = CLBLM_R_X3Y157_SLICE_X2Y157_CQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D5 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D6 = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_D1 = CLBLM_R_X5Y133_SLICE_X7Y133_BQ;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_T1 = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_D1 = CLBLM_R_X7Y133_SLICE_X9Y133_BQ;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_T1 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_B2 = CLBLL_L_X4Y132_SLICE_X4Y132_CQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_B3 = CLBLL_L_X4Y137_SLICE_X4Y137_AO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A4 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO2;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A5 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A6 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B2 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B3 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B4 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B5 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B6 = 1'b1;
  assign LIOI3_X0Y211_ILOGIC_X0Y212_D = LIOB33_X0Y211_IOB_X0Y212_I;
  assign LIOI3_X0Y211_ILOGIC_X0Y211_D = LIOB33_X0Y211_IOB_X0Y211_I;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C2 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_A3 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C3 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_A4 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_A5 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_A6 = 1'b1;
  assign LIOI3_X0Y89_ILOGIC_X0Y90_D = LIOB33_X0Y89_IOB_X0Y90_I;
  assign LIOI3_X0Y89_ILOGIC_X0Y89_D = LIOB33_X0Y89_IOB_X0Y89_I;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_AX = LIOB33_X0Y207_IOB_X0Y208_I;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A1 = BRAM_R_X17Y135_RAMB18_X1Y54_DO22;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A2 = CLBLM_R_X3Y132_SLICE_X2Y132_DQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A3 = BRAM_L_X6Y135_RAMB18_X0Y54_DO23;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_B1 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A4 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO7;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A5 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO7;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A6 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO6;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_B2 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B1 = BRAM_L_X6Y135_RAMB18_X0Y54_DO22;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B2 = CLBLL_L_X4Y133_SLICE_X5Y133_AQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B3 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO7;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_B3 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B4 = BRAM_R_X17Y135_RAMB18_X1Y54_DO23;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B5 = BRAM_L_X6Y135_RAMB18_X0Y54_DO23;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B6 = BRAM_L_X6Y130_RAMB18_X0Y53_DOADO6;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_B4 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y231_ILOGIC_X0Y232_D = LIOB33_X0Y231_IOB_X0Y232_I;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C1 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO4;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C3 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO4;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C4 = CLBLM_R_X5Y131_SLICE_X6Y131_A5Q;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C5 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO3;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C6 = BRAM_L_X6Y140_RAMB18_X0Y56_DO20;
  assign LIOI3_TBYTESRC_X0Y231_ILOGIC_X0Y231_D = LIOB33_X0Y231_IOB_X0Y231_I;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_B5 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C2 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO3;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_B6 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D1 = CLBLM_R_X7Y135_SLICE_X9Y135_AO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D2 = CLBLM_R_X3Y132_SLICE_X2Y132_DQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D3 = CLBLL_L_X4Y156_SLICE_X5Y156_CQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D4 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D5 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D6 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_BX = LIOB33_X0Y227_IOB_X0Y228_I;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A1 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A2 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO7;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A3 = CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A4 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO7;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A5 = CLBLM_R_X3Y147_SLICE_X2Y147_AQ;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_C1 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A6 = CLBLM_R_X5Y131_SLICE_X6Y131_A5Q;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_C2 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B1 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B2 = CLBLM_R_X7Y134_SLICE_X9Y134_CO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B3 = CLBLL_L_X4Y131_SLICE_X5Y131_AQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B4 = CLBLM_R_X3Y158_SLICE_X2Y158_AQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B5 = BRAM_L_X6Y135_RAMB18_X0Y54_DO23;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B6 = BRAM_L_X6Y125_RAMB18_X0Y51_DOADO7;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_C3 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_C4 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C1 = CLBLM_R_X3Y130_SLICE_X3Y130_AQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C2 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C3 = CLBLM_R_X3Y157_SLICE_X2Y157_AQ;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_C5 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C4 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C5 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C6 = CLBLM_R_X7Y134_SLICE_X8Y134_BO6;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_C6 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_CE = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D1 = CLBLM_R_X3Y158_SLICE_X3Y158_DQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D2 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D3 = CLBLM_R_X7Y132_SLICE_X9Y132_BO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D4 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D5 = CLBLL_L_X4Y129_SLICE_X5Y129_AQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D6 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_CX = LIOB33_X0Y229_IOB_X0Y229_I;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_D1 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_D2 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_D3 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A1 = BRAM_R_X17Y135_RAMB18_X1Y54_DO2;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A2 = CLBLM_R_X7Y129_SLICE_X8Y129_B5Q;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A3 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO2;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A4 = BRAM_L_X6Y135_RAMB18_X0Y54_DO1;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A5 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO1;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A6 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO2;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B1 = BRAM_R_X17Y135_RAMB18_X1Y54_DO0;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B2 = BRAM_R_X17Y135_RAMB18_X1Y55_DOBDO0;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B3 = BRAM_L_X6Y135_RAMB18_X0Y54_DO0;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B4 = CLBLM_R_X7Y127_SLICE_X8Y127_A5Q;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B5 = BRAM_R_X17Y135_RAMB18_X1Y54_DO7;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B6 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO7;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C1 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C2 = CLBLL_L_X4Y156_SLICE_X5Y156_AQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C3 = CLBLL_L_X4Y133_SLICE_X5Y133_AQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C4 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C5 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C6 = CLBLM_R_X7Y135_SLICE_X9Y135_BO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D1 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D2 = CLBLM_R_X7Y129_SLICE_X8Y129_B5Q;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D3 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D4 = CLBLM_R_X7Y136_SLICE_X9Y136_AO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D5 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D6 = CLBLM_R_X25Y151_SLICE_X36Y151_AQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A1 = BRAM_L_X6Y125_RAMB18_X0Y50_DO17;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A2 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A3 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A4 = BRAM_L_X6Y135_RAMB18_X0Y54_DO1;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A5 = CLBLM_R_X7Y136_SLICE_X8Y136_A5Q;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A6 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B1 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B2 = BRAM_L_X6Y140_RAMB18_X0Y56_DO4;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B3 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B4 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B5 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B6 = CLBLM_R_X3Y133_SLICE_X3Y133_BQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C1 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C2 = BRAM_L_X6Y140_RAMB18_X0Y57_DOBDO7;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C3 = CLBLM_L_X8Y136_SLICE_X10Y136_DO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C4 = BRAM_R_X17Y135_RAMB18_X1Y54_DO7;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C5 = CLBLM_R_X7Y125_SLICE_X8Y125_B5Q;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C6 = CLBLL_L_X4Y156_SLICE_X5Y156_A5Q;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D1 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D2 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D3 = CLBLM_R_X7Y136_SLICE_X9Y136_BO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D4 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D5 = CLBLL_L_X4Y156_SLICE_X5Y156_DQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D6 = CLBLM_R_X7Y127_SLICE_X8Y127_A5Q;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_D2 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_D3 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_D4 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_D5 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_D6 = 1'b1;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_D1 = CLBLM_R_X5Y135_SLICE_X7Y135_AQ;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_T1 = 1'b1;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_D1 = CLBLM_R_X7Y137_SLICE_X9Y137_AQ;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_T1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A2 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A3 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A4 = CLBLM_R_X5Y126_SLICE_X6Y126_BQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A5 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A6 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO3;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B2 = CLBLM_R_X5Y131_SLICE_X6Y131_CQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B3 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO0;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B4 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B5 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B6 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C2 = BRAM_L_X6Y140_RAMB18_X0Y56_DO1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C3 = CLBLL_L_X4Y132_SLICE_X4Y132_CQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C4 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C5 = 1'b1;
  assign BRAM_R_X17Y135_RAMB18_X1Y55_DIADI0 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C6 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D1 = BRAM_L_X6Y140_RAMB18_X0Y56_DO7;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D2 = CLBLM_R_X3Y132_SLICE_X3Y132_CQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D3 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D4 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D5 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D6 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A1 = LIOB33_X0Y129_IOB_X0Y130_I;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A2 = CLBLM_R_X7Y137_SLICE_X8Y137_A5Q;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A3 = BRAM_L_X6Y135_RAMB18_X0Y54_DO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A4 = BRAM_L_X6Y125_RAMB18_X0Y50_DO22;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A5 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A6 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B2 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B3 = BRAM_L_X6Y125_RAMB18_X0Y51_DOBDO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B4 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B5 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B6 = CLBLL_L_X4Y127_SLICE_X5Y127_AQ;
  assign LIOI3_X0Y215_ILOGIC_X0Y216_D = LIOB33_X0Y215_IOB_X0Y216_I;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C1 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO4;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C2 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO4;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C3 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO5;
  assign LIOI3_X0Y215_ILOGIC_X0Y215_D = LIOB33_X0Y215_IOB_X0Y215_I;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C5 = BRAM_L_X6Y140_RAMB18_X0Y56_DO21;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C6 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO5;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C4 = CLBLL_L_X4Y130_SLICE_X5Y130_A5Q;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D1 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D2 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D3 = CLBLM_R_X3Y147_SLICE_X3Y147_BQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D4 = CLBLM_R_X7Y137_SLICE_X8Y137_CO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D5 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D6 = CLBLL_L_X4Y130_SLICE_X5Y130_A5Q;
  assign LIOI3_X0Y91_ILOGIC_X0Y92_D = LIOB33_X0Y91_IOB_X0Y92_I;
  assign LIOI3_X0Y91_ILOGIC_X0Y91_D = LIOB33_X0Y91_IOB_X0Y91_I;
  assign LIOI3_TBYTESRC_X0Y243_ILOGIC_X0Y244_D = LIOB33_X0Y243_IOB_X0Y244_I;
  assign RIOB33_SING_X105Y50_IOB_X1Y50_O = CLBLM_R_X5Y130_SLICE_X7Y130_AQ;
  assign LIOI3_TBYTESRC_X0Y243_ILOGIC_X0Y243_D = LIOB33_X0Y243_IOB_X0Y243_I;
  assign RIOB33_SING_X105Y99_IOB_X1Y99_O = CLBLM_R_X7Y126_SLICE_X8Y126_DQ;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_A1 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_A2 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_A3 = CLBLM_R_X5Y129_SLICE_X7Y129_BQ;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_A4 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO0;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_A5 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_A6 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_B1 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_B2 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO1;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_B3 = CLBLM_R_X5Y129_SLICE_X6Y129_BQ;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_B4 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_B5 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_B6 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_C1 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_C2 = CLBLL_L_X4Y129_SLICE_X5Y129_CQ;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_C3 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_C4 = BRAM_L_X6Y135_RAMB18_X0Y55_DOADO2;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_C5 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_C6 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_D1 = CLBLL_L_X4Y130_SLICE_X4Y130_BQ;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_D2 = BRAM_L_X6Y130_RAMB18_X0Y53_DOBDO1;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_D3 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_D4 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_D5 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_D6 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_A1 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO7;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_A2 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO7;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_A3 = CLBLM_R_X3Y147_SLICE_X3Y147_AQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_A4 = CLBLM_R_X7Y138_SLICE_X8Y138_BO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_A5 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_A6 = CLBLM_R_X5Y130_SLICE_X7Y130_A5Q;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_B1 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO3;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_B2 = BRAM_L_X6Y140_RAMB18_X0Y56_DO20;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_B3 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO4;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_B4 = CLBLM_R_X5Y130_SLICE_X7Y130_A5Q;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_B5 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO4;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_B6 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO3;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_C1 = BRAM_L_X6Y140_RAMB18_X0Y57_DOADO4;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_C2 = BRAM_R_X17Y135_RAMB18_X1Y55_DOADO5;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_C3 = BRAM_L_X6Y140_RAMB18_X0Y56_DO21;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_C4 = CLBLM_R_X5Y127_SLICE_X7Y127_B5Q;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_C5 = BRAM_L_X6Y135_RAMB18_X0Y55_DOBDO5;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_C6 = BRAM_L_X6Y140_RAMB18_X0Y56_DO20;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_D1 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_D2 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_D3 = CLBLM_R_X3Y145_SLICE_X2Y145_BQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_D4 = CLBLM_R_X7Y138_SLICE_X8Y138_CO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_D5 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_D6 = CLBLM_R_X5Y127_SLICE_X7Y127_B5Q;
  assign RIOB33_SING_X105Y100_IOB_X1Y100_O = CLBLL_L_X54Y116_SLICE_X82Y116_AQ;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_DIADI11 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_DIADI12 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_DIADI13 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_DIADI14 = 1'b0;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_DIADI15 = 1'b0;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_B1 = CLBLM_L_X8Y137_SLICE_X10Y137_B5Q;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_DIBDI1 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_B2 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_DIBDI2 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_B3 = CLBLM_L_X16Y154_SLICE_X22Y154_BQ;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_DIBDI3 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_B4 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_C1 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_C2 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_C3 = 1'b1;
  assign BRAM_L_X6Y125_RAMB18_X0Y50_DIBDI14 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_C4 = 1'b1;
endmodule
