module top(
  input RIOB33_SING_X105Y50_IOB_X1Y50_IPAD,
  input RIOB33_X105Y51_IOB_X1Y51_IPAD,
  input RIOB33_X105Y51_IOB_X1Y52_IPAD,
  input RIOB33_X105Y53_IOB_X1Y53_IPAD,
  input RIOB33_X105Y53_IOB_X1Y54_IPAD,
  input RIOB33_X105Y55_IOB_X1Y55_IPAD,
  input RIOB33_X105Y55_IOB_X1Y56_IPAD,
  input RIOB33_X105Y57_IOB_X1Y57_IPAD,
  input RIOB33_X105Y57_IOB_X1Y58_IPAD,
  input RIOB33_X105Y59_IOB_X1Y59_IPAD,
  input RIOB33_X105Y59_IOB_X1Y60_IPAD,
  input RIOB33_X105Y61_IOB_X1Y61_IPAD,
  input RIOB33_X105Y61_IOB_X1Y62_IPAD,
  input RIOB33_X105Y77_IOB_X1Y78_IPAD,
  output LIOB33_SING_X0Y100_IOB_X0Y100_OPAD,
  output LIOB33_SING_X0Y149_IOB_X0Y149_OPAD,
  output LIOB33_SING_X0Y150_IOB_X0Y150_OPAD,
  output LIOB33_SING_X0Y199_IOB_X0Y199_OPAD,
  output LIOB33_SING_X0Y50_IOB_X0Y50_OPAD,
  output LIOB33_SING_X0Y99_IOB_X0Y99_OPAD,
  output LIOB33_X0Y101_IOB_X0Y101_OPAD,
  output LIOB33_X0Y101_IOB_X0Y102_OPAD,
  output LIOB33_X0Y103_IOB_X0Y103_OPAD,
  output LIOB33_X0Y103_IOB_X0Y104_OPAD,
  output LIOB33_X0Y105_IOB_X0Y105_OPAD,
  output LIOB33_X0Y105_IOB_X0Y106_OPAD,
  output LIOB33_X0Y107_IOB_X0Y107_OPAD,
  output LIOB33_X0Y107_IOB_X0Y108_OPAD,
  output LIOB33_X0Y109_IOB_X0Y109_OPAD,
  output LIOB33_X0Y109_IOB_X0Y110_OPAD,
  output LIOB33_X0Y111_IOB_X0Y111_OPAD,
  output LIOB33_X0Y111_IOB_X0Y112_OPAD,
  output LIOB33_X0Y113_IOB_X0Y113_OPAD,
  output LIOB33_X0Y113_IOB_X0Y114_OPAD,
  output LIOB33_X0Y115_IOB_X0Y115_OPAD,
  output LIOB33_X0Y115_IOB_X0Y116_OPAD,
  output LIOB33_X0Y117_IOB_X0Y117_OPAD,
  output LIOB33_X0Y117_IOB_X0Y118_OPAD,
  output LIOB33_X0Y119_IOB_X0Y119_OPAD,
  output LIOB33_X0Y119_IOB_X0Y120_OPAD,
  output LIOB33_X0Y121_IOB_X0Y121_OPAD,
  output LIOB33_X0Y121_IOB_X0Y122_OPAD,
  output LIOB33_X0Y123_IOB_X0Y123_OPAD,
  output LIOB33_X0Y123_IOB_X0Y124_OPAD,
  output LIOB33_X0Y125_IOB_X0Y125_OPAD,
  output LIOB33_X0Y125_IOB_X0Y126_OPAD,
  output LIOB33_X0Y127_IOB_X0Y127_OPAD,
  output LIOB33_X0Y127_IOB_X0Y128_OPAD,
  output LIOB33_X0Y129_IOB_X0Y129_OPAD,
  output LIOB33_X0Y129_IOB_X0Y130_OPAD,
  output LIOB33_X0Y131_IOB_X0Y131_OPAD,
  output LIOB33_X0Y131_IOB_X0Y132_OPAD,
  output LIOB33_X0Y133_IOB_X0Y133_OPAD,
  output LIOB33_X0Y133_IOB_X0Y134_OPAD,
  output LIOB33_X0Y135_IOB_X0Y135_OPAD,
  output LIOB33_X0Y135_IOB_X0Y136_OPAD,
  output LIOB33_X0Y137_IOB_X0Y137_OPAD,
  output LIOB33_X0Y137_IOB_X0Y138_OPAD,
  output LIOB33_X0Y139_IOB_X0Y139_OPAD,
  output LIOB33_X0Y139_IOB_X0Y140_OPAD,
  output LIOB33_X0Y141_IOB_X0Y141_OPAD,
  output LIOB33_X0Y141_IOB_X0Y142_OPAD,
  output LIOB33_X0Y143_IOB_X0Y143_OPAD,
  output LIOB33_X0Y145_IOB_X0Y145_OPAD,
  output LIOB33_X0Y145_IOB_X0Y146_OPAD,
  output LIOB33_X0Y147_IOB_X0Y147_OPAD,
  output LIOB33_X0Y147_IOB_X0Y148_OPAD,
  output LIOB33_X0Y151_IOB_X0Y151_OPAD,
  output LIOB33_X0Y151_IOB_X0Y152_OPAD,
  output LIOB33_X0Y153_IOB_X0Y153_OPAD,
  output LIOB33_X0Y153_IOB_X0Y154_OPAD,
  output LIOB33_X0Y155_IOB_X0Y155_OPAD,
  output LIOB33_X0Y155_IOB_X0Y156_OPAD,
  output LIOB33_X0Y157_IOB_X0Y157_OPAD,
  output LIOB33_X0Y157_IOB_X0Y158_OPAD,
  output LIOB33_X0Y159_IOB_X0Y159_OPAD,
  output LIOB33_X0Y159_IOB_X0Y160_OPAD,
  output LIOB33_X0Y161_IOB_X0Y161_OPAD,
  output LIOB33_X0Y161_IOB_X0Y162_OPAD,
  output LIOB33_X0Y163_IOB_X0Y163_OPAD,
  output LIOB33_X0Y163_IOB_X0Y164_OPAD,
  output LIOB33_X0Y165_IOB_X0Y165_OPAD,
  output LIOB33_X0Y165_IOB_X0Y166_OPAD,
  output LIOB33_X0Y167_IOB_X0Y167_OPAD,
  output LIOB33_X0Y167_IOB_X0Y168_OPAD,
  output LIOB33_X0Y169_IOB_X0Y169_OPAD,
  output LIOB33_X0Y169_IOB_X0Y170_OPAD,
  output LIOB33_X0Y171_IOB_X0Y171_OPAD,
  output LIOB33_X0Y171_IOB_X0Y172_OPAD,
  output LIOB33_X0Y173_IOB_X0Y173_OPAD,
  output LIOB33_X0Y173_IOB_X0Y174_OPAD,
  output LIOB33_X0Y175_IOB_X0Y175_OPAD,
  output LIOB33_X0Y175_IOB_X0Y176_OPAD,
  output LIOB33_X0Y177_IOB_X0Y177_OPAD,
  output LIOB33_X0Y177_IOB_X0Y178_OPAD,
  output LIOB33_X0Y179_IOB_X0Y179_OPAD,
  output LIOB33_X0Y179_IOB_X0Y180_OPAD,
  output LIOB33_X0Y181_IOB_X0Y181_OPAD,
  output LIOB33_X0Y181_IOB_X0Y182_OPAD,
  output LIOB33_X0Y183_IOB_X0Y183_OPAD,
  output LIOB33_X0Y183_IOB_X0Y184_OPAD,
  output LIOB33_X0Y185_IOB_X0Y185_OPAD,
  output LIOB33_X0Y185_IOB_X0Y186_OPAD,
  output LIOB33_X0Y187_IOB_X0Y187_OPAD,
  output LIOB33_X0Y187_IOB_X0Y188_OPAD,
  output LIOB33_X0Y189_IOB_X0Y189_OPAD,
  output LIOB33_X0Y189_IOB_X0Y190_OPAD,
  output LIOB33_X0Y191_IOB_X0Y191_OPAD,
  output LIOB33_X0Y191_IOB_X0Y192_OPAD,
  output LIOB33_X0Y193_IOB_X0Y193_OPAD,
  output LIOB33_X0Y193_IOB_X0Y194_OPAD,
  output LIOB33_X0Y195_IOB_X0Y195_OPAD,
  output LIOB33_X0Y195_IOB_X0Y196_OPAD,
  output LIOB33_X0Y197_IOB_X0Y197_OPAD,
  output LIOB33_X0Y197_IOB_X0Y198_OPAD,
  output LIOB33_X0Y51_IOB_X0Y51_OPAD,
  output LIOB33_X0Y51_IOB_X0Y52_OPAD,
  output LIOB33_X0Y53_IOB_X0Y53_OPAD,
  output LIOB33_X0Y53_IOB_X0Y54_OPAD,
  output LIOB33_X0Y55_IOB_X0Y55_OPAD,
  output LIOB33_X0Y55_IOB_X0Y56_OPAD,
  output LIOB33_X0Y57_IOB_X0Y57_OPAD,
  output LIOB33_X0Y57_IOB_X0Y58_OPAD,
  output LIOB33_X0Y59_IOB_X0Y59_OPAD,
  output LIOB33_X0Y59_IOB_X0Y60_OPAD,
  output LIOB33_X0Y61_IOB_X0Y61_OPAD,
  output LIOB33_X0Y61_IOB_X0Y62_OPAD,
  output LIOB33_X0Y63_IOB_X0Y63_OPAD,
  output LIOB33_X0Y63_IOB_X0Y64_OPAD,
  output LIOB33_X0Y65_IOB_X0Y65_OPAD,
  output LIOB33_X0Y65_IOB_X0Y66_OPAD,
  output LIOB33_X0Y67_IOB_X0Y67_OPAD,
  output LIOB33_X0Y67_IOB_X0Y68_OPAD,
  output LIOB33_X0Y69_IOB_X0Y69_OPAD,
  output LIOB33_X0Y69_IOB_X0Y70_OPAD,
  output LIOB33_X0Y71_IOB_X0Y71_OPAD,
  output LIOB33_X0Y71_IOB_X0Y72_OPAD,
  output LIOB33_X0Y73_IOB_X0Y73_OPAD,
  output LIOB33_X0Y73_IOB_X0Y74_OPAD,
  output LIOB33_X0Y75_IOB_X0Y75_OPAD,
  output LIOB33_X0Y75_IOB_X0Y76_OPAD,
  output LIOB33_X0Y77_IOB_X0Y77_OPAD,
  output LIOB33_X0Y77_IOB_X0Y78_OPAD,
  output LIOB33_X0Y79_IOB_X0Y79_OPAD,
  output LIOB33_X0Y79_IOB_X0Y80_OPAD,
  output LIOB33_X0Y81_IOB_X0Y81_OPAD,
  output LIOB33_X0Y81_IOB_X0Y82_OPAD,
  output LIOB33_X0Y83_IOB_X0Y83_OPAD,
  output LIOB33_X0Y83_IOB_X0Y84_OPAD,
  output LIOB33_X0Y85_IOB_X0Y85_OPAD,
  output LIOB33_X0Y85_IOB_X0Y86_OPAD,
  output LIOB33_X0Y87_IOB_X0Y87_OPAD,
  output LIOB33_X0Y87_IOB_X0Y88_OPAD,
  output LIOB33_X0Y89_IOB_X0Y89_OPAD,
  output LIOB33_X0Y89_IOB_X0Y90_OPAD,
  output LIOB33_X0Y91_IOB_X0Y91_OPAD,
  output LIOB33_X0Y91_IOB_X0Y92_OPAD,
  output LIOB33_X0Y93_IOB_X0Y93_OPAD,
  output LIOB33_X0Y93_IOB_X0Y94_OPAD,
  output LIOB33_X0Y95_IOB_X0Y95_OPAD,
  output LIOB33_X0Y95_IOB_X0Y96_OPAD,
  output LIOB33_X0Y97_IOB_X0Y97_OPAD,
  output LIOB33_X0Y97_IOB_X0Y98_OPAD,
  output RIOB33_SING_X105Y100_IOB_X1Y100_OPAD,
  output RIOB33_SING_X105Y149_IOB_X1Y149_OPAD,
  output RIOB33_SING_X105Y150_IOB_X1Y150_OPAD,
  output RIOB33_SING_X105Y199_IOB_X1Y199_OPAD,
  output RIOB33_X105Y101_IOB_X1Y101_OPAD,
  output RIOB33_X105Y101_IOB_X1Y102_OPAD,
  output RIOB33_X105Y103_IOB_X1Y103_OPAD,
  output RIOB33_X105Y103_IOB_X1Y104_OPAD,
  output RIOB33_X105Y105_IOB_X1Y105_OPAD,
  output RIOB33_X105Y105_IOB_X1Y106_OPAD,
  output RIOB33_X105Y107_IOB_X1Y107_OPAD,
  output RIOB33_X105Y107_IOB_X1Y108_OPAD,
  output RIOB33_X105Y109_IOB_X1Y109_OPAD,
  output RIOB33_X105Y109_IOB_X1Y110_OPAD,
  output RIOB33_X105Y111_IOB_X1Y111_OPAD,
  output RIOB33_X105Y111_IOB_X1Y112_OPAD,
  output RIOB33_X105Y113_IOB_X1Y113_OPAD,
  output RIOB33_X105Y113_IOB_X1Y114_OPAD,
  output RIOB33_X105Y115_IOB_X1Y115_OPAD,
  output RIOB33_X105Y115_IOB_X1Y116_OPAD,
  output RIOB33_X105Y117_IOB_X1Y117_OPAD,
  output RIOB33_X105Y117_IOB_X1Y118_OPAD,
  output RIOB33_X105Y119_IOB_X1Y119_OPAD,
  output RIOB33_X105Y119_IOB_X1Y120_OPAD,
  output RIOB33_X105Y121_IOB_X1Y121_OPAD,
  output RIOB33_X105Y121_IOB_X1Y122_OPAD,
  output RIOB33_X105Y123_IOB_X1Y123_OPAD,
  output RIOB33_X105Y123_IOB_X1Y124_OPAD,
  output RIOB33_X105Y125_IOB_X1Y125_OPAD,
  output RIOB33_X105Y125_IOB_X1Y126_OPAD,
  output RIOB33_X105Y127_IOB_X1Y127_OPAD,
  output RIOB33_X105Y127_IOB_X1Y128_OPAD,
  output RIOB33_X105Y129_IOB_X1Y129_OPAD,
  output RIOB33_X105Y129_IOB_X1Y130_OPAD,
  output RIOB33_X105Y131_IOB_X1Y131_OPAD,
  output RIOB33_X105Y131_IOB_X1Y132_OPAD,
  output RIOB33_X105Y133_IOB_X1Y133_OPAD,
  output RIOB33_X105Y133_IOB_X1Y134_OPAD,
  output RIOB33_X105Y135_IOB_X1Y135_OPAD,
  output RIOB33_X105Y135_IOB_X1Y136_OPAD,
  output RIOB33_X105Y137_IOB_X1Y137_OPAD,
  output RIOB33_X105Y137_IOB_X1Y138_OPAD,
  output RIOB33_X105Y139_IOB_X1Y139_OPAD,
  output RIOB33_X105Y139_IOB_X1Y140_OPAD,
  output RIOB33_X105Y141_IOB_X1Y141_OPAD,
  output RIOB33_X105Y141_IOB_X1Y142_OPAD,
  output RIOB33_X105Y143_IOB_X1Y143_OPAD,
  output RIOB33_X105Y143_IOB_X1Y144_OPAD,
  output RIOB33_X105Y145_IOB_X1Y145_OPAD,
  output RIOB33_X105Y145_IOB_X1Y146_OPAD,
  output RIOB33_X105Y147_IOB_X1Y147_OPAD,
  output RIOB33_X105Y147_IOB_X1Y148_OPAD,
  output RIOB33_X105Y151_IOB_X1Y151_OPAD,
  output RIOB33_X105Y151_IOB_X1Y152_OPAD,
  output RIOB33_X105Y153_IOB_X1Y153_OPAD,
  output RIOB33_X105Y153_IOB_X1Y154_OPAD,
  output RIOB33_X105Y155_IOB_X1Y155_OPAD,
  output RIOB33_X105Y155_IOB_X1Y156_OPAD,
  output RIOB33_X105Y157_IOB_X1Y157_OPAD,
  output RIOB33_X105Y157_IOB_X1Y158_OPAD,
  output RIOB33_X105Y159_IOB_X1Y159_OPAD,
  output RIOB33_X105Y159_IOB_X1Y160_OPAD,
  output RIOB33_X105Y161_IOB_X1Y161_OPAD,
  output RIOB33_X105Y161_IOB_X1Y162_OPAD,
  output RIOB33_X105Y163_IOB_X1Y163_OPAD,
  output RIOB33_X105Y163_IOB_X1Y164_OPAD,
  output RIOB33_X105Y165_IOB_X1Y165_OPAD,
  output RIOB33_X105Y165_IOB_X1Y166_OPAD,
  output RIOB33_X105Y167_IOB_X1Y167_OPAD,
  output RIOB33_X105Y167_IOB_X1Y168_OPAD,
  output RIOB33_X105Y169_IOB_X1Y169_OPAD,
  output RIOB33_X105Y169_IOB_X1Y170_OPAD,
  output RIOB33_X105Y171_IOB_X1Y171_OPAD,
  output RIOB33_X105Y171_IOB_X1Y172_OPAD,
  output RIOB33_X105Y173_IOB_X1Y173_OPAD,
  output RIOB33_X105Y173_IOB_X1Y174_OPAD,
  output RIOB33_X105Y175_IOB_X1Y175_OPAD,
  output RIOB33_X105Y175_IOB_X1Y176_OPAD,
  output RIOB33_X105Y177_IOB_X1Y177_OPAD,
  output RIOB33_X105Y177_IOB_X1Y178_OPAD,
  output RIOB33_X105Y179_IOB_X1Y179_OPAD,
  output RIOB33_X105Y179_IOB_X1Y180_OPAD,
  output RIOB33_X105Y181_IOB_X1Y181_OPAD,
  output RIOB33_X105Y181_IOB_X1Y182_OPAD,
  output RIOB33_X105Y183_IOB_X1Y183_OPAD,
  output RIOB33_X105Y183_IOB_X1Y184_OPAD,
  output RIOB33_X105Y185_IOB_X1Y185_OPAD,
  output RIOB33_X105Y185_IOB_X1Y186_OPAD,
  output RIOB33_X105Y187_IOB_X1Y187_OPAD,
  output RIOB33_X105Y187_IOB_X1Y188_OPAD,
  output RIOB33_X105Y189_IOB_X1Y189_OPAD,
  output RIOB33_X105Y189_IOB_X1Y190_OPAD,
  output RIOB33_X105Y191_IOB_X1Y191_OPAD,
  output RIOB33_X105Y191_IOB_X1Y192_OPAD,
  output RIOB33_X105Y193_IOB_X1Y193_OPAD,
  output RIOB33_X105Y193_IOB_X1Y194_OPAD,
  output RIOB33_X105Y195_IOB_X1Y195_OPAD,
  output RIOB33_X105Y195_IOB_X1Y196_OPAD,
  output RIOB33_X105Y197_IOB_X1Y197_OPAD,
  output RIOB33_X105Y197_IOB_X1Y198_OPAD,
  output RIOB33_X105Y63_IOB_X1Y63_OPAD,
  output RIOB33_X105Y63_IOB_X1Y64_OPAD,
  output RIOB33_X105Y65_IOB_X1Y65_OPAD,
  output RIOB33_X105Y65_IOB_X1Y66_OPAD,
  output RIOB33_X105Y67_IOB_X1Y67_OPAD,
  output RIOB33_X105Y67_IOB_X1Y68_OPAD,
  output RIOB33_X105Y69_IOB_X1Y69_OPAD,
  output RIOB33_X105Y69_IOB_X1Y70_OPAD,
  output RIOB33_X105Y71_IOB_X1Y71_OPAD,
  output RIOB33_X105Y71_IOB_X1Y72_OPAD,
  output RIOB33_X105Y73_IOB_X1Y73_OPAD,
  output RIOB33_X105Y73_IOB_X1Y74_OPAD,
  output RIOB33_X105Y75_IOB_X1Y75_OPAD,
  output RIOB33_X105Y75_IOB_X1Y76_OPAD,
  output RIOB33_X105Y77_IOB_X1Y77_OPAD,
  output RIOB33_X105Y79_IOB_X1Y79_OPAD,
  output RIOB33_X105Y79_IOB_X1Y80_OPAD,
  output RIOB33_X105Y81_IOB_X1Y81_OPAD,
  output RIOB33_X105Y81_IOB_X1Y82_OPAD,
  output RIOB33_X105Y83_IOB_X1Y83_OPAD,
  output RIOB33_X105Y83_IOB_X1Y84_OPAD,
  output RIOB33_X105Y85_IOB_X1Y85_OPAD,
  output RIOB33_X105Y85_IOB_X1Y86_OPAD,
  output RIOB33_X105Y87_IOB_X1Y87_OPAD,
  output RIOB33_X105Y87_IOB_X1Y88_OPAD,
  output RIOB33_X105Y89_IOB_X1Y89_OPAD,
  output RIOB33_X105Y89_IOB_X1Y90_OPAD,
  output RIOB33_X105Y91_IOB_X1Y91_OPAD
  );
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_AO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_AO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_BO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_BO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_CO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_CO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_DO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_DO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_AO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_AO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_BO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_BO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_CO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_CO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_DO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_DO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D_XOR;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_A;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_A1;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_A2;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_A3;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_A4;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_A5;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_A6;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_AO5;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_AO6;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_A_CY;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_A_XOR;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_B;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_B1;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_B2;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_B3;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_B4;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_B5;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_B6;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_BO5;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_BO6;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_B_CY;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_B_XOR;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_C;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_C1;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_C2;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_C3;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_C4;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_C5;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_C6;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_CO5;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_CO6;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_C_CY;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_C_XOR;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_D;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_D1;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_D2;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_D3;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_D4;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_D5;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_D6;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_DO5;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_DO6;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_D_CY;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_D_XOR;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_A;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_A1;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_A2;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_A3;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_A4;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_A5;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_A6;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_AO5;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_AO6;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_A_CY;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_A_XOR;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_B;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_B1;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_B2;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_B3;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_B4;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_B5;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_B6;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_BO5;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_BO6;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_B_CY;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_B_XOR;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_C;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_C1;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_C2;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_C3;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_C4;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_C5;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_C6;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_CO5;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_CO6;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_C_CY;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_C_XOR;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_D;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_D1;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_D2;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_D3;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_D4;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_D5;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_D6;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_DO5;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_DO6;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_D_CY;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_D_XOR;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_A;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_A1;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_A2;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_A3;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_A4;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_A5;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_A6;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_AO5;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_AO6;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_A_CY;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_A_XOR;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_B;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_B1;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_B2;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_B3;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_B4;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_B5;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_B6;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_BO5;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_BO6;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_B_CY;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_B_XOR;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_C;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_C1;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_C2;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_C3;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_C4;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_C5;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_C6;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_CO5;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_CO6;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_C_CY;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_C_XOR;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_D;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_D1;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_D2;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_D3;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_D4;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_D5;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_D6;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_DO5;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_DO6;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_D_CY;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_D_XOR;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_A;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_A1;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_A2;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_A3;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_A4;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_A5;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_A6;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_AO5;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_AO6;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_A_CY;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_A_XOR;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_B;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_B1;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_B2;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_B3;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_B4;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_B5;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_B6;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_BO5;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_BO6;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_B_CY;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_B_XOR;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_C;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_C1;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_C2;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_C3;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_C4;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_C5;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_C6;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_CO5;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_CO6;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_C_CY;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_C_XOR;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_D;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_D1;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_D2;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_D3;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_D4;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_D5;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_D6;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_DO5;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_DO6;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_D_CY;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_D_XOR;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_A;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_A1;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_A2;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_A3;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_A4;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_A5;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_A6;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_AO5;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_A_CY;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_A_XOR;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_B;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_B1;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_B2;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_B3;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_B4;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_B5;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_B6;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_BO5;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_BO6;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_B_CY;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_B_XOR;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_C;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_C1;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_C2;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_C3;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_C4;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_C5;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_C6;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_CO5;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_CO6;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_C_CY;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_C_XOR;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_D;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_D1;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_D2;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_D3;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_D4;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_D5;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_D6;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_DO5;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_DO6;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_D_CY;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_D_XOR;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_A;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_A1;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_A2;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_A3;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_A4;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_A5;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_A6;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_AO5;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_AO6;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_A_CY;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_A_XOR;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_B;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_B1;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_B2;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_B3;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_B4;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_B5;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_B6;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_BO5;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_BO6;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_B_CY;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_B_XOR;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_C;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_C1;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_C2;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_C3;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_C4;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_C5;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_C6;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_CO5;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_CO6;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_C_CY;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_C_XOR;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_D;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_D1;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_D2;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_D3;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_D4;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_D5;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_D6;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_DO5;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_DO6;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_D_CY;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_D_XOR;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_A;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_A1;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_A2;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_A3;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_A4;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_A5;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_A6;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_AMUX;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_AO5;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_AO6;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_A_CY;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_A_XOR;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_B;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_B1;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_B2;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_B3;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_B4;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_B5;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_B6;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_BO5;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_BO6;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_BQ;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_B_CY;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_B_XOR;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_C;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_C1;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_C2;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_C3;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_C4;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_C5;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_C6;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_CLK;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_CO5;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_CO6;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_C_CY;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_C_XOR;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_D;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_D1;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_D2;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_D3;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_D4;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_D5;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_D6;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_DO5;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_DO6;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_D_CY;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_D_XOR;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X106Y100_SR;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_A;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_A1;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_A2;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_A3;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_A4;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_A5;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_A6;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_AO5;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_AO6;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_A_CY;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_A_XOR;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_B;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_B1;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_B2;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_B3;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_B4;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_B5;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_B6;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_BO5;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_BO6;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_B_CY;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_B_XOR;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_C;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_C1;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_C2;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_C3;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_C4;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_C5;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_C6;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_CO5;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_CO6;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_C_CY;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_C_XOR;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_D;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_D1;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_D2;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_D3;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_D4;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_D5;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_D6;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_DO5;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_DO6;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_D_CY;
  wire [0:0] CLBLL_R_X71Y100_SLICE_X107Y100_D_XOR;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_A;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_A1;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_A2;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_A3;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_A4;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_A5;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_A6;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_AO5;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_AO6;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_AQ;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_A_CY;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_A_XOR;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_B;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_B1;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_B2;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_B3;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_B4;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_B5;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_B6;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_BO5;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_BO6;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_BQ;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_B_CY;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_B_XOR;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_C;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_C1;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_C2;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_C3;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_C4;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_C5;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_C6;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_CLK;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_CO5;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_CO6;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_CQ;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_C_CY;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_C_XOR;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_D;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_D1;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_D2;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_D3;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_D4;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_D5;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_D6;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_DO5;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_DO6;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_D_CY;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_D_XOR;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X106Y101_SR;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_A;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_A1;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_A2;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_A3;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_A4;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_A5;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_A6;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_AO5;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_AO6;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_AQ;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_A_CY;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_A_XOR;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_B;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_B1;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_B2;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_B3;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_B4;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_B5;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_B6;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_BO5;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_BO6;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_B_CY;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_B_XOR;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_C;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_C1;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_C2;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_C3;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_C4;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_C5;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_C6;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_CLK;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_CO5;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_CO6;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_C_CY;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_C_XOR;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_D;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_D1;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_D2;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_D3;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_D4;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_D5;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_D6;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_DO5;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_DO6;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_D_CY;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_D_XOR;
  wire [0:0] CLBLL_R_X71Y101_SLICE_X107Y101_SR;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_A;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_A1;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_A2;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_A3;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_A4;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_A5;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_A6;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_AO5;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_AO6;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_AQ;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_A_CY;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_A_XOR;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_B;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_B1;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_B2;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_B3;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_B4;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_B5;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_B6;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_BO5;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_BO6;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_BQ;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_B_CY;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_B_XOR;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_C;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_C1;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_C2;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_C3;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_C4;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_C5;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_C6;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_CLK;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_CO5;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_CO6;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_CQ;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_C_CY;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_C_XOR;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_D;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_D1;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_D2;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_D3;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_D4;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_D5;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_D6;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_DO5;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_DO6;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_D_CY;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_D_XOR;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X106Y102_SR;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_A;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_A1;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_A2;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_A3;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_A4;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_A5;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_A6;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_AO5;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_AO6;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_A_CY;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_A_XOR;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_B;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_B1;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_B2;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_B3;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_B4;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_B5;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_B6;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_BO5;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_BO6;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_B_CY;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_B_XOR;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_C;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_C1;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_C2;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_C3;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_C4;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_C5;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_C6;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_CO5;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_CO6;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_C_CY;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_C_XOR;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_D;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_D1;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_D2;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_D3;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_D4;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_D5;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_D6;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_DO5;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_DO6;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_D_CY;
  wire [0:0] CLBLL_R_X71Y102_SLICE_X107Y102_D_XOR;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_A;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_A1;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_A2;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_A3;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_A4;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_A5;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_A6;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_AO5;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_AO6;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_AQ;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_A_CY;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_A_XOR;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_B;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_B1;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_B2;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_B3;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_B4;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_B5;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_B6;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_BMUX;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_BO5;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_BO6;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_B_CY;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_B_XOR;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_C;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_C1;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_C2;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_C3;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_C4;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_C5;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_C6;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_CLK;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_CO5;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_CO6;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_C_CY;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_C_XOR;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_D;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_D1;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_D2;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_D3;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_D4;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_D5;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_D6;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_DO5;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_DO6;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_D_CY;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_D_XOR;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X106Y103_SR;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_A;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_A1;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_A2;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_A3;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_A4;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_A5;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_A6;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_AO5;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_AO6;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_A_CY;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_A_XOR;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_B;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_B1;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_B2;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_B3;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_B4;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_B5;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_B6;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_BO5;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_BO6;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_B_CY;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_B_XOR;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_C;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_C1;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_C2;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_C3;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_C4;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_C5;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_C6;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_CO5;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_CO6;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_C_CY;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_C_XOR;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_D;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_D1;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_D2;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_D3;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_D4;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_D5;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_D6;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_DO5;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_DO6;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_D_CY;
  wire [0:0] CLBLL_R_X71Y103_SLICE_X107Y103_D_XOR;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_A;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_A1;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_A2;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_A3;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_A4;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_A5;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_A6;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_AO5;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_AO6;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_AQ;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_A_CY;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_A_XOR;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_B;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_B1;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_B2;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_B3;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_B4;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_B5;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_B6;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_BMUX;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_BO5;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_BO6;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_B_CY;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_B_XOR;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_C;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_C1;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_C2;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_C3;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_C4;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_C5;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_C5Q;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_C6;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_CLK;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_CMUX;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_CO5;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_CO6;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_CQ;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_C_CY;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_C_XOR;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_D;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_D1;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_D2;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_D3;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_D4;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_D5;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_D6;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_DO5;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_DO6;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_D_CY;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_D_XOR;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X106Y107_SR;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_A;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_A1;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_A2;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_A3;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_A4;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_A5;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_A6;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_AO5;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_AO6;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_AQ;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_A_CY;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_A_XOR;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_B;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_B1;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_B2;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_B3;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_B4;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_B5;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_B6;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_BO5;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_BO6;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_BQ;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_B_CY;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_B_XOR;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_C;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_C1;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_C2;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_C3;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_C4;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_C5;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_C5Q;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_C6;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_CLK;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_CMUX;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_CO5;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_CO6;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_CQ;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_C_CY;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_C_XOR;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_D;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_D1;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_D2;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_D3;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_D4;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_D5;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_D6;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_DO5;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_DO6;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_D_CY;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_D_XOR;
  wire [0:0] CLBLL_R_X71Y107_SLICE_X107Y107_SR;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_A;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_A1;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_A2;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_A3;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_A4;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_A5;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_A6;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_AO5;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_AO6;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_AQ;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_A_CY;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_A_XOR;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_B;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_B1;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_B2;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_B3;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_B4;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_B5;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_B6;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_BO5;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_BO6;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_BQ;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_B_CY;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_B_XOR;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_C;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_C1;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_C2;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_C3;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_C4;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_C5;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_C6;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_CLK;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_CO5;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_CO6;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_CQ;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_C_CY;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_C_XOR;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_D;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_D1;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_D2;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_D3;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_D4;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_D5;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_D5Q;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_D6;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_DMUX;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_DO5;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_DO6;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_DQ;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_D_CY;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_D_XOR;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X106Y108_SR;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_A;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_A1;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_A2;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_A3;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_A4;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_A5;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_A5Q;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_A6;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_AMUX;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_AO5;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_AO6;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_AQ;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_AX;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_A_CY;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_A_XOR;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_B;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_B1;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_B2;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_B3;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_B4;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_B5;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_B6;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_BO5;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_BO6;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_B_CY;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_B_XOR;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_C;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_C1;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_C2;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_C3;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_C4;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_C5;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_C6;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_CLK;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_CO5;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_CO6;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_C_CY;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_C_XOR;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_D;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_D1;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_D2;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_D3;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_D4;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_D5;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_D6;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_DO5;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_DO6;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_D_CY;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_D_XOR;
  wire [0:0] CLBLL_R_X71Y108_SLICE_X107Y108_SR;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_A;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_A1;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_A2;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_A3;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_A4;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_A5;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_A6;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_AO5;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_AO6;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_AQ;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_A_CY;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_A_XOR;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_B;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_B1;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_B2;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_B3;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_B4;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_B5;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_B5Q;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_B6;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_BMUX;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_BO5;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_BO6;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_BQ;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_B_CY;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_B_XOR;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_C;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_C1;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_C2;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_C3;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_C4;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_C5;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_C6;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_CLK;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_CMUX;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_CO5;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_CO6;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_C_CY;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_C_XOR;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_D;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_D1;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_D2;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_D3;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_D4;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_D5;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_D6;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_DO5;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_DO6;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_D_CY;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_D_XOR;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X106Y109_SR;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_A;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_A1;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_A2;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_A3;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_A4;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_A5;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_A6;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_AO5;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_AO6;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_A_CY;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_A_XOR;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_B;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_B1;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_B2;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_B3;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_B4;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_B5;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_B6;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_BO5;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_BO6;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_B_CY;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_B_XOR;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_C;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_C1;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_C2;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_C3;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_C4;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_C5;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_C6;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_CO5;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_CO6;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_C_CY;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_C_XOR;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_D;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_D1;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_D2;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_D3;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_D4;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_D5;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_D6;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_DO5;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_DO6;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_D_CY;
  wire [0:0] CLBLL_R_X71Y109_SLICE_X107Y109_D_XOR;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_A;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_A1;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_A2;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_A3;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_A4;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_A5;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_A5Q;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_A6;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_AMUX;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_AO5;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_AO6;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_AQ;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_A_CY;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_A_XOR;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_B;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_B1;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_B2;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_B3;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_B4;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_B5;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_B6;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_BO5;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_BO6;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_BQ;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_B_CY;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_B_XOR;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_C;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_C1;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_C2;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_C3;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_C4;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_C5;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_C6;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_CLK;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_CO5;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_CO6;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_C_CY;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_C_XOR;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_D;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_D1;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_D2;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_D3;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_D4;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_D5;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_D6;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_DO5;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_DO6;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_D_CY;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_D_XOR;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X106Y110_SR;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_A;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_A1;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_A2;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_A3;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_A4;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_A5;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_A6;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_AO5;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_AO6;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_A_CY;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_A_XOR;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_B;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_B1;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_B2;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_B3;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_B4;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_B5;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_B6;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_BO5;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_BO6;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_B_CY;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_B_XOR;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_C;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_C1;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_C2;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_C3;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_C4;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_C5;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_C6;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_CO5;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_CO6;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_C_CY;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_C_XOR;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_D;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_D1;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_D2;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_D3;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_D4;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_D5;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_D6;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_DO5;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_DO6;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_D_CY;
  wire [0:0] CLBLL_R_X71Y110_SLICE_X107Y110_D_XOR;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_A;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_A1;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_A2;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_A3;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_A4;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_A5;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_A5Q;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_A6;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_AMUX;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_AO5;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_AO6;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_AQ;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_A_CY;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_A_XOR;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_B;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_B1;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_B2;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_B3;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_B4;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_B5;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_B6;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_BO5;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_BO6;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_BQ;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_B_CY;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_B_XOR;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_C;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_C1;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_C2;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_C3;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_C4;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_C5;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_C6;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_CLK;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_CO5;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_CO6;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_CQ;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_C_CY;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_C_XOR;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_D;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_D1;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_D2;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_D3;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_D4;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_D5;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_D6;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_DO5;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_DO6;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_D_CY;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_D_XOR;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X106Y111_SR;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_A;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_A1;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_A2;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_A3;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_A4;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_A5;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_A6;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_AO5;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_AO6;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_AQ;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_A_CY;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_A_XOR;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_B;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_B1;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_B2;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_B3;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_B4;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_B5;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_B6;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_BO5;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_BO6;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_B_CY;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_B_XOR;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_C;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_C1;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_C2;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_C3;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_C4;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_C5;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_C6;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_CLK;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_CO5;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_CO6;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_C_CY;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_C_XOR;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_D;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_D1;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_D2;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_D3;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_D4;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_D5;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_D6;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_DO5;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_DO6;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_D_CY;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_D_XOR;
  wire [0:0] CLBLL_R_X71Y111_SLICE_X107Y111_SR;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_A;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_A1;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_A2;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_A3;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_A4;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_A5;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_A6;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_AO5;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_AO6;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_AQ;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_A_CY;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_A_XOR;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_B;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_B1;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_B2;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_B3;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_B4;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_B5;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_B5Q;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_B6;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_BMUX;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_BO5;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_BO6;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_BQ;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_B_CY;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_B_XOR;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_C;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_C1;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_C2;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_C3;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_C4;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_C5;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_C6;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_CLK;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_CO5;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_CO6;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_C_CY;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_C_XOR;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_D;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_D1;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_D2;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_D3;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_D4;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_D5;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_D6;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_DO5;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_DO6;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_D_CY;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_D_XOR;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X106Y112_SR;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_A;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_A1;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_A2;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_A3;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_A4;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_A5;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_A6;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_AO5;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_AO6;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_A_CY;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_A_XOR;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_B;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_B1;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_B2;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_B3;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_B4;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_B5;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_B6;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_BO5;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_BO6;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_B_CY;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_B_XOR;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_C;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_C1;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_C2;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_C3;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_C4;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_C5;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_C6;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_CO5;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_CO6;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_C_CY;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_C_XOR;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_D;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_D1;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_D2;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_D3;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_D4;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_D5;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_D6;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_DO5;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_DO6;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_D_CY;
  wire [0:0] CLBLL_R_X71Y112_SLICE_X107Y112_D_XOR;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_A;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_A1;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_A2;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_A3;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_A4;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_A5;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_A6;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_AO5;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_AO6;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_AQ;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_AX;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_A_CY;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_A_XOR;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_B;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_B1;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_B2;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_B3;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_B4;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_B5;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_B6;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_BO5;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_BO6;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_B_CY;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_B_XOR;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_C;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_C1;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_C2;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_C3;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_C4;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_C5;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_C6;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_CLK;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_CO5;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_CO6;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_C_CY;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_C_XOR;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_D;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_D1;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_D2;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_D3;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_D4;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_D5;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_D6;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_DO5;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_DO6;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_D_CY;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_D_XOR;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X106Y114_SR;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_A;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_A1;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_A2;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_A3;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_A4;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_A5;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_A6;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_AO5;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_AO6;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_A_CY;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_A_XOR;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_B;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_B1;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_B2;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_B3;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_B4;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_B5;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_B6;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_BO5;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_BO6;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_B_CY;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_B_XOR;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_C;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_C1;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_C2;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_C3;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_C4;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_C5;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_C6;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_CO5;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_CO6;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_C_CY;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_C_XOR;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_D;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_D1;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_D2;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_D3;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_D4;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_D5;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_D6;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_DO5;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_DO6;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_D_CY;
  wire [0:0] CLBLL_R_X71Y114_SLICE_X107Y114_D_XOR;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_A;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_A1;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_A2;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_A3;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_A4;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_A5;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_A5Q;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_A6;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_AMUX;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_AO5;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_AO6;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_AQ;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_A_CY;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_A_XOR;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_B;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_B1;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_B2;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_B3;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_B4;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_B5;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_B5Q;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_B6;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_BMUX;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_BO5;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_BO6;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_BQ;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_B_CY;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_B_XOR;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_C;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_C1;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_C2;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_C3;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_C4;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_C5;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_C6;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_CLK;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_CO5;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_CO6;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_C_CY;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_C_XOR;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_D;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_D1;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_D2;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_D3;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_D4;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_D5;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_D6;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_DO5;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_DO6;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_D_CY;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_D_XOR;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_SR;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_A;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_A1;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_A2;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_A3;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_A4;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_A5;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_A6;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_AO5;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_AO6;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_A_CY;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_A_XOR;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_B;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_B1;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_B2;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_B3;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_B4;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_B5;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_B6;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_BO5;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_BO6;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_B_CY;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_B_XOR;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_C;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_C1;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_C2;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_C3;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_C4;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_C5;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_C6;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_CO5;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_CO6;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_C_CY;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_C_XOR;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_D;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_D1;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_D2;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_D3;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_D4;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_D5;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_D6;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_DO5;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_DO6;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_D_CY;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_D_XOR;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_A;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_A1;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_A2;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_A3;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_A4;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_A5;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_A5Q;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_A6;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_AMUX;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_AO5;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_AO6;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_AQ;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_A_CY;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_A_XOR;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_B;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_B1;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_B2;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_B3;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_B4;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_B5;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_B6;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_BO5;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_BO6;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_B_CY;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_B_XOR;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_C;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_C1;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_C2;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_C3;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_C4;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_C5;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_C6;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_CLK;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_CO5;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_CO6;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_C_CY;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_C_XOR;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_D;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_D1;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_D2;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_D3;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_D4;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_D5;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_D6;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_DO5;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_DO6;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_D_CY;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_D_XOR;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_SR;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_A;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_A1;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_A2;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_A3;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_A4;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_A5;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_A6;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_AO5;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_AO6;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_A_CY;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_A_XOR;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_B;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_B1;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_B2;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_B3;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_B4;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_B5;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_B6;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_BO5;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_BO6;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_B_CY;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_B_XOR;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_C;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_C1;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_C2;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_C3;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_C4;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_C5;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_C6;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_CO5;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_CO6;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_C_CY;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_C_XOR;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_D;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_D1;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_D2;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_D3;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_D4;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_D5;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_D6;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_DO5;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_DO6;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_D_CY;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_D_XOR;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_A;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_A1;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_A2;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_A3;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_A4;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_A5;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_A5Q;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_A6;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_AMUX;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_AO5;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_AO6;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_AQ;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_AX;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_A_CY;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_A_XOR;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_B;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_B1;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_B2;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_B3;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_B4;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_B5;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_B6;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_BMUX;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_BO5;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_BO6;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_B_CY;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_B_XOR;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_C;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_C1;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_C2;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_C3;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_C4;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_C5;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_C6;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_CLK;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_CO5;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_CO6;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_C_CY;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_C_XOR;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_D;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_D1;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_D2;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_D3;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_D4;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_D5;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_D6;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_DO5;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_DO6;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_D_CY;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_D_XOR;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_SR;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_A;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_A1;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_A2;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_A3;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_A4;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_A5;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_A6;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_AO5;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_AO6;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_A_CY;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_A_XOR;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_B;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_B1;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_B2;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_B3;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_B4;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_B5;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_B6;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_BO5;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_BO6;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_B_CY;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_B_XOR;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_C;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_C1;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_C2;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_C3;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_C4;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_C5;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_C6;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_CO5;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_CO6;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_C_CY;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_C_XOR;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_D;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_D1;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_D2;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_D3;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_D4;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_D5;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_D6;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_DO5;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_DO6;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_D_CY;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_D_XOR;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_A;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_A1;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_A2;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_A3;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_A4;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_A5;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_A5Q;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_A6;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_AMUX;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_AO5;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_AO6;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_AQ;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_A_CY;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_A_XOR;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_B;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_B1;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_B2;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_B3;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_B4;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_B5;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_B6;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_BO5;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_BO6;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_BQ;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_B_CY;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_B_XOR;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_C;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_C1;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_C2;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_C3;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_C4;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_C5;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_C6;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_CLK;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_CO5;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_CO6;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_C_CY;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_C_XOR;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_D;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_D1;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_D2;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_D3;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_D4;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_D5;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_D6;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_DO5;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_DO6;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_D_CY;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_D_XOR;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X106Y124_SR;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_A;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_A1;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_A2;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_A3;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_A4;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_A5;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_A6;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_AO5;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_AO6;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_A_CY;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_A_XOR;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_B;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_B1;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_B2;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_B3;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_B4;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_B5;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_B6;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_BO5;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_BO6;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_B_CY;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_B_XOR;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_C;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_C1;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_C2;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_C3;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_C4;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_C5;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_C6;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_CO5;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_CO6;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_C_CY;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_C_XOR;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_D;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_D1;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_D2;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_D3;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_D4;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_D5;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_D6;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_DO5;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_DO6;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_D_CY;
  wire [0:0] CLBLL_R_X71Y124_SLICE_X107Y124_D_XOR;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_A;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_A1;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_A2;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_A3;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_A4;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_A5;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_A6;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_AO5;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_AO6;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_AQ;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_A_CY;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_A_XOR;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_B;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_B1;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_B2;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_B3;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_B4;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_B5;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_B6;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_BO5;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_BO6;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_BQ;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_B_CY;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_B_XOR;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_C;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_C1;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_C2;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_C3;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_C4;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_C5;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_C6;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_CLK;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_CO5;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_CO6;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_CQ;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_C_CY;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_C_XOR;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_D;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_D1;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_D2;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_D3;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_D4;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_D5;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_D6;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_DO5;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_DO6;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_D_CY;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_D_XOR;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_SR;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_A;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_A1;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_A2;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_A3;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_A4;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_A5;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_A6;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_AO5;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_AO6;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_AQ;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_A_CY;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_A_XOR;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_B;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_B1;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_B2;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_B3;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_B4;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_B5;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_B6;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_BO5;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_BO6;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_B_CY;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_B_XOR;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_C;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_C1;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_C2;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_C3;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_C4;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_C5;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_C6;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_CLK;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_CO5;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_CO6;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_C_CY;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_C_XOR;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_D;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_D1;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_D2;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_D3;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_D4;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_D5;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_D6;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_DO5;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_DO6;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_D_CY;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_D_XOR;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_SR;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_A;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_A1;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_A2;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_A3;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_A4;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_A5;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_A6;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_AO5;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_AO6;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_AQ;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_A_CY;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_A_XOR;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_B;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_B1;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_B2;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_B3;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_B4;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_B5;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_B6;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_BO5;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_BO6;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_BQ;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_B_CY;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_B_XOR;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_C;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_C1;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_C2;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_C3;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_C4;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_C5;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_C6;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_CLK;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_CO5;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_CO6;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_C_CY;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_C_XOR;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_D;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_D1;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_D2;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_D3;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_D4;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_D5;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_D6;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_DO5;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_DO6;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_D_CY;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_D_XOR;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_SR;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_A;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_A1;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_A2;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_A3;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_A4;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_A5;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_A6;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_AMUX;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_AO5;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_AO6;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_AQ;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_A_CY;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_A_XOR;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_B;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_B1;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_B2;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_B3;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_B4;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_B5;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_B6;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_BMUX;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_BO5;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_BO6;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_BQ;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_B_CY;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_B_XOR;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_C;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_C1;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_C2;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_C3;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_C4;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_C5;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_C6;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_CLK;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_CO5;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_CO6;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_C_CY;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_C_XOR;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_D;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_D1;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_D2;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_D3;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_D4;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_D5;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_D6;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_DO5;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_DO6;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_D_CY;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_D_XOR;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_SR;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_A;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_A1;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_A2;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_A3;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_A4;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_A5;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_A6;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_AO5;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_AO6;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_A_CY;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_A_XOR;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_B;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_B1;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_B2;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_B3;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_B4;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_B5;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_B6;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_BO5;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_BO6;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_B_CY;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_B_XOR;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_C;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_C1;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_C2;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_C3;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_C4;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_C5;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_C6;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_CO5;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_CO6;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_C_CY;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_C_XOR;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_D;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_D1;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_D2;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_D3;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_D4;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_D5;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_D6;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_DO5;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_DO6;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_D_CY;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_D_XOR;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_A;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_A1;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_A2;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_A3;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_A4;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_A5;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_A6;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_AMUX;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_AO5;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_AO6;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_AQ;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_A_CY;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_A_XOR;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_B;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_B1;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_B2;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_B3;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_B4;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_B5;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_B6;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_BO5;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_BO6;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_BQ;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_B_CY;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_B_XOR;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_C;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_C1;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_C2;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_C3;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_C4;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_C5;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_C6;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_CLK;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_CO5;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_CO6;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_CQ;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_C_CY;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_C_XOR;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_D;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_D1;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_D2;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_D3;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_D4;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_D5;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_D6;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_DO5;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_DO6;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_DQ;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_D_CY;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_D_XOR;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_SR;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_A;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_A1;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_A2;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_A3;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_A4;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_A5;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_A6;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_AO5;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_AO6;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_AQ;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_A_CY;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_A_XOR;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_B;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_B1;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_B2;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_B3;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_B4;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_B5;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_B6;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_BO5;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_BO6;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_BQ;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_B_CY;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_B_XOR;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_C;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_C1;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_C2;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_C3;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_C4;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_C5;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_C6;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_CLK;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_CO5;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_CO6;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_C_CY;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_C_XOR;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_D;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_D1;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_D2;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_D3;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_D4;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_D5;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_D6;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_DO5;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_DO6;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_D_CY;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_D_XOR;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_SR;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_A;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_A1;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_A2;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_A3;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_A4;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_A5;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_A6;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_AO5;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_AO6;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_A_CY;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_A_XOR;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_B;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_B1;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_B2;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_B3;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_B4;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_B5;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_B6;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_BO5;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_BO6;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_B_CY;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_B_XOR;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_C;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_C1;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_C2;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_C3;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_C4;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_C5;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_C6;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_CO5;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_CO6;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_C_CY;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_C_XOR;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_D;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_D1;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_D2;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_D3;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_D4;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_D5;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_D6;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_DO5;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_DO6;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_D_CY;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_D_XOR;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_A;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_A1;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_A2;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_A3;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_A4;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_A5;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_A6;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_AMUX;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_AO5;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_AO6;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_AQ;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_A_CY;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_A_XOR;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_B;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_B1;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_B2;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_B3;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_B4;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_B5;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_B6;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_BO5;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_BO6;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_BQ;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_B_CY;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_B_XOR;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_C;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_C1;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_C2;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_C3;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_C4;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_C5;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_C6;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_CLK;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_CO5;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_CO6;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_CQ;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_C_CY;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_C_XOR;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_D;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_D1;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_D2;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_D3;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_D4;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_D5;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_D6;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_DO5;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_DO6;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_D_CY;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_D_XOR;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_SR;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_A;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_A1;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_A2;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_A3;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_A4;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_A5;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_A6;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_AO5;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_AO6;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_AQ;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_AX;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_A_CY;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_A_XOR;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_B;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_B1;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_B2;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_B3;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_B4;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_B5;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_B6;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_BO5;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_BO6;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_BQ;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_BX;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_B_CY;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_B_XOR;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_C;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_C1;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_C2;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_C3;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_C4;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_C5;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_C6;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_CE;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_CLK;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_CO5;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_CO6;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_C_CY;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_C_XOR;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_D;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_D1;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_D2;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_D3;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_D4;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_D5;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_D6;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_DO5;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_DO6;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_D_CY;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_D_XOR;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_SR;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_A;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_A1;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_A2;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_A3;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_A4;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_A5;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_A6;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_AO5;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_AO6;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_AQ;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_A_CY;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_A_XOR;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_B;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_B1;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_B2;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_B3;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_B4;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_B5;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_B6;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_BO5;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_BO6;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_BQ;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_B_CY;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_B_XOR;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_C;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_C1;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_C2;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_C3;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_C4;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_C5;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_C6;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_CLK;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_CO5;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_CO6;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_CQ;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_C_CY;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_C_XOR;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_D;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_D1;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_D2;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_D3;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_D4;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_D5;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_D6;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_DMUX;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_DO5;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_DO6;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_D_CY;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_D_XOR;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X106Y130_SR;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_A;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_A1;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_A2;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_A3;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_A4;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_A5;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_A6;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_AO5;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_AO6;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_AQ;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_AX;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_A_CY;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_A_XOR;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_B;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_B1;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_B2;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_B3;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_B4;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_B5;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_B6;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_BO5;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_BO6;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_BQ;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_BX;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_B_CY;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_B_XOR;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_C;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_C1;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_C2;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_C3;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_C4;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_C5;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_C6;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_CE;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_CLK;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_CO5;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_CO6;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_C_CY;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_C_XOR;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_D;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_D1;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_D2;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_D3;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_D4;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_D5;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_D6;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_DO5;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_DO6;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_D_CY;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_D_XOR;
  wire [0:0] CLBLL_R_X71Y130_SLICE_X107Y130_SR;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_A;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_A1;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_A2;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_A3;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_A4;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_A5;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_A6;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_AO5;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_AO6;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_AQ;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_A_CY;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_A_XOR;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_B;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_B1;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_B2;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_B3;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_B4;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_B5;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_B6;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_BO5;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_BO6;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_BQ;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_B_CY;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_B_XOR;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_C;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_C1;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_C2;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_C3;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_C4;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_C5;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_C6;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_CLK;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_CO5;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_CO6;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_CQ;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_C_CY;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_C_XOR;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_D;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_D1;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_D2;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_D3;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_D4;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_D5;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_D6;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_DO5;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_DO6;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_D_CY;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_D_XOR;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_SR;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_A;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_A1;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_A2;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_A3;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_A4;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_A5;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_A5Q;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_A6;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_AMUX;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_AO5;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_AO6;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_AQ;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_AX;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_A_CY;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_A_XOR;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_B;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_B1;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_B2;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_B3;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_B4;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_B5;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_B6;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_BO5;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_BO6;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_BQ;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_B_CY;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_B_XOR;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_C;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_C1;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_C2;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_C3;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_C4;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_C5;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_C6;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_CLK;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_CO5;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_CO6;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_CQ;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_C_CY;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_C_XOR;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_D;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_D1;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_D2;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_D3;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_D4;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_D5;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_D6;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_DMUX;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_DO5;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_DO6;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_D_CY;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_D_XOR;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_SR;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_A;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_A1;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_A2;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_A3;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_A4;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_A5;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_A6;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_AMUX;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_AO5;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_AO6;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_AQ;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_A_CY;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_A_XOR;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_B;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_B1;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_B2;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_B3;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_B4;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_B5;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_B6;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_BO5;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_BO6;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_BQ;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_B_CY;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_B_XOR;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_C;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_C1;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_C2;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_C3;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_C4;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_C5;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_C6;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_CLK;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_CO5;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_CO6;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_CQ;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_C_CY;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_C_XOR;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_D;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_D1;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_D2;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_D3;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_D4;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_D5;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_D6;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_DO5;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_DO6;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_DQ;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_D_CY;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_D_XOR;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X106Y132_SR;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_A;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_A1;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_A2;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_A3;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_A4;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_A5;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_A6;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_AO5;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_AO6;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_AQ;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_A_CY;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_A_XOR;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_B;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_B1;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_B2;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_B3;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_B4;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_B5;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_B6;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_BO5;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_BO6;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_BQ;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_B_CY;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_B_XOR;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_C;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_C1;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_C2;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_C3;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_C4;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_C5;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_C6;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_CLK;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_CO5;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_CO6;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_CQ;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_C_CY;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_C_XOR;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_D;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_D1;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_D2;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_D3;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_D4;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_D5;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_D6;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_DO5;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_DO6;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_DQ;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_D_CY;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_D_XOR;
  wire [0:0] CLBLL_R_X71Y132_SLICE_X107Y132_SR;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_A;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_A1;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_A2;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_A3;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_A4;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_A5;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_A6;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_AO5;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_AO6;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_AQ;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_A_CY;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_A_XOR;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_B;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_B1;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_B2;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_B3;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_B4;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_B5;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_B6;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_BO5;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_BO6;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_BQ;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_B_CY;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_B_XOR;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_C;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_C1;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_C2;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_C3;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_C4;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_C5;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_C6;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_CLK;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_CO5;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_CO6;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_CQ;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_C_CY;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_C_XOR;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_D;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_D1;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_D2;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_D3;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_D4;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_D5;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_D6;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_DO5;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_DO6;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_DQ;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_D_CY;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_D_XOR;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X106Y133_SR;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_A;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_A1;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_A2;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_A3;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_A4;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_A5;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_A6;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_AO5;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_AO6;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_AQ;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_A_CY;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_A_XOR;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_B;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_B1;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_B2;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_B3;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_B4;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_B5;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_B6;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_BO5;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_BO6;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_BQ;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_B_CY;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_B_XOR;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_C;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_C1;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_C2;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_C3;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_C4;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_C5;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_C6;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_CLK;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_CMUX;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_CO5;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_CO6;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_C_CY;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_C_XOR;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_D;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_D1;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_D2;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_D3;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_D4;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_D5;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_D6;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_DO5;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_DO6;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_D_CY;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_D_XOR;
  wire [0:0] CLBLL_R_X71Y133_SLICE_X107Y133_SR;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_A;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_A1;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_A2;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_A3;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_A4;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_A5;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_A6;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_AO5;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_AO6;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_AQ;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_A_CY;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_A_XOR;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_B;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_B1;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_B2;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_B3;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_B4;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_B5;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_B6;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_BO5;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_BO6;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_BQ;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_B_CY;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_B_XOR;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_C;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_C1;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_C2;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_C3;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_C4;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_C5;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_C6;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_CLK;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_CO5;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_CO6;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_C_CY;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_C_XOR;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_D;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_D1;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_D2;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_D3;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_D4;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_D5;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_D6;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_DO5;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_DO6;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_D_CY;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_D_XOR;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X106Y134_SR;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_A;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_A1;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_A2;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_A3;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_A4;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_A5;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_A6;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_AO5;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_AO6;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_AQ;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_A_CY;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_A_XOR;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_B;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_B1;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_B2;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_B3;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_B4;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_B5;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_B6;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_BO5;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_BO6;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_BQ;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_B_CY;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_B_XOR;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_C;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_C1;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_C2;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_C3;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_C4;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_C5;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_C6;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_CLK;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_CO5;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_CO6;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_CQ;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_C_CY;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_C_XOR;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_D;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_D1;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_D2;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_D3;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_D4;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_D5;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_D6;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_DO5;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_DO6;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_D_CY;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_D_XOR;
  wire [0:0] CLBLL_R_X71Y134_SLICE_X107Y134_SR;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_A;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_A1;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_A2;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_A3;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_A4;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_A5;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_A5Q;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_A6;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_AMUX;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_AO5;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_AO6;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_AQ;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_A_CY;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_A_XOR;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_B;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_B1;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_B2;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_B3;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_B4;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_B5;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_B6;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_BO5;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_BO6;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_B_CY;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_B_XOR;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_C;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_C1;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_C2;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_C3;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_C4;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_C5;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_C6;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_CLK;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_CO5;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_CO6;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_C_CY;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_C_XOR;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_D;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_D1;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_D2;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_D3;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_D4;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_D5;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_D6;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_DO5;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_DO6;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_D_CY;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_D_XOR;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X106Y98_SR;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_A;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_A1;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_A2;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_A3;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_A4;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_A5;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_A6;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_AO5;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_AO6;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_A_CY;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_A_XOR;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_B;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_B1;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_B2;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_B3;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_B4;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_B5;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_B6;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_BO5;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_BO6;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_B_CY;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_B_XOR;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_C;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_C1;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_C2;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_C3;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_C4;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_C5;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_C6;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_CO5;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_CO6;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_C_CY;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_C_XOR;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_D;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_D1;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_D2;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_D3;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_D4;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_D5;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_D6;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_DO5;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_DO6;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_D_CY;
  wire [0:0] CLBLL_R_X71Y98_SLICE_X107Y98_D_XOR;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_A;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_A1;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_A2;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_A3;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_A4;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_A5;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_A6;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_AO5;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_AO6;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_AQ;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_A_CY;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_A_XOR;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_B;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_B1;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_B2;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_B3;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_B4;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_B5;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_B6;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_BO5;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_BO6;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_B_CY;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_B_XOR;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_C;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_C1;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_C2;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_C3;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_C4;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_C5;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_C6;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_CLK;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_CO5;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_CO6;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_C_CY;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_C_XOR;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_D;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_D1;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_D2;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_D3;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_D4;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_D5;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_D6;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_DO5;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_DO6;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_D_CY;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_D_XOR;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X110Y101_SR;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_A;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_A1;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_A2;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_A3;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_A4;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_A5;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_A6;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_AO5;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_AO6;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_A_CY;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_A_XOR;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_B;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_B1;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_B2;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_B3;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_B4;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_B5;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_B6;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_BO5;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_BO6;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_B_CY;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_B_XOR;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_C;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_C1;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_C2;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_C3;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_C4;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_C5;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_C6;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_CO5;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_CO6;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_C_CY;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_C_XOR;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_D;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_D1;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_D2;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_D3;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_D4;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_D5;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_D6;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_DO5;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_DO6;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_D_CY;
  wire [0:0] CLBLL_R_X73Y101_SLICE_X111Y101_D_XOR;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_A;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_A1;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_A2;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_A3;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_A4;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_A5;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_A5Q;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_A6;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_AMUX;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_AO5;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_AO6;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_AQ;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_AX;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_A_CY;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_A_XOR;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_B;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_B1;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_B2;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_B3;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_B4;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_B5;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_B6;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_BO5;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_BO6;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_BQ;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_B_CY;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_B_XOR;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_C;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_C1;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_C2;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_C3;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_C4;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_C5;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_C6;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_CLK;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_CO5;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_CO6;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_CQ;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_C_CY;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_C_XOR;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_D;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_D1;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_D2;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_D3;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_D4;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_D5;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_D6;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_DO5;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_DO6;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_D_CY;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_D_XOR;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X110Y102_SR;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_A;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_A1;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_A2;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_A3;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_A4;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_A5;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_A5Q;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_A6;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_AMUX;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_AO5;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_AO6;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_AQ;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_AX;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_A_CY;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_A_XOR;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_B;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_B1;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_B2;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_B3;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_B4;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_B5;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_B6;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_BO5;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_BO6;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_B_CY;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_B_XOR;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_C;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_C1;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_C2;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_C3;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_C4;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_C5;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_C6;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_CLK;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_CO5;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_CO6;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_C_CY;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_C_XOR;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_D;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_D1;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_D2;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_D3;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_D4;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_D5;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_D6;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_DO5;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_DO6;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_D_CY;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_D_XOR;
  wire [0:0] CLBLL_R_X73Y102_SLICE_X111Y102_SR;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_A;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_A1;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_A2;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_A3;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_A4;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_A5;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_A5Q;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_A6;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_AMUX;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_AO5;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_AO6;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_AQ;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_AX;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_A_CY;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_A_XOR;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_B;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_B1;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_B2;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_B3;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_B4;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_B5;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_B5Q;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_B6;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_BMUX;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_BO5;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_BO6;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_BQ;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_BX;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_B_CY;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_B_XOR;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_C;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_C1;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_C2;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_C3;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_C4;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_C5;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_C6;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_CLK;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_CMUX;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_CO5;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_CO6;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_C_CY;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_C_XOR;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_D;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_D1;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_D2;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_D3;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_D4;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_D5;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_D6;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_DMUX;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_DO5;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_DO6;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_D_CY;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_D_XOR;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X110Y103_SR;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_A;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_A1;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_A2;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_A3;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_A4;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_A5;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_A5Q;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_A6;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_AMUX;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_AO5;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_AO6;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_AQ;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_AX;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_A_CY;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_A_XOR;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_B;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_B1;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_B2;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_B3;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_B4;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_B5;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_B6;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_BO5;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_BO6;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_B_CY;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_B_XOR;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_C;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_C1;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_C2;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_C3;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_C4;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_C5;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_C6;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_CLK;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_CO5;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_CO6;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_C_CY;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_C_XOR;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_D;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_D1;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_D2;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_D3;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_D4;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_D5;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_D6;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_DO5;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_DO6;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_D_CY;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_D_XOR;
  wire [0:0] CLBLL_R_X73Y103_SLICE_X111Y103_SR;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_A;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_A1;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_A2;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_A3;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_A4;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_A5;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_A5Q;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_A6;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_AMUX;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_AO5;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_AO6;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_AQ;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_A_CY;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_A_XOR;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_B;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_B1;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_B2;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_B3;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_B4;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_B5;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_B6;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_BMUX;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_BO5;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_BO6;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_BQ;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_B_CY;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_B_XOR;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_C;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_C1;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_C2;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_C3;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_C4;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_C5;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_C6;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_CLK;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_CO5;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_CO6;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_CQ;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_C_CY;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_C_XOR;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_D;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_D1;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_D2;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_D3;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_D4;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_D5;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_D6;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_DMUX;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_DO5;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_DO6;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_D_CY;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_D_XOR;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X110Y104_SR;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_A;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_A1;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_A2;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_A3;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_A4;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_A5;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_A6;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_AO5;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_AO6;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_AQ;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_A_CY;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_A_XOR;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_B;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_B1;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_B2;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_B3;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_B4;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_B5;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_B6;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_BO5;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_BO6;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_BQ;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_B_CY;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_B_XOR;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_C;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_C1;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_C2;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_C3;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_C4;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_C5;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_C6;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_CLK;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_CO5;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_CO6;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_C_CY;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_C_XOR;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_D;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_D1;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_D2;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_D3;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_D4;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_D5;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_D6;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_DMUX;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_DO5;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_DO6;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_D_CY;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_D_XOR;
  wire [0:0] CLBLL_R_X73Y104_SLICE_X111Y104_SR;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_A;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_A1;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_A2;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_A3;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_A4;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_A5;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_A6;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_AO5;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_AO6;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_A_CY;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_A_XOR;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_B;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_B1;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_B2;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_B3;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_B4;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_B5;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_B6;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_BO5;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_BO6;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_B_CY;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_B_XOR;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_C;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_C1;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_C2;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_C3;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_C4;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_C5;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_C6;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_CO5;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_CO6;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_C_CY;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_C_XOR;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_D;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_D1;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_D2;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_D3;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_D4;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_D5;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_D6;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_DO5;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_DO6;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_D_CY;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X110Y106_D_XOR;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_A;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_A1;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_A2;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_A3;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_A4;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_A5;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_A6;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_AO5;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_AO6;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_A_CY;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_A_XOR;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_B;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_B1;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_B2;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_B3;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_B4;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_B5;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_B6;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_BO5;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_BO6;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_B_CY;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_B_XOR;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_C;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_C1;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_C2;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_C3;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_C4;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_C5;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_C6;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_CO5;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_CO6;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_C_CY;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_C_XOR;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_D;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_D1;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_D2;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_D3;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_D4;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_D5;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_D6;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_DO5;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_DO6;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_D_CY;
  wire [0:0] CLBLL_R_X73Y106_SLICE_X111Y106_D_XOR;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_A;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_A1;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_A2;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_A3;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_A4;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_A5;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_A6;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_AO5;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_AO6;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_AQ;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_A_CY;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_A_XOR;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_B;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_B1;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_B2;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_B3;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_B4;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_B5;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_B6;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_BO5;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_BO6;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_BQ;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_B_CY;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_B_XOR;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_C;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_C1;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_C2;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_C3;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_C4;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_C5;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_C6;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_CLK;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_CO5;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_CO6;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_C_CY;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_C_XOR;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_D;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_D1;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_D2;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_D3;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_D4;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_D5;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_D6;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_DO5;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_DO6;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_D_CY;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_D_XOR;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X110Y107_SR;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_A;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_A1;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_A2;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_A3;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_A4;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_A5;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_A6;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_AO5;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_AO6;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_AQ;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_A_CY;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_A_XOR;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_B;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_B1;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_B2;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_B3;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_B4;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_B5;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_B6;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_BO5;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_BO6;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_BQ;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_B_CY;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_B_XOR;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_C;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_C1;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_C2;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_C3;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_C4;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_C5;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_C6;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_CLK;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_CO5;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_CO6;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_CQ;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_C_CY;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_C_XOR;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_D;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_D1;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_D2;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_D3;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_D4;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_D5;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_D6;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_DO5;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_DO6;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_DQ;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_D_CY;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_D_XOR;
  wire [0:0] CLBLL_R_X73Y107_SLICE_X111Y107_SR;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_A;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_A1;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_A2;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_A3;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_A4;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_A5;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_A5Q;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_A6;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_AMUX;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_AO5;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_AO6;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_AQ;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_A_CY;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_A_XOR;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_B;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_B1;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_B2;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_B3;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_B4;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_B5;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_B6;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_BO5;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_BO6;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_BQ;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_B_CY;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_B_XOR;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_C;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_C1;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_C2;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_C3;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_C4;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_C5;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_C6;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_CLK;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_CO5;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_CO6;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_C_CY;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_C_XOR;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_D;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_D1;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_D2;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_D3;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_D4;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_D5;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_D6;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_DO5;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_DO6;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_D_CY;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_D_XOR;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X110Y108_SR;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_A;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_A1;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_A2;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_A3;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_A4;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_A5;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_A6;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_AO5;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_AO6;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_A_CY;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_A_XOR;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_B;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_B1;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_B2;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_B3;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_B4;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_B5;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_B6;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_BO5;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_BO6;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_B_CY;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_B_XOR;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_C;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_C1;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_C2;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_C3;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_C4;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_C5;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_C6;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_CO5;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_CO6;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_C_CY;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_C_XOR;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_D;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_D1;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_D2;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_D3;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_D4;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_D5;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_D6;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_DO5;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_DO6;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_D_CY;
  wire [0:0] CLBLL_R_X73Y108_SLICE_X111Y108_D_XOR;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_A;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_A1;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_A2;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_A3;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_A4;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_A5;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_A6;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_AO5;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_AO6;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_AQ;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_A_CY;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_A_XOR;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_B;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_B1;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_B2;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_B3;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_B4;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_B5;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_B6;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_BO5;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_BO6;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_B_CY;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_B_XOR;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_C;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_C1;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_C2;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_C3;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_C4;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_C5;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_C6;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_CLK;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_CO5;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_CO6;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_C_CY;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_C_XOR;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_D;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_D1;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_D2;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_D3;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_D4;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_D5;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_D6;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_DO5;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_DO6;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_D_CY;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_D_XOR;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X110Y109_SR;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_A;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_A1;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_A2;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_A3;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_A4;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_A5;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_A6;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_AO5;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_AO6;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_A_CY;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_A_XOR;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_B;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_B1;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_B2;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_B3;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_B4;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_B5;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_B6;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_BO5;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_BO6;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_B_CY;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_B_XOR;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_C;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_C1;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_C2;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_C3;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_C4;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_C5;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_C6;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_CO5;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_CO6;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_C_CY;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_C_XOR;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_D;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_D1;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_D2;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_D3;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_D4;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_D5;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_D6;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_DO5;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_DO6;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_D_CY;
  wire [0:0] CLBLL_R_X73Y109_SLICE_X111Y109_D_XOR;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_A;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_A1;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_A2;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_A3;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_A4;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_A5;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_A5Q;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_A6;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_AMUX;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_AO5;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_AO6;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_AQ;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_AX;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_A_CY;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_A_XOR;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_B;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_B1;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_B2;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_B3;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_B4;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_B5;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_B6;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_BO5;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_BO6;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_B_CY;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_B_XOR;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_C;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_C1;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_C2;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_C3;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_C4;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_C5;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_C6;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_CLK;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_CO5;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_CO6;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_C_CY;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_C_XOR;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_D;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_D1;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_D2;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_D3;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_D4;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_D5;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_D6;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_DO5;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_DO6;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_D_CY;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_D_XOR;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X110Y111_SR;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_A;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_A1;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_A2;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_A3;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_A4;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_A5;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_A6;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_AO5;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_AO6;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_A_CY;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_A_XOR;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_B;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_B1;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_B2;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_B3;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_B4;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_B5;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_B6;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_BO5;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_BO6;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_B_CY;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_B_XOR;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_C;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_C1;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_C2;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_C3;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_C4;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_C5;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_C6;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_CO5;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_CO6;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_C_CY;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_C_XOR;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_D;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_D1;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_D2;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_D3;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_D4;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_D5;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_D6;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_DO5;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_DO6;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_D_CY;
  wire [0:0] CLBLL_R_X73Y111_SLICE_X111Y111_D_XOR;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_A;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_A1;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_A2;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_A3;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_A4;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_A5;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_A5Q;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_A6;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_AMUX;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_AO5;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_AO6;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_AQ;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_AX;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_A_CY;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_A_XOR;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_B;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_B1;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_B2;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_B3;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_B4;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_B5;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_B6;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_BO5;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_BO6;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_B_CY;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_B_XOR;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_C;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_C1;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_C2;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_C3;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_C4;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_C5;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_C6;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_CLK;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_CO5;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_CO6;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_C_CY;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_C_XOR;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_D;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_D1;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_D2;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_D3;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_D4;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_D5;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_D6;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_DO5;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_DO6;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_D_CY;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_D_XOR;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X110Y113_SR;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_A;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_A1;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_A2;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_A3;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_A4;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_A5;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_A6;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_AO5;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_AO6;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_A_CY;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_A_XOR;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_B;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_B1;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_B2;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_B3;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_B4;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_B5;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_B6;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_BO5;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_BO6;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_B_CY;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_B_XOR;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_C;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_C1;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_C2;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_C3;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_C4;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_C5;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_C6;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_CO5;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_CO6;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_C_CY;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_C_XOR;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_D;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_D1;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_D2;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_D3;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_D4;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_D5;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_D6;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_DO5;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_DO6;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_D_CY;
  wire [0:0] CLBLL_R_X73Y113_SLICE_X111Y113_D_XOR;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_A;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_A1;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_A2;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_A3;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_A4;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_A5;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_A6;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_AO5;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_AO6;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_AQ;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_A_CY;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_A_XOR;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_B;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_B1;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_B2;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_B3;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_B4;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_B5;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_B5Q;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_B6;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_BMUX;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_BO5;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_BO6;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_BQ;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_B_CY;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_B_XOR;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_C;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_C1;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_C2;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_C3;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_C4;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_C5;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_C6;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_CLK;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_CO5;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_CO6;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_C_CY;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_C_XOR;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_D;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_D1;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_D2;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_D3;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_D4;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_D5;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_D6;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_DO5;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_DO6;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_D_CY;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_D_XOR;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_SR;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_A;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_A1;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_A2;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_A3;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_A4;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_A5;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_A5Q;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_A6;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_AMUX;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_AO5;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_AO6;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_AQ;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_A_CY;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_A_XOR;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_B;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_B1;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_B2;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_B3;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_B4;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_B5;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_B6;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_BO5;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_BO6;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_BQ;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_BX;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_B_CY;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_B_XOR;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_C;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_C1;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_C2;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_C3;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_C4;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_C5;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_C6;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_CLK;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_CO5;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_CO6;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_C_CY;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_C_XOR;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_D;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_D1;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_D2;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_D3;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_D4;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_D5;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_D6;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_DO5;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_DO6;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_D_CY;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_D_XOR;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_SR;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_A;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_A1;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_A2;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_A3;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_A4;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_A5;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_A5Q;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_A6;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_AMUX;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_AO5;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_AO6;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_AQ;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_AX;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_A_CY;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_A_XOR;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_B;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_B1;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_B2;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_B3;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_B4;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_B5;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_B5Q;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_B6;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_BMUX;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_BO5;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_BO6;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_BQ;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_B_CY;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_B_XOR;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_C;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_C1;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_C2;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_C3;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_C4;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_C5;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_C6;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_CLK;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_CMUX;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_CO5;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_CO6;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_C_CY;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_C_XOR;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_D;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_D1;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_D2;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_D3;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_D4;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_D5;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_D6;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_DO5;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_DO6;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_D_CY;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_D_XOR;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_SR;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_A;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_A1;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_A2;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_A3;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_A4;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_A5;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_A6;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_AO5;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_AO6;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_AQ;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_AX;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_A_CY;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_A_XOR;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_B;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_B1;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_B2;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_B3;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_B4;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_B5;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_B6;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_BO5;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_BO6;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_B_CY;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_B_XOR;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_C;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_C1;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_C2;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_C3;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_C4;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_C5;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_C6;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_CLK;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_CO5;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_CO6;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_C_CY;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_C_XOR;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_D;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_D1;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_D2;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_D3;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_D4;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_D5;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_D6;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_DO5;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_D_CY;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_D_XOR;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_SR;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_A;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_A1;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_A2;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_A3;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_A4;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_A5;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_A6;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_AO5;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_AO6;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_AQ;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_A_CY;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_A_XOR;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_B;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_B1;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_B2;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_B3;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_B4;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_B5;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_B6;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_BO5;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_BO6;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_BQ;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_B_CY;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_B_XOR;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_C;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_C1;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_C2;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_C3;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_C4;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_C5;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_C6;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_CLK;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_CO5;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_CO6;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_C_CY;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_C_XOR;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_D;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_D1;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_D2;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_D3;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_D4;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_D5;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_D6;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_DO5;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_DO6;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_D_CY;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_D_XOR;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_SR;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_A;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_A1;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_A2;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_A3;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_A4;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_A5;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_A6;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_AO5;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_AO6;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_AQ;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_A_CY;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_A_XOR;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_B;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_B1;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_B2;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_B3;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_B4;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_B5;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_B6;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_BO5;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_BO6;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_BQ;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_B_CY;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_B_XOR;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_C;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_C1;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_C2;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_C3;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_C4;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_C5;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_C6;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_CLK;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_CO5;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_CO6;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_C_CY;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_C_XOR;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_D;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_D1;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_D2;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_D3;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_D4;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_D5;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_D6;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_DO5;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_DO6;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_D_CY;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_D_XOR;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_SR;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_A;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_A1;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_A2;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_A3;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_A4;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_A5;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_A6;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_AMUX;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_AO5;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_AO6;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_A_CY;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_A_XOR;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_B;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_B1;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_B2;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_B3;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_B4;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_B5;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_B6;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_BO5;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_BO6;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_BQ;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_B_CY;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_B_XOR;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_C;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_C1;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_C2;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_C3;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_C4;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_C5;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_C6;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_CLK;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_CO5;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_CO6;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_CQ;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_C_CY;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_C_XOR;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_D;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_D1;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_D2;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_D3;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_D4;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_D5;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_D6;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_DMUX;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_DO5;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_DO6;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_D_CY;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_D_XOR;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_SR;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_A;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_A1;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_A2;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_A3;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_A4;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_A5;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_A6;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_AO5;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_AO6;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_AQ;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_A_CY;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_A_XOR;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_B;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_B1;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_B2;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_B3;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_B4;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_B5;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_B6;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_BO5;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_BO6;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_BQ;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_B_CY;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_B_XOR;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_C;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_C1;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_C2;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_C3;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_C4;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_C5;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_C6;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_CLK;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_CO5;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_CO6;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_CQ;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_C_CY;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_C_XOR;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_D;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_D1;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_D2;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_D3;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_D4;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_D5;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_D6;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_DO5;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_DO6;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_DQ;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_D_CY;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_D_XOR;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_SR;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_A;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_A1;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_A2;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_A3;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_A4;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_A5;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_A6;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_AO5;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_AO6;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_AQ;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_AX;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_A_CY;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_A_XOR;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_B;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_B1;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_B2;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_B3;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_B4;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_B5;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_B6;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_BO5;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_BO6;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_BQ;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_BX;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_B_CY;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_B_XOR;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_C;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_C1;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_C2;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_C3;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_C4;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_C5;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_C6;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_CE;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_CLK;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_CO5;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_CO6;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_CQ;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_CX;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_C_CY;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_C_XOR;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_D;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_D1;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_D2;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_D3;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_D4;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_D5;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_D6;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_DO5;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_DO6;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_D_CY;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_D_XOR;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_SR;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_A;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_A1;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_A2;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_A3;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_A4;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_A5;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_A6;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_AMUX;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_AO5;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_AO6;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_AQ;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_A_CY;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_A_XOR;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_B;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_B1;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_B2;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_B3;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_B4;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_B5;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_B6;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_BO5;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_BO6;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_BQ;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_B_CY;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_B_XOR;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_C;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_C1;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_C2;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_C3;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_C4;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_C5;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_C6;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_CLK;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_CO5;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_CO6;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_CQ;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_C_CY;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_C_XOR;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_D;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_D1;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_D2;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_D3;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_D4;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_D5;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_D6;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_DO5;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_DO6;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_DQ;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_D_CY;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_D_XOR;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_SR;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_A;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_A1;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_A2;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_A3;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_A4;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_A5;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_A5Q;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_A6;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_AMUX;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_AO5;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_AO6;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_AQ;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_AX;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_A_CY;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_A_XOR;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_B;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_B1;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_B2;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_B3;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_B4;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_B5;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_B6;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_BO5;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_BO6;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_BQ;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_B_CY;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_B_XOR;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_C;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_C1;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_C2;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_C3;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_C4;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_C5;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_C6;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_CLK;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_CMUX;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_CO5;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_CO6;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_C_CY;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_C_XOR;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_D;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_D1;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_D2;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_D3;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_D4;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_D5;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_D6;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_DO5;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_DO6;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_D_CY;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_D_XOR;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_SR;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_A;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_A1;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_A2;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_A3;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_A4;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_A5;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_A6;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_AO5;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_AO6;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_AQ;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_A_CY;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_A_XOR;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_B;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_B1;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_B2;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_B3;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_B4;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_B5;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_B6;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_BO5;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_BO6;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_BQ;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_B_CY;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_B_XOR;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_C;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_C1;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_C2;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_C3;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_C4;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_C5;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_C6;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_CLK;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_CO5;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_CO6;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_C_CY;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_C_XOR;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_D;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_D1;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_D2;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_D3;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_D4;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_D5;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_D6;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_DO5;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_DO6;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_D_CY;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_D_XOR;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_SR;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_A;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_A1;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_A2;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_A3;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_A4;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_A5;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_A6;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_AO5;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_AO6;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_AQ;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_AX;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_A_CY;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_A_XOR;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_B;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_B1;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_B2;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_B3;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_B4;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_B5;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_B6;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_BMUX;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_BO5;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_BO6;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_B_CY;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_B_XOR;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_C;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_C1;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_C2;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_C3;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_C4;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_C5;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_C6;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_CE;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_CLK;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_CO5;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_CO6;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_C_CY;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_C_XOR;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_D;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_D1;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_D2;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_D3;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_D4;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_D5;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_D6;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_DO5;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_DO6;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_D_CY;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_D_XOR;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_SR;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_A;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_A1;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_A2;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_A3;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_A4;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_A5;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_A5Q;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_A6;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_AMUX;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_AO5;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_AO6;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_AQ;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_A_CY;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_A_XOR;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_B;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_B1;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_B2;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_B3;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_B4;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_B5;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_B6;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_BO5;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_BO6;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_BQ;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_B_CY;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_B_XOR;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_C;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_C1;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_C2;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_C3;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_C4;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_C5;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_C6;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_CLK;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_CO5;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_CO6;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_CQ;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_C_CY;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_C_XOR;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_D;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_D1;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_D2;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_D3;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_D4;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_D5;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_D6;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_DO5;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_DO6;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_DQ;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_D_CY;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_D_XOR;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_SR;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_A;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_A1;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_A2;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_A3;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_A4;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_A5;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_A5Q;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_A6;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_AMUX;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_AO5;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_AO6;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_AQ;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_AX;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_A_CY;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_A_XOR;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_B;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_B1;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_B2;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_B3;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_B4;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_B5;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_B6;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_BO5;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_BO6;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_BQ;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_B_CY;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_B_XOR;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_C;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_C1;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_C2;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_C3;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_C4;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_C5;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_C6;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_CLK;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_CMUX;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_CO5;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_CO6;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_C_CY;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_C_XOR;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_D;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_D1;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_D2;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_D3;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_D4;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_D5;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_D6;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_DO5;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_DO6;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_DQ;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_D_CY;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_D_XOR;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_SR;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_A;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_A1;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_A2;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_A3;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_A4;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_A5;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_A6;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_AO5;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_AO6;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_AQ;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_A_CY;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_A_XOR;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_B;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_B1;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_B2;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_B3;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_B4;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_B5;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_B6;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_BMUX;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_BO5;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_BO6;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_B_CY;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_B_XOR;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_C;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_C1;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_C2;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_C3;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_C4;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_C5;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_C6;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_CLK;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_CO5;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_CO6;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_CQ;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_C_CY;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_C_XOR;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_D;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_D1;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_D2;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_D3;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_D4;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_D5;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_D6;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_DO5;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_DO6;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_DQ;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_D_CY;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_D_XOR;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_SR;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_A;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_A1;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_A2;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_A3;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_A4;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_A5;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_A5Q;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_A6;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_AMUX;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_AO5;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_AO6;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_AQ;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_AX;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_A_CY;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_A_XOR;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_B;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_B1;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_B2;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_B3;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_B4;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_B5;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_B6;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_BO5;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_BO6;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_BQ;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_B_CY;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_B_XOR;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_C;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_C1;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_C2;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_C3;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_C4;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_C5;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_C6;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_CLK;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_CMUX;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_CO5;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_CO6;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_C_CY;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_C_XOR;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_D;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_D1;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_D2;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_D3;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_D4;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_D5;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_D6;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_DO5;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_DO6;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_DQ;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_D_CY;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_D_XOR;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_SR;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_A;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_A1;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_A2;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_A3;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_A4;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_A5;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_A6;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_AO5;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_AO6;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_AQ;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_A_CY;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_A_XOR;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_B;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_B1;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_B2;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_B3;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_B4;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_B5;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_B6;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_BMUX;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_BO5;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_BO6;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_B_CY;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_B_XOR;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_C;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_C1;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_C2;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_C3;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_C4;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_C5;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_C6;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_CLK;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_CO5;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_CO6;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_CQ;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_C_CY;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_C_XOR;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_D;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_D1;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_D2;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_D3;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_D4;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_D5;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_D6;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_DO5;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_DO6;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_D_CY;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_D_XOR;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_SR;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_A;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_A1;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_A2;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_A3;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_A4;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_A5;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_A6;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_AO5;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_AO6;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_AQ;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_A_CY;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_A_XOR;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_B;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_B1;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_B2;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_B3;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_B4;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_B5;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_B6;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_BO5;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_BO6;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_B_CY;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_B_XOR;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_C;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_C1;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_C2;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_C3;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_C4;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_C5;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_C6;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_CLK;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_CO5;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_CO6;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_C_CY;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_C_XOR;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_D;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_D1;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_D2;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_D3;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_D4;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_D5;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_D6;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_DO5;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_DO6;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_D_CY;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_D_XOR;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_SR;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_A;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_A1;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_A2;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_A3;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_A4;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_A5;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_A6;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_AO5;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_AO6;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_AQ;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_A_CY;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_A_XOR;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_B;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_B1;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_B2;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_B3;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_B4;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_B5;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_B6;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_BO5;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_BO6;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_BQ;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_B_CY;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_B_XOR;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_C;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_C1;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_C2;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_C3;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_C4;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_C5;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_C6;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_CLK;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_CO5;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_CO6;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_C_CY;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_C_XOR;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_D;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_D1;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_D2;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_D3;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_D4;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_D5;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_D6;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_DO5;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_DO6;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_D_CY;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_D_XOR;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_SR;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_A;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_A1;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_A2;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_A3;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_A4;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_A5;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_A6;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_AO5;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_AO6;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_AQ;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_AX;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_A_CY;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_A_XOR;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_B;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_B1;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_B2;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_B3;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_B4;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_B5;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_B6;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_BO5;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_BO6;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_B_CY;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_B_XOR;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_C;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_C1;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_C2;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_C3;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_C4;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_C5;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_C6;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_CLK;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_CO5;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_CO6;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_C_CY;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_C_XOR;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_D;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_D1;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_D2;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_D3;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_D4;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_D5;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_D6;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_DO5;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_DO6;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_D_CY;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_D_XOR;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X110Y131_SR;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_A;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_A1;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_A2;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_A3;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_A4;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_A5;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_A6;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_AO5;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_AO6;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_AQ;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_A_CY;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_A_XOR;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_B;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_B1;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_B2;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_B3;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_B4;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_B5;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_B6;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_BO5;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_BO6;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_B_CY;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_B_XOR;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_C;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_C1;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_C2;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_C3;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_C4;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_C5;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_C6;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_CLK;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_CO5;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_CO6;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_C_CY;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_C_XOR;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_D;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_D1;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_D2;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_D3;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_D4;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_D5;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_D6;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_DO5;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_DO6;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_D_CY;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_D_XOR;
  wire [0:0] CLBLL_R_X73Y131_SLICE_X111Y131_SR;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_A;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_A1;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_A2;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_A3;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_A4;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_A5;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_A6;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_AMUX;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_AO5;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_AO6;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_A_CY;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_A_XOR;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_B;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_B1;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_B2;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_B3;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_B4;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_B5;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_B6;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_BO5;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_BO6;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_B_CY;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_B_XOR;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_C;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_C1;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_C2;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_C3;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_C4;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_C5;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_C6;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_CO5;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_CO6;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_C_CY;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_C_XOR;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_D;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_D1;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_D2;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_D3;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_D4;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_D5;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_D6;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_DO5;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_DO6;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_D_CY;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X110Y132_D_XOR;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_A;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_A1;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_A2;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_A3;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_A4;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_A5;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_A6;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_AMUX;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_AO5;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_AO6;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_A_CY;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_A_XOR;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_B;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_B1;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_B2;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_B3;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_B4;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_B5;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_B6;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_BO5;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_BO6;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_B_CY;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_B_XOR;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_C;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_C1;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_C2;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_C3;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_C4;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_C5;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_C6;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_CMUX;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_CO5;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_CO6;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_C_CY;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_C_XOR;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_D;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_D1;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_D2;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_D3;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_D4;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_D5;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_D6;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_DO5;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_DO6;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_D_CY;
  wire [0:0] CLBLL_R_X73Y132_SLICE_X111Y132_D_XOR;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_A;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_A1;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_A2;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_A3;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_A4;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_A5;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_A5Q;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_A6;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_AMUX;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_AO5;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_AO6;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_AQ;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_A_CY;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_A_XOR;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_B;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_B1;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_B2;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_B3;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_B4;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_B5;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_B6;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_BO5;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_BO6;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_BQ;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_B_CY;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_B_XOR;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_C;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_C1;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_C2;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_C3;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_C4;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_C5;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_C6;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_CLK;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_CO5;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_CO6;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_CQ;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_C_CY;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_C_XOR;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_D;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_D1;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_D2;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_D3;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_D4;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_D5;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_D6;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_DO5;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_DO6;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_D_CY;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_D_XOR;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X110Y133_SR;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_A;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_A1;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_A2;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_A3;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_A4;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_A5;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_A5Q;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_A6;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_AMUX;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_AO5;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_AO6;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_AQ;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_AX;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_A_CY;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_A_XOR;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_B;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_B1;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_B2;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_B3;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_B4;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_B5;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_B6;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_BMUX;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_BO5;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_BO6;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_B_CY;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_B_XOR;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_C;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_C1;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_C2;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_C3;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_C4;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_C5;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_C6;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_CLK;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_CO5;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_CO6;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_C_CY;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_C_XOR;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_D;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_D1;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_D2;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_D3;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_D4;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_D5;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_D6;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_DO5;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_DO6;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_D_CY;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_D_XOR;
  wire [0:0] CLBLL_R_X73Y133_SLICE_X111Y133_SR;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_A;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_A1;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_A2;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_A3;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_A4;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_A5;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_A6;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_AMUX;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_AO5;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_AO6;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_A_CY;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_A_XOR;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_B;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_B1;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_B2;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_B3;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_B4;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_B5;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_B6;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_BO5;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_BO6;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_B_CY;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_B_XOR;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_C;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_C1;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_C2;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_C3;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_C4;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_C5;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_C6;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_CO5;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_CO6;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_C_CY;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_C_XOR;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_D;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_D1;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_D2;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_D3;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_D4;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_D5;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_D6;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_DO5;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_DO6;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_D_CY;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X110Y134_D_XOR;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_A;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_A1;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_A2;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_A3;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_A4;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_A5;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_A6;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_AO5;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_AO6;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_AQ;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_A_CY;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_A_XOR;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_B;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_B1;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_B2;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_B3;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_B4;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_B5;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_B6;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_BO5;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_BO6;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_B_CY;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_B_XOR;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_C;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_C1;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_C2;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_C3;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_C4;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_C5;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_C6;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_CLK;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_CO5;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_CO6;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_C_CY;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_C_XOR;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_D;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_D1;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_D2;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_D3;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_D4;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_D5;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_D6;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_DO5;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_DO6;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_D_CY;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_D_XOR;
  wire [0:0] CLBLL_R_X73Y134_SLICE_X111Y134_SR;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_A;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_A1;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_A2;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_A3;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_A4;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_A5;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_A6;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_AO5;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_AO6;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_A_CY;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_A_XOR;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_B;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_B1;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_B2;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_B3;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_B4;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_B5;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_B6;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_BO5;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_BO6;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_B_CY;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_B_XOR;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_C;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_C1;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_C2;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_C3;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_C4;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_C5;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_C6;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_CO5;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_CO6;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_C_CY;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_C_XOR;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_D;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_D1;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_D2;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_D3;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_D4;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_D5;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_D6;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_DO5;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_DO6;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_D_CY;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X114Y103_D_XOR;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_A;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_A1;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_A2;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_A3;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_A4;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_A5;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_A6;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_AO5;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_AO6;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_AQ;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_A_CY;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_A_XOR;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_B;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_B1;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_B2;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_B3;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_B4;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_B5;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_B6;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_BO5;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_BO6;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_B_CY;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_B_XOR;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_C;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_C1;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_C2;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_C3;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_C4;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_C5;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_C6;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_CLK;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_CO5;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_CO6;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_C_CY;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_C_XOR;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_D;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_D1;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_D2;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_D3;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_D4;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_D5;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_D6;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_DO5;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_DO6;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_D_CY;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_D_XOR;
  wire [0:0] CLBLL_R_X75Y103_SLICE_X115Y103_SR;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_A;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_A1;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_A2;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_A3;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_A4;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_A5;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_A6;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_AO5;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_AO6;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_AQ;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_AX;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_A_CY;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_A_XOR;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_B;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_B1;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_B2;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_B3;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_B4;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_B5;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_B6;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_BO5;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_BO6;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_B_CY;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_B_XOR;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_C;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_C1;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_C2;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_C3;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_C4;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_C5;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_C6;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_CLK;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_CO5;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_CO6;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_C_CY;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_C_XOR;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_D;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_D1;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_D2;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_D3;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_D4;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_D5;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_D6;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_DO5;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_DO6;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_D_CY;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_D_XOR;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X114Y107_SR;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_A;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_A1;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_A2;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_A3;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_A4;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_A5;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_A6;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_AO5;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_AO6;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_A_CY;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_A_XOR;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_B;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_B1;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_B2;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_B3;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_B4;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_B5;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_B6;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_BO5;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_BO6;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_B_CY;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_B_XOR;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_C;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_C1;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_C2;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_C3;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_C4;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_C5;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_C6;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_CO5;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_CO6;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_C_CY;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_C_XOR;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_D;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_D1;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_D2;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_D3;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_D4;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_D5;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_D6;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_DO5;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_DO6;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_D_CY;
  wire [0:0] CLBLL_R_X75Y107_SLICE_X115Y107_D_XOR;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_A;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_A1;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_A2;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_A3;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_A4;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_A5;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_A6;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_AO5;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_AO6;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_AQ;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_AX;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_A_CY;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_A_XOR;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_B;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_B1;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_B2;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_B3;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_B4;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_B5;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_B6;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_BO5;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_BO6;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_B_CY;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_B_XOR;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_C;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_C1;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_C2;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_C3;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_C4;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_C5;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_C6;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_CLK;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_CO5;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_CO6;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_C_CY;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_C_XOR;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_D;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_D1;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_D2;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_D3;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_D4;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_D5;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_D6;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_DO5;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_DO6;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_D_CY;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_D_XOR;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X114Y113_SR;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_A;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_A1;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_A2;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_A3;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_A4;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_A5;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_A6;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_AO5;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_AO6;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_A_CY;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_A_XOR;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_B;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_B1;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_B2;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_B3;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_B4;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_B5;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_B6;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_BO5;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_BO6;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_B_CY;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_B_XOR;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_C;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_C1;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_C2;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_C3;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_C4;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_C5;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_C6;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_CO5;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_CO6;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_C_CY;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_C_XOR;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_D;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_D1;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_D2;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_D3;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_D4;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_D5;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_D6;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_DO5;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_DO6;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_D_CY;
  wire [0:0] CLBLL_R_X75Y113_SLICE_X115Y113_D_XOR;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_A;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_A1;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_A2;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_A3;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_A4;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_A5;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_A6;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_AMUX;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_AO5;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_AO6;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_AQ;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_A_CY;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_A_XOR;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_B;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_B1;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_B2;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_B3;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_B4;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_B5;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_B6;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_BO5;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_BO6;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_BQ;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_B_CY;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_B_XOR;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_C;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_C1;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_C2;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_C3;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_C4;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_C5;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_C6;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_CLK;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_CO5;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_CO6;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_C_CY;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_C_XOR;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_D;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_D1;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_D2;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_D3;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_D4;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_D5;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_D6;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_DO5;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_DO6;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_D_CY;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_D_XOR;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X114Y121_SR;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_A;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_A1;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_A2;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_A3;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_A4;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_A5;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_A6;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_AO5;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_AO6;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_A_CY;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_A_XOR;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_B;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_B1;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_B2;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_B3;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_B4;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_B5;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_B6;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_BO5;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_BO6;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_B_CY;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_B_XOR;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_C;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_C1;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_C2;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_C3;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_C4;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_C5;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_C6;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_CO5;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_CO6;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_C_CY;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_C_XOR;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_D;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_D1;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_D2;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_D3;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_D4;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_D5;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_D6;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_DO5;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_DO6;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_D_CY;
  wire [0:0] CLBLL_R_X75Y121_SLICE_X115Y121_D_XOR;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_A;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_A1;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_A2;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_A3;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_A4;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_A5;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_A6;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_AO5;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_AO6;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_AQ;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_A_CY;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_A_XOR;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_B;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_B1;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_B2;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_B3;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_B4;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_B5;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_B6;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_BO5;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_BO6;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_BQ;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_B_CY;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_B_XOR;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_C;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_C1;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_C2;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_C3;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_C4;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_C5;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_C6;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_CLK;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_CO5;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_CO6;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_CQ;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_C_CY;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_C_XOR;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_D;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_D1;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_D2;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_D3;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_D4;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_D5;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_D6;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_DO5;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_DO6;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_D_CY;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_D_XOR;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X114Y122_SR;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_A;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_A1;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_A2;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_A3;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_A4;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_A5;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_A5Q;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_A6;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_AMUX;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_AO5;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_AO6;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_AQ;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_A_CY;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_A_XOR;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_B;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_B1;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_B2;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_B3;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_B4;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_B5;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_B6;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_BO5;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_BO6;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_BQ;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_B_CY;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_B_XOR;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_C;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_C1;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_C2;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_C3;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_C4;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_C5;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_C6;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_CLK;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_CO5;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_CO6;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_C_CY;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_C_XOR;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_D;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_D1;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_D2;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_D3;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_D4;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_D5;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_D6;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_DO5;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_DO6;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_D_CY;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_D_XOR;
  wire [0:0] CLBLL_R_X75Y122_SLICE_X115Y122_SR;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_A;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_A1;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_A2;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_A3;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_A4;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_A5;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_A6;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_AMUX;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_AO5;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_AO6;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_A_CY;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_A_XOR;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_B;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_B1;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_B2;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_B3;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_B4;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_B5;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_B6;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_BO5;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_BO6;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_BQ;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_B_CY;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_B_XOR;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_C;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_C1;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_C2;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_C3;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_C4;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_C5;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_C6;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_CLK;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_CO5;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_CO6;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_C_CY;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_C_XOR;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_D;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_D1;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_D2;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_D3;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_D4;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_D5;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_D6;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_DO5;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_DO6;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_D_CY;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_D_XOR;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_SR;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_A;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_A1;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_A2;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_A3;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_A4;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_A5;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_A6;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_AMUX;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_AO5;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_AO6;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_AQ;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_AX;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_A_CY;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_A_XOR;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_B;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_B1;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_B2;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_B3;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_B4;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_B5;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_B6;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_BO5;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_BO6;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_B_CY;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_B_XOR;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_C;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_C1;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_C2;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_C3;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_C4;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_C5;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_C6;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_CE;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_CLK;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_CO5;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_CO6;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_C_CY;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_C_XOR;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_D;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_D1;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_D2;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_D3;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_D4;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_D5;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_D6;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_DO5;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_DO6;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_D_CY;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_D_XOR;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_SR;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_A;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_A1;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_A2;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_A3;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_A4;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_A5;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_A6;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_AO5;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_AO6;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_AQ;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_A_CY;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_A_XOR;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_B;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_B1;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_B2;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_B3;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_B4;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_B5;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_B6;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_BO5;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_BO6;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_BQ;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_B_CY;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_B_XOR;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_C;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_C1;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_C2;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_C3;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_C4;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_C5;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_C5Q;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_C6;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_CLK;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_CMUX;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_CO5;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_CO6;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_CQ;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_C_CY;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_C_XOR;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_D;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_D1;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_D2;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_D3;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_D4;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_D5;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_D5Q;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_D6;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_DMUX;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_DO5;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_DO6;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_DQ;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_D_CY;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_D_XOR;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_SR;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_A;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_A1;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_A2;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_A3;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_A4;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_A5;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_A6;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_AO5;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_AO6;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_AQ;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_A_CY;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_A_XOR;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_B;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_B1;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_B2;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_B3;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_B4;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_B5;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_B5Q;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_B6;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_BMUX;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_BO5;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_BO6;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_BQ;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_B_CY;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_B_XOR;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_C;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_C1;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_C2;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_C3;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_C4;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_C5;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_C6;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_CLK;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_CO5;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_CO6;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_CQ;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_C_CY;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_C_XOR;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_D;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_D1;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_D2;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_D3;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_D4;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_D5;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_D6;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_DO5;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_DO6;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_DQ;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_D_CY;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_D_XOR;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_SR;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_A;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_A1;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_A2;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_A3;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_A4;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_A5;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_A5Q;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_A6;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_AMUX;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_AO5;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_AO6;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_AQ;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_A_CY;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_A_XOR;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_B;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_B1;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_B2;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_B3;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_B4;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_B5;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_B6;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_BO5;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_BO6;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_BQ;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_B_CY;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_B_XOR;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_C;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_C1;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_C2;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_C3;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_C4;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_C5;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_C6;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_CLK;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_CMUX;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_CO5;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_CO6;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_C_CY;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_C_XOR;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_D;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_D1;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_D2;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_D3;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_D4;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_D5;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_D6;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_DO5;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_DO6;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_DQ;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_D_CY;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_D_XOR;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_SR;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_A;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_A1;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_A2;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_A3;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_A4;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_A5;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_A6;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_AO5;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_AO6;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_AQ;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_A_CY;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_A_XOR;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_B;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_B1;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_B2;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_B3;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_B4;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_B5;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_B6;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_BO5;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_BO6;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_BQ;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_B_CY;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_B_XOR;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_C;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_C1;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_C2;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_C3;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_C4;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_C5;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_C6;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_CLK;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_CO5;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_CO6;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_CQ;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_C_CY;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_C_XOR;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_D;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_D1;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_D2;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_D3;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_D4;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_D5;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_D6;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_DO5;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_DO6;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_DQ;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_D_CY;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_D_XOR;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_SR;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_A;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_A1;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_A2;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_A3;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_A4;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_A5;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_A6;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_AMUX;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_AO5;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_AO6;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_A_CY;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_A_XOR;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_B;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_B1;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_B2;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_B3;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_B4;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_B5;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_B6;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_BMUX;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_BO5;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_BO6;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_B_CY;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_B_XOR;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_C;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_C1;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_C2;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_C3;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_C4;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_C5;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_C6;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_CLK;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_CO5;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_CO6;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_CQ;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_C_CY;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_C_XOR;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_D;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_D1;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_D2;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_D3;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_D4;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_D5;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_D6;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_DMUX;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_DO5;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_DO6;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_D_CY;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_D_XOR;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_SR;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_A;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_A1;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_A2;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_A3;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_A4;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_A5;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_A6;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_AO5;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_AO6;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_A_CY;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_A_XOR;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_B;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_B1;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_B2;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_B3;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_B4;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_B5;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_B6;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_BO5;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_BO6;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_B_CY;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_B_XOR;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_C;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_C1;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_C2;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_C3;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_C4;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_C5;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_C6;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_CO5;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_CO6;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_C_CY;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_C_XOR;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_D;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_D1;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_D2;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_D3;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_D4;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_D5;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_D6;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_DO5;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_DO6;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_D_CY;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_D_XOR;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_A;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_A1;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_A2;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_A3;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_A4;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_A5;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_A6;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_AO5;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_AO6;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_AQ;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_A_CY;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_A_XOR;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_B;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_B1;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_B2;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_B3;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_B4;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_B5;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_B6;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_BO5;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_BO6;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_BQ;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_B_CY;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_B_XOR;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_C;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_C1;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_C2;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_C3;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_C4;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_C5;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_C6;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_CLK;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_CMUX;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_CO5;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_CO6;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_C_CY;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_C_XOR;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_D;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_D1;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_D2;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_D3;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_D4;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_D5;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_D6;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_DO5;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_DO6;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_DQ;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_D_CY;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_D_XOR;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X114Y129_SR;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_A;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_A1;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_A2;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_A3;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_A4;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_A5;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_A6;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_AO5;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_AO6;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_AQ;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_A_CY;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_A_XOR;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_B;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_B1;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_B2;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_B3;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_B4;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_B5;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_B6;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_BO5;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_BO6;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_B_CY;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_B_XOR;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_C;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_C1;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_C2;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_C3;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_C4;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_C5;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_C6;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_CLK;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_CO5;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_CO6;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_C_CY;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_C_XOR;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_D;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_D1;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_D2;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_D3;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_D4;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_D5;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_D6;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_DO5;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_DO6;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_D_CY;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_D_XOR;
  wire [0:0] CLBLL_R_X75Y129_SLICE_X115Y129_SR;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_A;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_A1;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_A2;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_A3;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_A4;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_A5;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_A6;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_AO5;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_AO6;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_AQ;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_A_CY;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_A_XOR;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_B;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_B1;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_B2;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_B3;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_B4;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_B5;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_B6;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_BO5;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_BO6;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_B_CY;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_B_XOR;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_C;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_C1;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_C2;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_C3;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_C4;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_C5;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_C6;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_CLK;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_CO5;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_CO6;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_C_CY;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_C_XOR;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_D;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_D1;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_D2;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_D3;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_D4;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_D5;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_D6;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_DO5;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_DO6;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_D_CY;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_D_XOR;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X114Y130_SR;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_A;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_A1;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_A2;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_A3;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_A4;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_A5;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_A6;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_AO5;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_AO6;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_AQ;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_A_CY;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_A_XOR;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_B;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_B1;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_B2;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_B3;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_B4;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_B5;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_B6;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_BMUX;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_BO5;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_BO6;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_B_CY;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_B_XOR;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_C;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_C1;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_C2;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_C3;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_C4;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_C5;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_C6;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_CLK;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_CO5;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_CO6;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_CQ;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_C_CY;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_C_XOR;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_D;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_D1;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_D2;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_D3;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_D4;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_D5;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_D6;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_DO5;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_DO6;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_D_CY;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_D_XOR;
  wire [0:0] CLBLL_R_X75Y130_SLICE_X115Y130_SR;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_A;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_A1;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_A2;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_A3;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_A4;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_A5;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_A6;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_AO5;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_AO6;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_AQ;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_A_CY;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_A_XOR;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_B;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_B1;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_B2;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_B3;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_B4;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_B5;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_B6;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_BO5;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_BO6;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_BQ;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_B_CY;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_B_XOR;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_C;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_C1;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_C2;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_C3;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_C4;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_C5;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_C6;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_CLK;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_CMUX;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_CO5;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_CO6;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_C_CY;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_C_XOR;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_D;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_D1;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_D2;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_D3;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_D4;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_D5;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_D6;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_DO5;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_DO6;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_D_CY;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_D_XOR;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X114Y133_SR;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_A;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_A1;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_A2;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_A3;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_A4;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_A5;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_A6;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_AO5;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_AO6;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_AQ;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_A_CY;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_A_XOR;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_B;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_B1;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_B2;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_B3;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_B4;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_B5;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_B6;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_BO5;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_BO6;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_BQ;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_BX;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_B_CY;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_B_XOR;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_C;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_C1;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_C2;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_C3;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_C4;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_C5;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_C6;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_CLK;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_CO5;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_CO6;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_C_CY;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_C_XOR;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_D;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_D1;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_D2;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_D3;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_D4;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_D5;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_D6;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_DO5;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_DO6;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_D_CY;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_D_XOR;
  wire [0:0] CLBLL_R_X75Y133_SLICE_X115Y133_SR;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_A;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_A1;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_A2;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_A3;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_A4;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_A5;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_A5Q;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_A6;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_AMUX;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_AO5;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_AO6;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_AQ;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_AX;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_A_CY;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_A_XOR;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_B;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_B1;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_B2;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_B3;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_B4;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_B5;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_B6;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_BMUX;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_BO5;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_BO6;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_B_CY;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_B_XOR;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_C;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_C1;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_C2;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_C3;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_C4;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_C5;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_C6;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_CLK;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_CMUX;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_CO5;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_CO6;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_C_CY;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_C_XOR;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_D;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_D1;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_D2;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_D3;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_D4;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_D5;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_D6;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_DO5;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_DO6;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_D_CY;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_D_XOR;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X114Y134_SR;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_A;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_A1;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_A2;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_A3;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_A4;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_A5;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_A6;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_AMUX;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_AO5;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_AO6;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_AQ;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_AX;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_A_CY;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_A_XOR;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_B;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_B1;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_B2;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_B3;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_B4;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_B5;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_B6;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_BO5;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_BO6;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_B_CY;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_B_XOR;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_C;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_C1;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_C2;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_C3;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_C4;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_C5;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_C6;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_CLK;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_CO5;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_CO6;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_C_CY;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_C_XOR;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_D;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_D1;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_D2;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_D3;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_D4;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_D5;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_D6;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_DMUX;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_DO5;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_DO6;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_D_CY;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_D_XOR;
  wire [0:0] CLBLL_R_X75Y134_SLICE_X115Y134_SR;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_A;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_A1;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_A2;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_A3;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_A4;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_A5;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_A6;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_AO5;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_AO6;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_AQ;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_AX;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_A_CY;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_A_XOR;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_B;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_B1;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_B2;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_B3;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_B4;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_B5;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_B6;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_BO5;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_BO6;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_BQ;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_BX;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_B_CY;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_B_XOR;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_C;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_C1;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_C2;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_C3;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_C4;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_C5;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_C6;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_CE;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_CLK;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_CO5;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_CO6;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_CQ;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_CX;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_C_CY;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_C_XOR;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_D;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_D1;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_D2;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_D3;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_D4;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_D5;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_D6;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_DO5;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_DO6;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_D_CY;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_D_XOR;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X118Y104_SR;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_A;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_A1;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_A2;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_A3;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_A4;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_A5;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_A5Q;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_A6;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_AMUX;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_AO5;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_AO6;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_AQ;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_A_CY;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_A_XOR;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_B;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_B1;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_B2;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_B3;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_B4;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_B5;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_B6;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_BO5;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_BO6;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_B_CY;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_B_XOR;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_C;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_C1;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_C2;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_C3;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_C4;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_C5;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_C6;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_CLK;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_CO5;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_CO6;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_C_CY;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_C_XOR;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_D;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_D1;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_D2;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_D3;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_D4;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_D5;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_D6;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_DO5;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_DO6;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_D_CY;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_D_XOR;
  wire [0:0] CLBLL_R_X77Y104_SLICE_X119Y104_SR;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_A;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_A1;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_A2;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_A3;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_A4;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_A5;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_A6;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_AO5;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_AO6;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_AQ;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_AX;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_A_CY;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_A_XOR;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_B;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_B1;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_B2;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_B3;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_B4;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_B5;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_B6;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_BO5;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_BO6;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_B_CY;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_B_XOR;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_C;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_C1;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_C2;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_C3;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_C4;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_C5;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_C6;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_CLK;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_CO5;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_CO6;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_C_CY;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_C_XOR;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_D;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_D1;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_D2;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_D3;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_D4;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_D5;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_D6;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_DO5;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_DO6;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_D_CY;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_D_XOR;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X118Y108_SR;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_A;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_A1;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_A2;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_A3;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_A4;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_A5;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_A6;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_AO5;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_AO6;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_A_CY;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_A_XOR;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_B;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_B1;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_B2;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_B3;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_B4;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_B5;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_B6;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_BO5;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_BO6;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_B_CY;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_B_XOR;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_C;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_C1;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_C2;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_C3;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_C4;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_C5;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_C6;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_CO5;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_CO6;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_C_CY;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_C_XOR;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_D;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_D1;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_D2;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_D3;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_D4;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_D5;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_D6;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_DO5;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_DO6;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_D_CY;
  wire [0:0] CLBLL_R_X77Y108_SLICE_X119Y108_D_XOR;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_A;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_A1;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_A2;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_A3;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_A4;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_A5;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_A6;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_AO5;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_AO6;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_AQ;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_AX;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_A_CY;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_A_XOR;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_B;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_B1;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_B2;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_B3;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_B4;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_B5;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_B6;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_BO5;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_BO6;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_B_CY;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_B_XOR;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_C;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_C1;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_C2;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_C3;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_C4;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_C5;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_C6;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_CLK;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_CO5;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_CO6;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_C_CY;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_C_XOR;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_D;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_D1;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_D2;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_D3;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_D4;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_D5;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_D6;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_DO5;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_DO6;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_D_CY;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_D_XOR;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_SR;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_A;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_A1;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_A2;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_A3;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_A4;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_A5;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_A6;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_AO5;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_AO6;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_A_CY;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_A_XOR;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_B;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_B1;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_B2;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_B3;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_B4;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_B5;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_B6;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_BO5;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_BO6;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_B_CY;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_B_XOR;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_C;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_C1;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_C2;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_C3;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_C4;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_C5;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_C6;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_CO5;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_CO6;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_C_CY;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_C_XOR;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_D;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_D1;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_D2;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_D3;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_D4;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_D5;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_D6;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_DO5;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_DO6;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_D_CY;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_D_XOR;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_A;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_A1;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_A2;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_A3;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_A4;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_A5;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_A6;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_AO5;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_AO6;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_A_CY;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_A_XOR;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_B;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_B1;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_B2;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_B3;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_B4;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_B5;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_B6;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_BO5;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_BO6;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_B_CY;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_B_XOR;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_C;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_C1;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_C2;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_C3;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_C4;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_C5;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_C6;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_CO5;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_CO6;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_C_CY;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_C_XOR;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_D;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_D1;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_D2;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_D3;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_D4;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_D5;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_D6;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_DO5;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_DO6;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_D_CY;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X118Y121_D_XOR;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_A;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_A1;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_A2;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_A3;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_A4;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_A5;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_A6;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_AO5;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_AO6;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_AQ;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_A_CY;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_A_XOR;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_B;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_B1;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_B2;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_B3;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_B4;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_B5;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_B6;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_BMUX;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_BO5;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_BO6;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_B_CY;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_B_XOR;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_C;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_C1;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_C2;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_C3;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_C4;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_C5;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_C6;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_CLK;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_CO5;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_CO6;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_CQ;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_C_CY;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_C_XOR;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_D;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_D1;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_D2;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_D3;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_D4;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_D5;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_D6;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_DO5;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_DO6;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_DQ;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_D_CY;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_D_XOR;
  wire [0:0] CLBLL_R_X77Y121_SLICE_X119Y121_SR;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_A;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_A1;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_A2;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_A3;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_A4;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_A5;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_A6;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_AO5;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_AO6;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_AQ;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_A_CY;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_A_XOR;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_B;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_B1;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_B2;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_B3;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_B4;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_B5;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_B6;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_BO5;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_BO6;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_BQ;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_B_CY;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_B_XOR;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_C;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_C1;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_C2;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_C3;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_C4;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_C5;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_C6;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_CLK;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_CO5;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_C_CY;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_C_XOR;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_D;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_D1;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_D2;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_D3;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_D4;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_D5;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_D6;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_DO5;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_DO6;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_D_CY;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_D_XOR;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_SR;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_A;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_A1;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_A2;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_A3;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_A4;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_A5;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_A6;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_AMUX;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_AO5;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_AO6;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_A_CY;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_A_XOR;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_B;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_B1;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_B2;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_B3;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_B4;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_B5;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_B6;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_BO5;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_BO6;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_BQ;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_B_CY;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_B_XOR;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_C;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_C1;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_C2;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_C3;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_C4;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_C5;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_C6;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_CLK;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_CO5;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_CO6;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_CQ;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_C_CY;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_C_XOR;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_D;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_D1;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_D2;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_D3;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_D4;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_D5;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_D6;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_DO5;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_DO6;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_DQ;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_D_CY;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_D_XOR;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_SR;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_A;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_A1;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_A2;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_A3;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_A4;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_A5;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_A6;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_AO5;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_AO6;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_AQ;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_A_CY;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_A_XOR;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_B;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_B1;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_B2;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_B3;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_B4;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_B5;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_B6;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_BMUX;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_BO5;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_BO6;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_B_CY;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_B_XOR;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_C;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_C1;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_C2;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_C3;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_C4;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_C5;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_C6;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_CLK;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_CO5;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_CO6;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_CQ;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_C_CY;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_C_XOR;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_D;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_D1;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_D2;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_D3;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_D4;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_D5;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_D6;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_DO5;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_DO6;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_D_CY;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_D_XOR;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X118Y123_SR;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_A;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_A1;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_A2;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_A3;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_A4;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_A5;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_A6;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_AO5;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_AO6;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_AQ;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_A_CY;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_A_XOR;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_B;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_B1;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_B2;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_B3;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_B4;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_B5;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_B6;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_BMUX;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_BO5;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_BO6;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_B_CY;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_B_XOR;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_C;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_C1;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_C2;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_C3;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_C4;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_C5;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_C6;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_CLK;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_CO5;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_CO6;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_CQ;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_C_CY;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_C_XOR;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_D;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_D1;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_D2;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_D3;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_D4;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_D5;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_D6;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_DO5;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_DO6;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_D_CY;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_D_XOR;
  wire [0:0] CLBLL_R_X77Y123_SLICE_X119Y123_SR;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_A;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_A1;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_A2;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_A3;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_A4;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_A5;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_A6;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_AMUX;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_AO5;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_AO6;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_A_CY;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_A_XOR;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_B;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_B1;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_B2;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_B3;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_B4;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_B5;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_B6;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_BO5;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_BO6;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_BQ;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_B_CY;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_B_XOR;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_C;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_C1;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_C2;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_C3;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_C4;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_C5;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_C6;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_CLK;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_CO5;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_CO6;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_C_CY;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_C_XOR;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_D;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_D1;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_D2;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_D3;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_D4;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_D5;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_D6;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_DO5;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_DO6;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_D_CY;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_D_XOR;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X118Y124_SR;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_A;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_A1;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_A2;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_A3;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_A4;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_A5;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_A6;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_AO5;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_AO6;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_AQ;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_A_CY;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_A_XOR;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_B;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_B1;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_B2;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_B3;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_B4;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_B5;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_B6;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_BO5;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_BO6;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_BQ;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_B_CY;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_B_XOR;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_C;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_C1;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_C2;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_C3;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_C4;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_C5;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_C6;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_CLK;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_CO5;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_CO6;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_CQ;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_C_CY;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_C_XOR;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_D;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_D1;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_D2;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_D3;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_D4;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_D5;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_D6;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_DO5;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_DO6;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_D_CY;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_D_XOR;
  wire [0:0] CLBLL_R_X77Y124_SLICE_X119Y124_SR;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_A;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_A1;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_A2;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_A3;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_A4;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_A5;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_A5Q;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_A6;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_AMUX;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_AO5;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_AO6;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_AQ;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_A_CY;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_A_XOR;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_B;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_B1;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_B2;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_B3;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_B4;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_B5;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_B6;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_BMUX;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_BO5;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_BO6;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_BQ;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_B_CY;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_B_XOR;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_C;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_C1;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_C2;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_C3;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_C4;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_C5;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_C6;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_CLK;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_CO5;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_CO6;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_CQ;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_C_CY;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_C_XOR;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_D;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_D1;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_D2;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_D3;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_D4;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_D5;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_D6;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_DO5;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_DO6;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_D_CY;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_D_XOR;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_SR;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_A;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_A1;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_A2;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_A3;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_A4;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_A5;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_A6;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_AO5;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_AO6;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_A_CY;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_A_XOR;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_B;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_B1;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_B2;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_B3;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_B4;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_B5;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_B6;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_BO5;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_BO6;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_B_CY;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_B_XOR;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_C;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_C1;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_C2;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_C3;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_C4;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_C5;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_C6;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_CO5;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_CO6;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_C_CY;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_C_XOR;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_D;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_D1;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_D2;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_D3;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_D4;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_D5;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_D6;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_DO5;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_DO6;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_D_CY;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_D_XOR;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_A;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_A1;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_A2;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_A3;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_A4;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_A5;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_A6;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_AMUX;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_AO5;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_AO6;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_AQ;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_AX;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_A_CY;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_A_XOR;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_B;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_B1;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_B2;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_B3;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_B4;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_B5;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_B6;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_BO5;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_BO6;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_BQ;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_BX;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_B_CY;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_B_XOR;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_C;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_C1;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_C2;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_C3;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_C4;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_C5;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_C6;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_CLK;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_CO5;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_CO6;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_C_CY;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_C_XOR;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_D;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_D1;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_D2;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_D3;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_D4;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_D5;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_D6;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_DO5;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_DO6;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_D_CY;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_D_XOR;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X118Y126_SR;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_A;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_A1;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_A2;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_A3;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_A4;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_A5;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_A6;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_AO5;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_AO6;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_A_CY;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_A_XOR;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_B;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_B1;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_B2;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_B3;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_B4;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_B5;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_B6;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_BO5;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_BO6;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_B_CY;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_B_XOR;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_C;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_C1;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_C2;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_C3;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_C4;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_C5;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_C6;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_CO5;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_CO6;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_C_CY;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_C_XOR;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_D;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_D1;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_D2;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_D3;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_D4;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_D5;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_D6;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_DO5;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_DO6;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_D_CY;
  wire [0:0] CLBLL_R_X77Y126_SLICE_X119Y126_D_XOR;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_A;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_A1;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_A2;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_A3;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_A4;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_A5;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_A6;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_AO5;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_AO6;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_AQ;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_A_CY;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_A_XOR;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_B;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_B1;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_B2;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_B3;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_B4;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_B5;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_B6;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_BO5;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_BO6;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_B_CY;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_B_XOR;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_C;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_C1;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_C2;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_C3;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_C4;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_C5;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_C6;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_CLK;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_CO5;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_CO6;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_C_CY;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_C_XOR;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_D;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_D1;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_D2;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_D3;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_D4;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_D5;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_D6;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_DO5;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_DO6;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_D_CY;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_D_XOR;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X118Y127_SR;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_A;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_A1;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_A2;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_A3;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_A4;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_A5;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_A6;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_AMUX;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_AO5;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_AO6;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_AQ;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_A_CY;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_A_XOR;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_B;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_B1;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_B2;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_B3;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_B4;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_B5;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_B6;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_BO5;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_BO6;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_B_CY;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_B_XOR;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_C;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_C1;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_C2;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_C3;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_C4;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_C5;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_C6;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_CLK;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_CO5;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_CO6;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_C_CY;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_C_XOR;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_D;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_D1;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_D2;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_D3;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_D4;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_D5;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_D6;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_DO5;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_DO6;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_D_CY;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_D_XOR;
  wire [0:0] CLBLL_R_X77Y127_SLICE_X119Y127_SR;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_A;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_A1;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_A2;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_A3;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_A4;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_A5;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_A6;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_AMUX;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_AO5;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_AO6;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_AQ;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_AX;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_A_CY;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_A_XOR;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_B;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_B1;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_B2;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_B3;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_B4;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_B5;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_B5Q;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_B6;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_BMUX;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_BO5;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_BO6;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_BQ;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_B_CY;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_B_XOR;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_C;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_C1;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_C2;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_C3;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_C4;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_C5;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_C6;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_CLK;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_CMUX;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_CO5;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_CO6;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_CQ;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_CX;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_C_CY;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_C_XOR;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_D;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_D1;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_D2;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_D3;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_D4;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_D5;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_D6;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_DO5;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_DO6;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_D_CY;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_D_XOR;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X118Y128_SR;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_A;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_A1;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_A2;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_A3;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_A4;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_A5;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_A5Q;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_A6;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_AMUX;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_AO5;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_AO6;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_AQ;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_AX;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_A_CY;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_A_XOR;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_B;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_B1;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_B2;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_B3;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_B4;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_B5;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_B6;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_BO5;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_BO6;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_BQ;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_B_CY;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_B_XOR;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_C;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_C1;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_C2;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_C3;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_C4;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_C5;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_C6;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_CLK;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_CO5;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_CO6;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_CQ;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_C_CY;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_C_XOR;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_D;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_D1;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_D2;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_D3;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_D4;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_D5;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_D6;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_DO5;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_DO6;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_DQ;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_D_CY;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_D_XOR;
  wire [0:0] CLBLL_R_X77Y128_SLICE_X119Y128_SR;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_A;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_A1;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_A2;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_A3;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_A4;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_A5;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_A6;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_AO5;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_AO6;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_AQ;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_A_CY;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_A_XOR;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_B;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_B1;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_B2;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_B3;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_B4;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_B5;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_B6;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_BO5;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_BO6;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_BQ;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_B_CY;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_B_XOR;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_C;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_C1;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_C2;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_C3;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_C4;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_C5;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_C6;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_CLK;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_CO5;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_CO6;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_CQ;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_C_CY;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_C_XOR;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_D;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_D1;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_D2;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_D3;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_D4;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_D5;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_D6;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_DO5;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_DO6;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_DQ;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_D_CY;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_D_XOR;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_SR;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_A;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_A1;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_A2;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_A3;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_A4;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_A5;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_A6;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_AMUX;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_AO5;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_AO6;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_A_CY;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_A_XOR;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_B;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_B1;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_B2;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_B3;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_B4;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_B5;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_B6;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_BO5;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_BO6;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_BQ;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_B_CY;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_B_XOR;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_C;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_C1;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_C2;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_C3;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_C4;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_C5;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_C6;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_CLK;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_CMUX;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_CO5;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_CO6;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_C_CY;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_C_XOR;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_D;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_D1;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_D2;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_D3;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_D4;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_D5;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_D6;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_DO5;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_DO6;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_D_CY;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_D_XOR;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_SR;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_A;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_A1;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_A2;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_A3;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_A4;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_A5;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_A6;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_AMUX;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_AO5;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_AO6;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_AQ;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_A_CY;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_A_XOR;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_B;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_B1;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_B2;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_B3;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_B4;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_B5;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_B6;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_BO5;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_BO6;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_BQ;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_B_CY;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_B_XOR;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_C;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_C1;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_C2;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_C3;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_C4;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_C5;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_C6;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_CLK;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_CO5;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_CO6;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_CQ;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_C_CY;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_C_XOR;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_D;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_D1;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_D2;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_D3;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_D4;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_D5;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_D6;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_DMUX;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_DO5;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_DO6;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_D_CY;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_D_XOR;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_SR;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_A;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_A1;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_A2;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_A3;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_A4;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_A5;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_A6;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_AMUX;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_AO5;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_AO6;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_AQ;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_AX;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_A_CY;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_A_XOR;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_B;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_B1;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_B2;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_B3;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_B4;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_B5;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_B6;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_BO5;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_BO6;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_BQ;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_B_CY;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_B_XOR;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_C;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_C1;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_C2;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_C3;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_C4;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_C5;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_C6;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_CLK;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_CO5;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_CO6;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_C_CY;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_C_XOR;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_D;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_D1;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_D2;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_D3;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_D4;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_D5;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_D6;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_DO5;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_DO6;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_D_CY;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_D_XOR;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_SR;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_A;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_A1;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_A2;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_A3;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_A4;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_A5;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_A6;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_AO5;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_AO6;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_A_CY;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_A_XOR;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_B;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_B1;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_B2;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_B3;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_B4;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_B5;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_B6;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_BO5;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_BO6;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_B_CY;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_B_XOR;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_C;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_C1;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_C2;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_C3;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_C4;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_C5;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_C6;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_CO5;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_CO6;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_C_CY;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_C_XOR;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_D;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_D1;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_D2;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_D3;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_D4;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_D5;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_D6;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_DO5;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_DO6;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_D_CY;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_D_XOR;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_A;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_A1;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_A2;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_A3;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_A4;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_A5;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_A6;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_AO5;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_AO6;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_AQ;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_A_CY;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_A_XOR;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_B;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_B1;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_B2;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_B3;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_B4;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_B5;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_B6;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_BO5;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_BO6;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_BQ;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_B_CY;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_B_XOR;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_C;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_C1;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_C2;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_C3;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_C4;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_C5;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_C6;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_CLK;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_CO5;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_CO6;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_C_CY;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_C_XOR;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_D;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_D1;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_D2;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_D3;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_D4;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_D5;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_D6;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_DO5;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_DO6;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_D_CY;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_D_XOR;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_SR;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_A;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_A1;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_A2;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_A3;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_A4;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_A5;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_A5Q;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_A6;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_AMUX;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_AO5;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_AO6;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_AQ;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_AX;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_A_CY;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_A_XOR;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_B;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_B1;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_B2;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_B3;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_B4;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_B5;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_B6;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_BO5;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_BO6;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_BQ;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_B_CY;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_B_XOR;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_C;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_C1;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_C2;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_C3;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_C4;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_C5;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_C6;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_CLK;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_CO5;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_CO6;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_C_CY;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_C_XOR;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_D;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_D1;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_D2;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_D3;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_D4;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_D5;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_D6;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_DO5;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_DO6;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_D_CY;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_D_XOR;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X122Y104_SR;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_A;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_A1;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_A2;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_A3;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_A4;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_A5;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_A6;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_AO5;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_AO6;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_A_CY;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_A_XOR;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_B;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_B1;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_B2;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_B3;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_B4;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_B5;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_B6;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_BO5;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_BO6;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_B_CY;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_B_XOR;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_C;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_C1;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_C2;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_C3;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_C4;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_C5;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_C6;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_CO5;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_CO6;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_C_CY;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_C_XOR;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_D;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_D1;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_D2;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_D3;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_D4;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_D5;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_D6;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_DO5;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_DO6;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_D_CY;
  wire [0:0] CLBLL_R_X79Y104_SLICE_X123Y104_D_XOR;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_A;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_A1;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_A2;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_A3;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_A4;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_A5;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_A5Q;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_A6;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_AMUX;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_AO5;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_AO6;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_AQ;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_AX;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_A_CY;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_A_XOR;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_B;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_B1;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_B2;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_B3;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_B4;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_B5;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_B6;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_BO5;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_BO6;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_BQ;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_B_CY;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_B_XOR;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_C;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_C1;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_C2;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_C3;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_C4;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_C5;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_C6;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_CLK;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_CO5;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_CO6;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_CQ;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_C_CY;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_C_XOR;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_D;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_D1;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_D2;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_D3;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_D4;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_D5;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_D6;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_DO5;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_DO6;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_D_CY;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_D_XOR;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X122Y127_SR;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_A;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_A1;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_A2;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_A3;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_A4;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_A5;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_A6;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_AO5;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_AO6;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_A_CY;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_A_XOR;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_B;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_B1;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_B2;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_B3;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_B4;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_B5;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_B6;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_BO5;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_BO6;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_B_CY;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_B_XOR;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_C;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_C1;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_C2;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_C3;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_C4;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_C5;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_C6;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_CO5;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_CO6;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_C_CY;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_C_XOR;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_D;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_D1;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_D2;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_D3;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_D4;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_D5;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_D6;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_DO5;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_DO6;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_D_CY;
  wire [0:0] CLBLL_R_X79Y127_SLICE_X123Y127_D_XOR;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_A;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_A1;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_A2;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_A3;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_A4;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_A5;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_A6;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_AO5;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_AO6;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_AQ;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_A_CY;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_A_XOR;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_B;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_B1;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_B2;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_B3;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_B4;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_B5;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_B6;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_BO5;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_BO6;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_BQ;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_B_CY;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_B_XOR;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_C;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_C1;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_C2;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_C3;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_C4;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_C5;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_C6;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_CLK;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_CO5;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_CO6;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_CQ;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_C_CY;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_C_XOR;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_D;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_D1;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_D2;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_D3;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_D4;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_D5;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_D6;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_DO5;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_DO6;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_DQ;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_D_CY;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_D_XOR;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X122Y128_SR;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_A;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_A1;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_A2;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_A3;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_A4;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_A5;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_A6;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_AO5;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_AO6;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_A_CY;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_A_XOR;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_B;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_B1;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_B2;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_B3;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_B4;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_B5;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_B6;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_BO5;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_BO6;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_B_CY;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_B_XOR;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_C;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_C1;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_C2;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_C3;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_C4;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_C5;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_C6;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_CO5;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_CO6;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_C_CY;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_C_XOR;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_D;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_D1;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_D2;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_D3;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_D4;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_D5;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_D6;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_DO5;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_DO6;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_D_CY;
  wire [0:0] CLBLL_R_X79Y128_SLICE_X123Y128_D_XOR;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_A;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_A1;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_A2;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_A3;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_A4;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_A5;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_A6;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_AO5;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_AO6;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_AQ;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_AX;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_A_CY;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_A_XOR;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_B;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_B1;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_B2;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_B3;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_B4;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_B5;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_B6;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_BO5;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_BO6;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_B_CY;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_B_XOR;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_C;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_C1;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_C2;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_C3;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_C4;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_C5;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_C6;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_CLK;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_CO5;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_CO6;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_C_CY;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_C_XOR;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_D;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_D1;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_D2;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_D3;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_D4;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_D5;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_D6;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_DO5;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_DO6;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_D_CY;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_D_XOR;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X122Y135_SR;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_A;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_A1;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_A2;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_A3;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_A4;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_A5;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_A6;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_AO5;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_AO6;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_A_CY;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_A_XOR;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_B;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_B1;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_B2;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_B3;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_B4;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_B5;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_B6;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_BO5;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_BO6;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_B_CY;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_B_XOR;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_C;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_C1;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_C2;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_C3;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_C4;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_C5;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_C6;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_CO5;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_CO6;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_C_CY;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_C_XOR;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_D;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_D1;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_D2;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_D3;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_D4;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_D5;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_D6;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_DO5;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_DO6;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_D_CY;
  wire [0:0] CLBLL_R_X79Y135_SLICE_X123Y135_D_XOR;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_A;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_A1;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_A2;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_A3;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_A4;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_A5;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_A6;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_AO5;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_A_CY;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_A_XOR;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_B;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_B1;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_B2;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_B3;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_B4;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_B5;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_B6;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_BO5;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_BO6;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_B_CY;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_B_XOR;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_C;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_C1;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_C2;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_C3;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_C4;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_C5;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_C6;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_CO5;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_CO6;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_C_CY;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_C_XOR;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_D;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_D1;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_D2;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_D3;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_D4;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_D5;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_D6;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_DO5;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_DO6;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_D_CY;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X122Y96_D_XOR;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_A;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_A1;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_A2;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_A3;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_A4;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_A5;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_A6;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_AO5;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_AO6;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_A_CY;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_A_XOR;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_B;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_B1;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_B2;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_B3;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_B4;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_B5;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_B6;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_BO5;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_BO6;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_B_CY;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_B_XOR;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_C;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_C1;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_C2;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_C3;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_C4;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_C5;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_C6;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_CO5;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_CO6;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_C_CY;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_C_XOR;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_D;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_D1;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_D2;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_D3;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_D4;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_D5;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_D6;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_DO5;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_DO6;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_D_CY;
  wire [0:0] CLBLL_R_X79Y96_SLICE_X123Y96_D_XOR;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_A;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_A1;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_A2;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_A3;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_A4;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_A5;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_A6;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_AO5;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_AO6;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_A_CY;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_A_XOR;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_B;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_B1;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_B2;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_B3;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_B4;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_B5;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_B6;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_BO5;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_BO6;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_B_CY;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_B_XOR;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_C;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_C1;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_C2;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_C3;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_C4;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_C5;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_C6;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_CO5;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_CO6;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_C_CY;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_C_XOR;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_D;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_D1;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_D2;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_D3;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_D4;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_D5;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_D6;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_DO5;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_DO6;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_D_CY;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X122Y99_D_XOR;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_A;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_A1;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_A2;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_A3;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_A4;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_A5;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_A6;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_AO5;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_AO6;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_A_CY;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_A_XOR;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_B;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_B1;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_B2;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_B3;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_B4;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_B5;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_B6;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_BO5;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_BO6;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_B_CY;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_B_XOR;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_C;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_C1;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_C2;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_C3;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_C4;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_C5;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_C6;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_CO5;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_CO6;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_C_CY;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_C_XOR;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_D;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_D1;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_D2;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_D3;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_D4;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_D5;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_D6;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_DO5;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_DO6;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_D_CY;
  wire [0:0] CLBLL_R_X79Y99_SLICE_X123Y99_D_XOR;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_A;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_A1;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_A2;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_A3;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_A4;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_A5;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_A6;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_AO5;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_AO6;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_AQ;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_AX;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_A_CY;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_A_XOR;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_B;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_B1;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_B2;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_B3;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_B4;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_B5;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_B6;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_BO5;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_BO6;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_BQ;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_BX;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_B_CY;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_B_XOR;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_C;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_C1;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_C2;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_C3;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_C4;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_C5;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_C6;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_CLK;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_CO5;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_CO6;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_CQ;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_CX;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_C_CY;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_C_XOR;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_D;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_D1;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_D2;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_D3;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_D4;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_D5;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_D6;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_DO5;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_DO6;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_DQ;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_DX;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_D_CY;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_D_XOR;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X130Y130_SR;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_A;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_A1;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_A2;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_A3;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_A4;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_A5;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_A6;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_AO5;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_AO6;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_A_CY;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_A_XOR;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_B;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_B1;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_B2;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_B3;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_B4;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_B5;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_B6;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_BO5;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_BO6;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_B_CY;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_B_XOR;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_C;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_C1;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_C2;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_C3;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_C4;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_C5;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_C6;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_CO5;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_CO6;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_C_CY;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_C_XOR;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_D;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_D1;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_D2;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_D3;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_D4;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_D5;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_D6;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_DO5;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_DO6;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_D_CY;
  wire [0:0] CLBLL_R_X83Y130_SLICE_X131Y130_D_XOR;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_A;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_A1;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_A2;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_A3;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_A4;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_A5;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_A6;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_AO5;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_AO6;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_AQ;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_AX;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_A_CY;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_A_XOR;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_B;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_B1;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_B2;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_B3;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_B4;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_B5;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_B6;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_BO5;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_BO6;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_B_CY;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_B_XOR;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_C;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_C1;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_C2;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_C3;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_C4;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_C5;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_C6;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_CLK;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_CO5;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_CO6;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_C_CY;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_C_XOR;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_D;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_D1;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_D2;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_D3;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_D4;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_D5;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_D6;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_DO5;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_DO6;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_D_CY;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_D_XOR;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X130Y132_SR;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_A;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_A1;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_A2;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_A3;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_A4;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_A5;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_A6;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_AO5;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_AO6;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_A_CY;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_A_XOR;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_B;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_B1;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_B2;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_B3;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_B4;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_B5;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_B6;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_BO5;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_BO6;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_B_CY;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_B_XOR;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_C;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_C1;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_C2;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_C3;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_C4;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_C5;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_C6;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_CO5;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_CO6;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_C_CY;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_C_XOR;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_D;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_D1;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_D2;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_D3;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_D4;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_D5;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_D6;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_DO5;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_DO6;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_D_CY;
  wire [0:0] CLBLL_R_X83Y132_SLICE_X131Y132_D_XOR;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_A;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_A1;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_A2;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_A3;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_A4;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_A5;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_A5Q;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_A6;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_AMUX;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_AO5;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_AO6;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_AQ;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_A_CY;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_A_XOR;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_B;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_B1;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_B2;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_B3;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_B4;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_B5;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_B6;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_BO5;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_BO6;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_BQ;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_BX;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_B_CY;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_B_XOR;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_C;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_C1;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_C2;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_C3;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_C4;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_C5;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_C6;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_CLK;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_CO5;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_CO6;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_C_CY;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_C_XOR;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_D;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_D1;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_D2;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_D3;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_D4;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_D5;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_D6;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_DO5;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_DO6;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_D_CY;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_D_XOR;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X130Y94_SR;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_A;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_A1;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_A2;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_A3;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_A4;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_A5;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_A6;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_AO5;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_AO6;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_A_CY;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_A_XOR;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_B;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_B1;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_B2;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_B3;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_B4;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_B5;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_B6;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_BO5;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_BO6;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_B_CY;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_B_XOR;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_C;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_C1;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_C2;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_C3;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_C4;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_C5;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_C6;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_CO5;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_CO6;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_C_CY;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_C_XOR;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_D;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_D1;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_D2;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_D3;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_D4;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_D5;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_D6;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_DO5;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_DO6;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_D_CY;
  wire [0:0] CLBLL_R_X83Y94_SLICE_X131Y94_D_XOR;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_A;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_A1;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_A2;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_A3;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_A4;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_A5;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_A6;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_AO5;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_AO6;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_AQ;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_AX;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_A_CY;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_A_XOR;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_B;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_B1;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_B2;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_B3;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_B4;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_B5;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_B6;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_BO5;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_BO6;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_BQ;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_BX;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_B_CY;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_B_XOR;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_C;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_C1;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_C2;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_C3;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_C4;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_C5;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_C6;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_CLK;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_CO5;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_CO6;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_C_CY;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_C_XOR;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_D;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_D1;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_D2;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_D3;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_D4;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_D5;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_D6;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_DO5;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_DO6;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_D_CY;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_D_XOR;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_SR;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_A;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_A1;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_A2;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_A3;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_A4;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_A5;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_A6;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_AO5;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_AO6;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_A_CY;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_A_XOR;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_B;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_B1;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_B2;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_B3;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_B4;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_B5;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_B6;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_BO5;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_BO6;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_B_CY;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_B_XOR;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_C;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_C1;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_C2;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_C3;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_C4;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_C5;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_C6;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_CO5;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_CO6;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_C_CY;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_C_XOR;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_D;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_D1;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_D2;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_D3;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_D4;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_D5;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_D6;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_DO5;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_DO6;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_D_CY;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_D_XOR;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_A;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_A1;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_A2;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_A3;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_A4;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_A5;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_A6;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_AO5;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_AO6;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_AQ;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_AX;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_A_CY;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_A_XOR;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_B;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_B1;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_B2;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_B3;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_B4;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_B5;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_B6;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_BO5;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_BO6;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_B_CY;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_B_XOR;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_C;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_C1;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_C2;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_C3;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_C4;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_C5;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_C6;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_CLK;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_CO5;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_CO6;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_C_CY;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_C_XOR;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_D;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_D1;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_D2;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_D3;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_D4;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_D5;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_D6;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_DO5;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_DO6;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_D_CY;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_D_XOR;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_SR;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_A;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_A1;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_A2;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_A3;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_A4;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_A5;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_A6;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_AO5;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_AO6;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_A_CY;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_A_XOR;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_B;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_B1;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_B2;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_B3;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_B4;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_B5;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_B6;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_BO5;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_BO6;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_B_CY;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_B_XOR;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_C;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_C1;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_C2;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_C3;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_C4;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_C5;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_C6;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_CO5;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_CO6;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_C_CY;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_C_XOR;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_D;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_D1;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_D2;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_D3;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_D4;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_D5;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_D6;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_DO5;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_DO6;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_D_CY;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_D_XOR;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_A;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_A1;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_A2;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_A3;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_A4;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_A5;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_A6;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_AO5;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_AO6;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_AQ;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_AX;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_A_CY;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_A_XOR;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_B;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_B1;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_B2;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_B3;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_B4;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_B5;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_B6;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_BO5;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_BO6;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_BQ;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_BX;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_B_CY;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_B_XOR;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_C;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_C1;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_C2;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_C3;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_C4;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_C5;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_C6;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_CLK;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_CO5;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_CO6;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_C_CY;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_C_XOR;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_D;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_D1;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_D2;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_D3;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_D4;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_D5;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_D6;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_DO5;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_DO6;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_D_CY;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_D_XOR;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X90Y92_SR;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_A;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_A1;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_A2;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_A3;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_A4;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_A5;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_A6;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_AO5;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_AO6;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_A_CY;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_A_XOR;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_B;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_B1;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_B2;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_B3;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_B4;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_B5;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_B6;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_BO5;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_BO6;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_B_CY;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_B_XOR;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_C;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_C1;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_C2;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_C3;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_C4;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_C5;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_C6;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_CO5;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_CO6;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_C_CY;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_C_XOR;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_D;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_D1;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_D2;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_D3;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_D4;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_D5;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_D6;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_DO5;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_DO6;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_D_CY;
  wire [0:0] CLBLM_L_X60Y92_SLICE_X91Y92_D_XOR;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_A;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_A1;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_A2;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_A3;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_A4;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_A5;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_A6;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_AO5;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_AO6;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_AQ;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_AX;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_A_CY;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_A_XOR;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_B;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_B1;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_B2;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_B3;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_B4;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_B5;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_B6;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_BO5;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_BO6;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_BQ;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_BX;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_B_CY;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_B_XOR;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_C;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_C1;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_C2;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_C3;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_C4;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_C5;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_C6;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_CLK;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_CO5;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_CO6;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_CQ;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_CX;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_C_CY;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_C_XOR;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_D;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_D1;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_D2;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_D3;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_D4;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_D5;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_D6;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_DO5;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_DO6;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_D_CY;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_D_XOR;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X90Y94_SR;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_A;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_A1;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_A2;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_A3;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_A4;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_A5;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_A6;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_AO5;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_AO6;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_A_CY;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_A_XOR;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_B;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_B1;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_B2;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_B3;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_B4;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_B5;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_B6;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_BO5;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_BO6;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_B_CY;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_B_XOR;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_C;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_C1;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_C2;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_C3;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_C4;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_C5;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_C6;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_CO5;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_CO6;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_C_CY;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_C_XOR;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_D;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_D1;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_D2;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_D3;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_D4;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_D5;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_D6;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_DO5;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_DO6;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_D_CY;
  wire [0:0] CLBLM_L_X60Y94_SLICE_X91Y94_D_XOR;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_A;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_A1;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_A2;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_A3;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_A4;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_A5;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_A6;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_AO5;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_AO6;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_AX;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_A_CY;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_A_XOR;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_B;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_B1;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_B2;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_B3;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_B4;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_B5;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_B6;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_BO5;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_BO6;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_BQ;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_BX;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_B_CY;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_B_XOR;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_C;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_C1;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_C2;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_C3;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_C4;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_C5;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_C6;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_CLK;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_CO5;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_CO6;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_CX;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_C_CY;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_C_XOR;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_D;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_D1;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_D2;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_D3;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_D4;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_D5;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_D6;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_DO5;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_DO6;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_DQ;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_DX;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_D_CY;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_D_XOR;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_SR;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_A;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_A1;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_A2;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_A3;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_A4;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_A5;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_A6;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_AO5;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_AO6;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_AQ;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_AX;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_A_CY;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_A_XOR;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_B;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_B1;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_B2;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_B3;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_B4;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_B5;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_B6;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_BO5;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_BO6;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_B_CY;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_B_XOR;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_C;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_C1;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_C2;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_C3;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_C4;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_C5;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_C6;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_CLK;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_CO5;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_CO6;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_C_CY;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_C_XOR;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_D;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_D1;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_D2;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_D3;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_D4;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_D5;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_D6;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_DO5;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_DO6;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_D_CY;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_D_XOR;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_SR;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_A;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_A1;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_A2;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_A3;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_A4;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_A5;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_A6;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_AO5;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_AO6;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_AQ;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_AX;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_A_CY;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_A_XOR;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_B;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_B1;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_B2;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_B3;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_B4;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_B5;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_B6;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_BO5;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_BO6;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_BQ;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_BX;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_B_CY;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_B_XOR;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_C;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_C1;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_C2;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_C3;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_C4;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_C5;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_C6;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_CLK;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_CO5;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_CO6;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_CQ;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_CX;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_C_CY;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_C_XOR;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_D;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_D1;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_D2;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_D3;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_D4;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_D5;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_D6;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_DO5;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_DO6;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_DQ;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_DX;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_D_CY;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_D_XOR;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_SR;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_A;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_A1;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_A2;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_A3;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_A4;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_A5;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_A6;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_AO5;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_AO6;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_A_CY;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_A_XOR;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_B;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_B1;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_B2;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_B3;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_B4;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_B5;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_B6;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_BO5;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_BO6;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_B_CY;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_B_XOR;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_C;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_C1;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_C2;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_C3;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_C4;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_C5;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_C6;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_CO5;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_CO6;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_C_CY;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_C_XOR;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_D;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_D1;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_D2;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_D3;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_D4;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_D5;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_D6;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_DO5;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_DO6;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_D_CY;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_D_XOR;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_A;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_A1;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_A2;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_A3;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_A4;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_A5;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_A6;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_AO5;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_AO6;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_AQ;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_A_CY;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_A_XOR;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_B;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_B1;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_B2;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_B3;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_B4;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_B5;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_B6;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_BO5;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_BO6;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_B_CY;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_B_XOR;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_C;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_C1;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_C2;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_C3;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_C4;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_C5;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_C6;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_CLK;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_CO5;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_CO6;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_C_CY;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_C_XOR;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_D;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_D1;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_D2;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_D3;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_D4;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_D5;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_D6;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_DO5;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_DO6;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_D_CY;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_D_XOR;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_SR;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_A;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_A1;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_A2;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_A3;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_A4;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_A5;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_A6;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_AO5;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_AO6;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_A_CY;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_A_XOR;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_B;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_B1;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_B2;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_B3;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_B4;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_B5;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_B6;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_BO5;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_BO6;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_B_CY;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_B_XOR;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_C;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_C1;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_C2;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_C3;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_C4;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_C5;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_C6;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_CO5;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_CO6;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_C_CY;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_C_XOR;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_D;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_D1;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_D2;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_D3;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_D4;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_D5;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_D6;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_DO5;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_DO6;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_D_CY;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_D_XOR;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_A;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_A1;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_A2;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_A3;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_A4;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_A5;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_A6;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_AO5;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_AO6;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_AQ;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_AX;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_A_CY;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_A_XOR;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_B;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_B1;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_B2;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_B3;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_B4;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_B5;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_B6;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_BO5;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_BO6;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_B_CY;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_B_XOR;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_C;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_C1;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_C2;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_C3;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_C4;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_C5;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_C6;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_CLK;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_CO5;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_CO6;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_C_CY;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_C_XOR;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_D;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_D1;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_D2;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_D3;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_D4;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_D5;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_D6;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_DO5;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_DO6;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_D_CY;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_D_XOR;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_SR;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_A;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_A1;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_A2;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_A3;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_A4;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_A5;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_A6;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_AMUX;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_AO5;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_AO6;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_A_CY;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_A_XOR;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_B;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_B1;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_B2;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_B3;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_B4;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_B5;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_B6;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_BO5;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_BO6;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_B_CY;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_B_XOR;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_C;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_C1;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_C2;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_C3;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_C4;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_C5;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_C6;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_CO5;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_CO6;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_C_CY;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_C_XOR;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_D;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_D1;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_D2;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_D3;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_D4;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_D5;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_D6;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_DO5;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_DO6;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_D_CY;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_D_XOR;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_A;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_A1;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_A2;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_A3;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_A4;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_A5;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_A6;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_AO5;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_AO6;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_AQ;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_A_CY;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_A_XOR;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_B;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_B1;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_B2;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_B3;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_B4;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_B5;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_B6;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_BO5;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_BO6;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_BQ;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_B_CY;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_B_XOR;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_C;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_C1;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_C2;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_C3;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_C4;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_C5;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_C6;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_CLK;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_CO5;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_CO6;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_CQ;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_C_CY;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_C_XOR;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_D;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_D1;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_D2;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_D3;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_D4;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_D5;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_D6;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_DO5;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_DO6;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_D_CY;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_D_XOR;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_SR;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_A;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_A1;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_A2;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_A3;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_A4;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_A5;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_A6;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_AO5;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_AO6;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_AQ;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_A_CY;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_A_XOR;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_B;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_B1;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_B2;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_B3;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_B4;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_B5;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_B6;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_BO5;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_BO6;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_BQ;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_B_CY;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_B_XOR;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_C;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_C1;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_C2;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_C3;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_C4;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_C5;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_C6;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_CLK;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_CO5;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_CO6;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_CQ;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_C_CY;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_C_XOR;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_D;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_D1;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_D2;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_D3;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_D4;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_D5;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_D6;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_DO5;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_DO6;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_DQ;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_D_CY;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_D_XOR;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_SR;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_A;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_A1;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_A2;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_A3;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_A4;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_A5;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_A5Q;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_A6;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_AMUX;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_AO5;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_AO6;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_AQ;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_AX;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_A_CY;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_A_XOR;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_B;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_B1;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_B2;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_B3;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_B4;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_B5;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_B5Q;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_B6;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_BMUX;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_BO5;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_BO6;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_BQ;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_BX;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_B_CY;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_B_XOR;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_C;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_C1;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_C2;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_C3;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_C4;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_C5;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_C6;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_CLK;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_CO5;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_CO6;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_C_CY;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_C_XOR;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_D;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_D1;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_D2;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_D3;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_D4;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_D5;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_D6;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_DO5;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_DO6;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_D_CY;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_D_XOR;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_SR;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_A;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_A1;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_A2;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_A3;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_A4;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_A5;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_A6;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_AO5;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_AO6;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_AQ;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_A_CY;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_A_XOR;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_B;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_B1;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_B2;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_B3;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_B4;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_B5;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_B6;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_BO5;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_BO6;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_BQ;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_B_CY;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_B_XOR;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_C;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_C1;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_C2;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_C3;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_C4;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_C5;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_C6;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_CLK;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_CO5;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_CO6;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_CQ;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_C_CY;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_C_XOR;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_D;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_D1;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_D2;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_D3;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_D4;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_D5;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_D6;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_DO5;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_DO6;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_DQ;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_D_CY;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_D_XOR;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_SR;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_A;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_A1;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_A2;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_A3;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_A4;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_A5;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_A6;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_AO5;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_AO6;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_A_CY;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_A_XOR;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_B;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_B1;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_B2;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_B3;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_B4;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_B5;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_B6;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_BO5;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_BO6;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_B_CY;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_B_XOR;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_C;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_C1;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_C2;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_C3;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_C4;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_C5;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_C6;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_CO5;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_CO6;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_C_CY;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_C_XOR;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_D;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_D1;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_D2;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_D3;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_D4;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_D5;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_D6;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_DO5;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_DO6;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_D_CY;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_D_XOR;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_A;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_A1;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_A2;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_A3;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_A4;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_A5;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_A5Q;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_A6;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_AMUX;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_AO5;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_AO6;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_AQ;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_AX;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_A_CY;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_A_XOR;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_B;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_B1;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_B2;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_B3;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_B4;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_B5;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_B6;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_BO5;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_BO6;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_BQ;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_B_CY;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_B_XOR;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_C;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_C1;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_C2;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_C3;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_C4;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_C5;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_C6;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_CLK;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_CO5;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_CO6;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_CQ;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_C_CY;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_C_XOR;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_D;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_D1;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_D2;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_D3;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_D4;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_D5;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_D6;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_DO5;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_DO6;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_D_CY;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_D_XOR;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_SR;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_A;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_A1;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_A2;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_A3;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_A4;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_A5;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_A6;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_AO5;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_AO6;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_AQ;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_AX;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_A_CY;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_A_XOR;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_B;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_B1;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_B2;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_B3;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_B4;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_B5;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_B6;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_BO5;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_BO6;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_BQ;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_BX;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_B_CY;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_B_XOR;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_C;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_C1;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_C2;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_C3;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_C4;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_C5;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_C6;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_CLK;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_CO5;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_CO6;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_C_CY;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_C_XOR;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_D;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_D1;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_D2;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_D3;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_D4;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_D5;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_D6;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_DO5;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_DO6;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_D_CY;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_D_XOR;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_SR;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_A;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_A1;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_A2;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_A3;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_A4;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_A5;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_A6;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_AMUX;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_AO5;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_AO6;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_AQ;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_AX;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_A_CY;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_A_XOR;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_B;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_B1;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_B2;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_B3;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_B4;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_B5;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_B6;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_BO5;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_BO6;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_BQ;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_B_CY;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_B_XOR;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_C;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_C1;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_C2;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_C3;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_C4;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_C5;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_C6;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_CLK;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_CO5;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_CO6;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_CQ;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_C_CY;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_C_XOR;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_D;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_D1;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_D2;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_D3;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_D4;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_D5;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_D6;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_DO5;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_DO6;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_D_CY;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_D_XOR;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_SR;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_A;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_A1;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_A2;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_A3;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_A4;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_A5;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_A6;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_AMUX;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_AO5;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_AO6;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_A_CY;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_A_XOR;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_B;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_B1;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_B2;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_B3;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_B4;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_B5;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_B6;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_BO5;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_BO6;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_B_CY;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_B_XOR;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_C;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_C1;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_C2;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_C3;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_C4;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_C5;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_C6;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_CO5;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_CO6;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_C_CY;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_C_XOR;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_D;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_D1;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_D2;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_D3;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_D4;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_D5;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_D6;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_DO5;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_DO6;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_D_CY;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_D_XOR;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_A;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_A1;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_A2;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_A3;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_A4;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_A5;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_A5Q;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_A6;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_AMUX;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_AO5;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_AQ;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_AX;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_A_CY;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_A_XOR;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_B;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_B1;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_B2;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_B3;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_B4;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_B5;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_B6;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_BO5;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_BQ;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_B_CY;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_B_XOR;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_C;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_C1;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_C2;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_C3;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_C4;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_C5;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_C6;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_CLK;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_CMUX;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_CO5;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_CO6;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_C_CY;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_C_XOR;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_D;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_D1;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_D2;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_D3;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_D4;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_D5;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_D6;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_DO5;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_DO6;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_D_CY;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_D_XOR;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_SR;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_A;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_A1;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_A2;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_A3;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_A4;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_A5;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_A6;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_AO5;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_AO6;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_AQ;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_AX;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_A_CY;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_A_XOR;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_B;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_B1;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_B2;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_B3;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_B4;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_B5;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_B6;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_BO5;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_BO6;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_B_CY;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_B_XOR;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_C;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_C1;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_C2;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_C3;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_C4;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_C5;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_C6;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_CLK;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_CO5;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_CO6;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_C_CY;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_C_XOR;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_D;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_D1;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_D2;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_D3;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_D4;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_D5;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_D6;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_DO5;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_DO6;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_D_CY;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_D_XOR;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X92Y90_SR;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_A;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_A1;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_A2;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_A3;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_A4;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_A5;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_A6;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_AO5;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_AO6;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_A_CY;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_A_XOR;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_B;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_B1;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_B2;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_B3;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_B4;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_B5;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_B6;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_BO5;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_BO6;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_B_CY;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_B_XOR;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_C;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_C1;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_C2;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_C3;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_C4;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_C5;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_C6;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_CO5;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_CO6;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_C_CY;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_C_XOR;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_D;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_D1;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_D2;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_D3;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_D4;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_D5;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_D6;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_DO5;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_DO6;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_D_CY;
  wire [0:0] CLBLM_L_X62Y90_SLICE_X93Y90_D_XOR;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_A;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_A1;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_A2;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_A3;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_A4;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_A5;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_A6;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_AO5;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_AO6;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_AQ;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_AX;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_A_CY;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_A_XOR;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_B;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_B1;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_B2;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_B3;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_B4;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_B5;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_B6;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_BO5;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_BO6;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_BQ;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_BX;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_B_CY;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_B_XOR;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_C;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_C1;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_C2;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_C3;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_C4;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_C5;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_C6;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_CLK;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_CO5;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_CO6;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_C_CY;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_C_XOR;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_D;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_D1;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_D2;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_D3;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_D4;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_D5;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_D6;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_DO5;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_DO6;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_D_CY;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_D_XOR;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X92Y92_SR;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_A;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_A1;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_A2;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_A3;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_A4;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_A5;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_A6;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_AO5;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_AO6;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_A_CY;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_A_XOR;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_B;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_B1;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_B2;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_B3;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_B4;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_B5;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_B6;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_BO5;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_BO6;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_B_CY;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_B_XOR;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_C;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_C1;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_C2;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_C3;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_C4;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_C5;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_C6;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_CO5;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_CO6;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_C_CY;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_C_XOR;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_D;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_D1;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_D2;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_D3;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_D4;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_D5;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_D6;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_DO5;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_DO6;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_D_CY;
  wire [0:0] CLBLM_L_X62Y92_SLICE_X93Y92_D_XOR;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_A;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_A1;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_A2;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_A3;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_A4;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_A5;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_A6;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_AO5;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_AO6;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_AQ;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_AX;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_A_CY;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_A_XOR;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_B;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_B1;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_B2;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_B3;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_B4;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_B5;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_B6;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_BO5;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_BO6;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_BQ;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_BX;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_B_CY;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_B_XOR;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_C;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_C1;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_C2;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_C3;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_C4;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_C5;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_C6;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_CLK;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_CO5;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_CO6;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_CQ;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_CX;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_C_CY;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_C_XOR;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_D;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_D1;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_D2;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_D3;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_D4;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_D5;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_D6;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_DO5;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_DO6;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_D_CY;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_D_XOR;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_SR;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_A;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_A1;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_A2;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_A3;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_A4;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_A5;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_A6;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_AO5;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_AO6;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_A_CY;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_A_XOR;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_B;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_B1;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_B2;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_B3;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_B4;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_B5;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_B6;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_BO5;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_BO6;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_B_CY;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_B_XOR;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_C;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_C1;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_C2;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_C3;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_C4;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_C5;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_C6;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_CO5;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_CO6;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_C_CY;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_C_XOR;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_D;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_D1;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_D2;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_D3;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_D4;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_D5;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_D6;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_DO5;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_DO6;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_D_CY;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_D_XOR;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_A;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_A1;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_A2;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_A3;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_A4;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_A5;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_A6;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_AO5;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_AO6;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_A_CY;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_A_XOR;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_B;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_B1;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_B2;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_B3;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_B4;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_B5;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_B6;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_BO5;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_BO6;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_B_CY;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_B_XOR;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_C;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_C1;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_C2;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_C3;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_C4;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_C5;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_C6;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_CO5;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_CO6;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_C_CY;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_C_XOR;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_D;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_D1;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_D2;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_D3;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_D4;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_D5;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_D6;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_DO5;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_DO6;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_D_CY;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_D_XOR;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_A;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_A1;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_A2;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_A3;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_A4;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_A5;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_A6;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_AO5;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_AO6;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_AQ;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_A_CY;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_A_XOR;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_B;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_B1;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_B2;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_B3;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_B4;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_B5;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_B6;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_BO5;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_BO6;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_BQ;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_B_CY;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_B_XOR;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_C;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_C1;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_C2;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_C3;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_C4;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_C5;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_C6;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_CLK;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_CO5;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_CO6;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_C_CY;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_C_XOR;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_D;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_D1;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_D2;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_D3;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_D4;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_D5;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_D6;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_DO5;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_DO6;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_D_CY;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_D_XOR;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_SR;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_A;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_A1;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_A2;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_A3;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_A4;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_A5;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_A6;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_AO5;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_AO6;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_A_CY;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_A_XOR;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_B;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_B1;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_B2;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_B3;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_B4;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_B5;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_B6;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_BO5;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_BO6;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_B_CY;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_B_XOR;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_C;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_C1;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_C2;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_C3;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_C4;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_C5;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_C6;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_CO5;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_CO6;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_C_CY;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_C_XOR;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_D;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_D1;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_D2;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_D3;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_D4;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_D5;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_D6;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_DO5;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_DO6;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_D_CY;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_D_XOR;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_A;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_A1;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_A2;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_A3;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_A4;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_A5;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_A6;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_AO5;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_AO6;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_AQ;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_A_CY;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_A_XOR;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_B;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_B1;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_B2;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_B3;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_B4;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_B5;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_B6;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_BO5;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_BO6;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_BQ;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_B_CY;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_B_XOR;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_C;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_C1;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_C2;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_C3;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_C4;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_C5;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_C6;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_CLK;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_CO5;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_CO6;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_CQ;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_C_CY;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_C_XOR;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_D;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_D1;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_D2;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_D3;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_D4;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_D5;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_D6;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_DO5;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_DO6;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_D_CY;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_D_XOR;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_SR;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_A;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_A1;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_A2;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_A3;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_A4;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_A5;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_A6;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_AO5;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_AO6;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_A_CY;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_A_XOR;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_B;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_B1;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_B2;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_B3;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_B4;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_B5;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_B6;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_BO5;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_BO6;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_B_CY;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_B_XOR;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_C;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_C1;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_C2;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_C3;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_C4;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_C5;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_C6;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_CO5;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_CO6;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_C_CY;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_C_XOR;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_D;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_D1;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_D2;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_D3;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_D4;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_D5;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_D6;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_DO5;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_DO6;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_D_CY;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_D_XOR;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_A;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_A1;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_A2;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_A3;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_A4;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_A5;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_A6;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_AO5;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_AO6;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_AQ;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_A_CY;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_A_XOR;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_B;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_B1;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_B2;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_B3;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_B4;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_B5;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_B6;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_BO5;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_BO6;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_B_CY;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_B_XOR;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_C;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_C1;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_C2;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_C3;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_C4;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_C5;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_C6;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_CLK;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_CO5;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_CO6;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_C_CY;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_C_XOR;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_D;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_D1;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_D2;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_D3;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_D4;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_D5;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_D6;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_DO5;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_DO6;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_D_CY;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_D_XOR;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_SR;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_A;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_A1;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_A2;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_A3;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_A4;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_A5;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_A6;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_AO5;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_AO6;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_A_CY;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_A_XOR;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_B;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_B1;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_B2;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_B3;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_B4;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_B5;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_B6;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_BO5;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_BO6;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_B_CY;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_B_XOR;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_C;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_C1;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_C2;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_C3;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_C4;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_C5;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_C6;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_CO5;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_CO6;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_C_CY;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_C_XOR;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_D;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_D1;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_D2;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_D3;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_D4;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_D5;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_D6;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_DO5;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_DO6;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_D_CY;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_D_XOR;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_A;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_A1;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_A2;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_A3;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_A4;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_A5;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_A6;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_AO5;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_AO6;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_AQ;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_A_CY;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_A_XOR;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_B;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_B1;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_B2;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_B3;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_B4;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_B5;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_B6;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_BO5;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_BO6;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_B_CY;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_B_XOR;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_C;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_C1;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_C2;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_C3;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_C4;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_C5;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_C6;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_CLK;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_CO5;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_CO6;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_C_CY;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_C_XOR;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_D;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_D1;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_D2;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_D3;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_D4;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_D5;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_D6;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_DO5;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_DO6;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_D_CY;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_D_XOR;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_SR;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_A;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_A1;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_A2;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_A3;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_A4;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_A5;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_A5Q;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_A6;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_AMUX;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_AO5;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_AO6;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_AQ;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_A_CY;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_A_XOR;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_B;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_B1;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_B2;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_B3;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_B4;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_B5;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_B5Q;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_B6;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_BMUX;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_BO5;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_BO6;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_BQ;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_B_CY;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_B_XOR;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_C;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_C1;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_C2;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_C3;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_C4;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_C5;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_C5Q;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_C6;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_CLK;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_CMUX;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_CO5;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_CO6;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_CQ;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_C_CY;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_C_XOR;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_D;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_D1;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_D2;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_D3;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_D4;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_D5;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_D6;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_DO5;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_DO6;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_D_CY;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_D_XOR;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_SR;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_A;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_A1;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_A2;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_A3;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_A4;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_A5;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_A6;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_AO5;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_AO6;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_A_CY;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_A_XOR;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_B;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_B1;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_B2;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_B3;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_B4;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_B5;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_B6;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_BO5;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_BO6;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_B_CY;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_B_XOR;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_C;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_C1;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_C2;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_C3;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_C4;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_C5;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_C6;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_CO5;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_CO6;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_C_CY;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_C_XOR;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_D;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_D1;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_D2;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_D3;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_D4;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_D5;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_D6;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_DO5;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_DO6;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_D_CY;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_D_XOR;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_A;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_A1;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_A2;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_A3;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_A4;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_A5;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_A5Q;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_A6;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_AMUX;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_AO5;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_AO6;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_AQ;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_A_CY;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_A_XOR;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_B;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_B1;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_B2;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_B3;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_B4;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_B5;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_B6;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_BMUX;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_BO5;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_BO6;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_B_CY;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_B_XOR;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_C;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_C1;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_C2;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_C3;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_C4;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_C5;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_C6;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_CLK;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_CO5;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_CO6;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_CQ;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_C_CY;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_C_XOR;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_D;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_D1;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_D2;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_D3;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_D4;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_D5;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_D6;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_DO5;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_DO6;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_D_CY;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_D_XOR;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_SR;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_A;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_A1;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_A2;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_A3;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_A4;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_A5;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_A6;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_AO5;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_AO6;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_AQ;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_A_CY;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_A_XOR;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_B;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_B1;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_B2;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_B3;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_B4;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_B5;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_B6;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_BO5;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_BO6;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_BQ;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_B_CY;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_B_XOR;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_C;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_C1;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_C2;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_C3;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_C4;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_C5;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_C6;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_CLK;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_CO5;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_CO6;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_C_CY;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_C_XOR;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_D;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_D1;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_D2;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_D3;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_D4;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_D5;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_D6;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_DO5;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_DO6;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_D_CY;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_D_XOR;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_SR;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_A;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_A1;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_A2;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_A3;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_A4;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_A5;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_A6;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_AO5;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_AO6;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_AQ;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_A_CY;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_A_XOR;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_B;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_B1;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_B2;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_B3;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_B4;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_B5;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_B6;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_BO5;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_BO6;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_B_CY;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_B_XOR;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_C;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_C1;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_C2;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_C3;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_C4;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_C5;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_C6;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_CLK;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_CO5;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_CO6;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_C_CY;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_C_XOR;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_D;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_D1;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_D2;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_D3;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_D4;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_D5;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_D6;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_DO5;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_DO6;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_D_CY;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_D_XOR;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_SR;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_A;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_A1;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_A2;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_A3;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_A4;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_A5;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_A6;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_AO5;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_AO6;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_AQ;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_A_CY;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_A_XOR;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_B;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_B1;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_B2;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_B3;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_B4;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_B5;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_B6;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_BO5;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_BO6;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_BQ;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_B_CY;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_B_XOR;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_C;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_C1;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_C2;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_C3;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_C4;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_C5;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_C6;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_CLK;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_CO5;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_CO6;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_C_CY;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_C_XOR;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_D;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_D1;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_D2;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_D3;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_D4;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_D5;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_D6;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_DMUX;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_DO5;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_DO6;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_D_CY;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_D_XOR;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_SR;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_A;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_A1;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_A2;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_A3;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_A4;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_A5;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_A6;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_AO5;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_AO6;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_AQ;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_A_CY;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_A_XOR;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_B;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_B1;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_B2;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_B3;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_B4;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_B5;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_B6;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_BO5;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_BO6;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_BQ;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_B_CY;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_B_XOR;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_C;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_C1;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_C2;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_C3;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_C4;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_C5;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_C6;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_CLK;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_CO5;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_CO6;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_CQ;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_C_CY;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_C_XOR;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_D;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_D1;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_D2;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_D3;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_D4;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_D5;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_D6;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_DO5;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_DO6;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_DQ;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_D_CY;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_D_XOR;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_SR;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_A;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_A1;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_A2;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_A3;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_A4;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_A5;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_A6;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_AO5;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_AO6;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_AQ;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_A_CY;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_A_XOR;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_B;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_B1;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_B2;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_B3;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_B4;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_B5;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_B6;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_BO5;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_BO6;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_B_CY;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_B_XOR;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_C;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_C1;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_C2;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_C3;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_C4;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_C5;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_C6;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_CLK;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_CO5;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_CO6;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_C_CY;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_C_XOR;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_D;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_D1;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_D2;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_D3;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_D4;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_D5;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_D6;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_DO5;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_DO6;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_D_CY;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_D_XOR;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_SR;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_A;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_A1;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_A2;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_A3;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_A4;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_A5;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_A6;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_AMUX;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_AO5;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_AO6;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_A_CY;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_A_XOR;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_B;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_B1;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_B2;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_B3;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_B4;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_B5;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_B6;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_BMUX;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_BO5;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_BO6;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_B_CY;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_B_XOR;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_C;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_C1;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_C2;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_C3;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_C4;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_C5;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_C5Q;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_C6;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_CLK;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_CMUX;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_CO5;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_CO6;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_CQ;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_C_CY;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_C_XOR;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_D;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_D1;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_D2;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_D3;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_D4;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_D5;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_D6;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_DO5;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_DO6;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_D_CY;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_D_XOR;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_SR;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_A;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_A1;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_A2;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_A3;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_A4;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_A5;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_A6;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_AO5;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_AO6;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_AQ;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_A_CY;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_A_XOR;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_B;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_B1;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_B2;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_B3;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_B4;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_B5;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_B6;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_BO5;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_BO6;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_BQ;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_B_CY;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_B_XOR;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_C;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_C1;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_C2;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_C3;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_C4;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_C5;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_C6;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_CLK;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_CO5;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_CO6;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_CQ;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_C_CY;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_C_XOR;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_D;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_D1;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_D2;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_D3;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_D4;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_D5;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_D6;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_DO5;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_DO6;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_D_CY;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_D_XOR;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_SR;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_A;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_A1;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_A2;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_A3;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_A4;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_A5;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_A5Q;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_A6;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_AMUX;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_AO5;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_AO6;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_AQ;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_AX;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_A_CY;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_A_XOR;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_B;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_B1;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_B2;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_B3;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_B4;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_B5;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_B6;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_BMUX;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_BO5;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_BO6;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_BQ;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_BX;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_B_CY;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_B_XOR;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_C;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_C1;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_C2;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_C3;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_C4;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_C5;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_C6;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_CLK;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_CO5;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_CO6;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_CQ;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_C_CY;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_C_XOR;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_D;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_D1;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_D2;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_D3;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_D4;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_D5;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_D6;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_DMUX;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_DO5;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_DO6;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_D_CY;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_D_XOR;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_SR;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_A;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_A1;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_A2;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_A3;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_A4;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_A5;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_A6;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_AO5;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_AO6;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_AQ;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_A_CY;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_A_XOR;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_B;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_B1;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_B2;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_B3;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_B4;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_B5;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_B5Q;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_B6;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_BMUX;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_BO5;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_BO6;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_BQ;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_B_CY;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_B_XOR;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_C;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_C1;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_C2;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_C3;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_C4;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_C5;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_C5Q;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_C6;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_CLK;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_CMUX;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_CO5;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_CO6;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_CQ;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_C_CY;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_C_XOR;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_D;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_D1;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_D2;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_D3;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_D4;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_D5;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_D6;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_DO5;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_DO6;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_D_CY;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_D_XOR;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_SR;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_A;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_A1;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_A2;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_A3;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_A4;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_A5;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_A6;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_AO5;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_AO6;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_AQ;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_AX;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_A_CY;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_A_XOR;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_B;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_B1;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_B2;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_B3;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_B4;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_B5;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_B6;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_BO5;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_BO6;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_B_CY;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_B_XOR;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_C;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_C1;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_C2;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_C3;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_C4;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_C5;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_C6;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_CE;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_CLK;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_CO5;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_CO6;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_C_CY;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_C_XOR;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_D;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_D1;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_D2;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_D3;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_D4;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_D5;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_D6;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_DO5;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_DO6;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_D_CY;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_D_XOR;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X96Y122_SR;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_A;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_A1;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_A2;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_A3;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_A4;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_A5;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_A6;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_AO5;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_AO6;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_A_CY;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_A_XOR;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_B;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_B1;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_B2;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_B3;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_B4;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_B5;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_B6;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_BO5;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_BO6;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_B_CY;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_B_XOR;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_C;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_C1;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_C2;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_C3;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_C4;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_C5;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_C6;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_CO5;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_CO6;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_C_CY;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_C_XOR;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_D;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_D1;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_D2;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_D3;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_D4;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_D5;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_D6;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_DO5;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_DO6;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_D_CY;
  wire [0:0] CLBLM_L_X64Y122_SLICE_X97Y122_D_XOR;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_A;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_A1;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_A2;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_A3;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_A4;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_A5;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_A6;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_AO5;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_AO6;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_A_CY;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_A_XOR;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_B;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_B1;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_B2;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_B3;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_B4;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_B5;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_B6;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_BO5;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_BO6;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_B_CY;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_B_XOR;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_C;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_C1;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_C2;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_C3;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_C4;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_C5;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_C6;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_CO5;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_CO6;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_C_CY;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_C_XOR;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_D;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_D1;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_D2;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_D3;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_D4;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_D5;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_D6;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_DO5;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_DO6;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_D_CY;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_D_XOR;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_A;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_A1;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_A2;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_A3;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_A4;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_A5;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_A5Q;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_A6;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_AMUX;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_AO5;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_AO6;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_AQ;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_AX;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_A_CY;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_A_XOR;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_B;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_B1;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_B2;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_B3;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_B4;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_B5;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_B6;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_BO5;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_BO6;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_B_CY;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_B_XOR;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_C;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_C1;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_C2;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_C3;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_C4;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_C5;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_C6;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_CLK;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_CO5;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_CO6;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_C_CY;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_C_XOR;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_D;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_D1;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_D2;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_D3;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_D4;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_D5;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_D6;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_DO5;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_DO6;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_D_CY;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_D_XOR;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_SR;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_A;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_A1;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_A2;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_A3;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_A4;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_A5;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_A6;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_AO5;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_AO6;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_AQ;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_A_CY;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_A_XOR;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_B;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_B1;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_B2;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_B3;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_B4;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_B5;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_B6;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_BO5;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_BO6;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_BQ;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_B_CY;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_B_XOR;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_C;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_C1;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_C2;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_C3;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_C4;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_C5;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_C6;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_CLK;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_CO5;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_CO6;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_CQ;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_C_CY;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_C_XOR;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_D;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_D1;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_D2;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_D3;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_D4;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_D5;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_D6;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_DO5;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_DO6;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_DQ;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_D_CY;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_D_XOR;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_SR;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_A;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_A1;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_A2;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_A3;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_A4;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_A5;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_A5Q;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_A6;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_AMUX;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_AO5;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_AO6;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_AQ;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_A_CY;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_A_XOR;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_B;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_B1;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_B2;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_B3;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_B4;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_B5;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_B6;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_BMUX;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_BO5;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_BO6;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_B_CY;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_B_XOR;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_C;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_C1;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_C2;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_C3;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_C4;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_C5;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_C6;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_CLK;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_CO5;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_CO6;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_CQ;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_C_CY;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_C_XOR;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_D;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_D1;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_D2;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_D3;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_D4;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_D5;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_D6;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_DO5;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_DO6;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_DQ;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_D_CY;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_D_XOR;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_SR;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_A;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_A1;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_A2;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_A3;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_A4;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_A5;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_A6;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_AMUX;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_AO5;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_AO6;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_A_CY;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_A_XOR;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_B;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_B1;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_B2;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_B3;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_B4;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_B5;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_B6;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_BO5;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_BO6;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_BQ;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_B_CY;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_B_XOR;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_C;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_C1;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_C2;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_C3;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_C4;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_C5;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_C6;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_CLK;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_CO5;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_CO6;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_C_CY;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_C_XOR;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_D;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_D1;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_D2;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_D3;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_D4;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_D5;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_D6;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_DO5;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_DO6;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_D_CY;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_D_XOR;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_SR;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_A;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_A1;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_A2;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_A3;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_A4;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_A5;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_A6;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_AO5;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_AO6;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_A_CY;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_A_XOR;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_B;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_B1;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_B2;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_B3;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_B4;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_B5;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_B6;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_BO5;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_BO6;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_B_CY;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_B_XOR;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_C;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_C1;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_C2;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_C3;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_C4;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_C5;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_C6;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_CO5;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_CO6;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_C_CY;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_C_XOR;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_D;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_D1;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_D2;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_D3;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_D4;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_D5;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_D6;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_DO5;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_DO6;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_D_CY;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_D_XOR;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_A;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_A1;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_A2;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_A3;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_A4;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_A5;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_A5Q;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_A6;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_AMUX;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_AO5;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_AO6;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_AQ;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_A_CY;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_A_XOR;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_B;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_B1;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_B2;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_B3;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_B4;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_B5;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_B6;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_BMUX;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_BO5;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_BO6;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_BQ;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_B_CY;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_B_XOR;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_C;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_C1;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_C2;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_C3;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_C4;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_C5;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_C6;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_CLK;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_CO5;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_CO6;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_CQ;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_C_CY;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_C_XOR;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_D;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_D1;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_D2;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_D3;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_D4;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_D5;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_D6;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_DO5;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_DO6;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_D_CY;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_D_XOR;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_SR;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_A;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_A1;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_A2;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_A3;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_A4;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_A5;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_A5Q;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_A6;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_AMUX;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_AO5;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_AO6;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_AQ;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_A_CY;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_A_XOR;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_B;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_B1;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_B2;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_B3;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_B4;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_B5;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_B5Q;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_B6;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_BMUX;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_BO5;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_BO6;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_BQ;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_B_CY;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_B_XOR;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_C;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_C1;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_C2;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_C3;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_C4;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_C5;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_C6;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_CLK;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_CO5;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_CO6;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_C_CY;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_C_XOR;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_D;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_D1;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_D2;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_D3;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_D4;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_D5;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_D6;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_DO5;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_DO6;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_D_CY;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_D_XOR;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_SR;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_A;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_A1;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_A2;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_A3;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_A4;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_A5;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_A6;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_AO5;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_AO6;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_A_CY;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_A_XOR;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_B;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_B1;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_B2;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_B3;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_B4;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_B5;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_B6;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_BO5;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_BO6;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_B_CY;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_B_XOR;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_C;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_C1;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_C2;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_C3;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_C4;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_C5;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_C6;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_CO5;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_CO6;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_C_CY;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_C_XOR;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_D;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_D1;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_D2;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_D3;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_D4;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_D5;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_D6;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_DO5;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_DO6;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_D_CY;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X102Y100_D_XOR;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_A;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_A1;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_A2;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_A3;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_A4;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_A5;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_A6;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_AO5;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_AO6;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_A_CY;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_A_XOR;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_B;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_B1;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_B2;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_B3;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_B4;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_B5;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_B6;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_BO5;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_BO6;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_B_CY;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_B_XOR;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_C;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_C1;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_C2;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_C3;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_C4;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_C5;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_C6;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_CO5;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_CO6;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_C_CY;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_C_XOR;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_D;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_D1;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_D2;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_D3;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_D4;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_D5;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_D6;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_DO5;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_DO6;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_D_CY;
  wire [0:0] CLBLM_L_X68Y100_SLICE_X103Y100_D_XOR;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_A;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_A1;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_A2;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_A3;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_A4;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_A5;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_A5Q;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_A6;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_AMUX;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_AO5;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_AO6;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_AQ;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_AX;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_A_CY;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_A_XOR;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_B;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_B1;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_B2;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_B3;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_B4;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_B5;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_B6;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_BMUX;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_BO5;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_BO6;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_BQ;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_B_CY;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_B_XOR;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_C;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_C1;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_C2;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_C3;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_C4;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_C5;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_C6;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_CLK;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_CO5;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_CO6;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_CQ;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_C_CY;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_C_XOR;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_D;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_D1;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_D2;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_D3;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_D4;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_D5;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_D6;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_DO5;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_DO6;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_D_CY;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_D_XOR;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X102Y101_SR;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_A;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_A1;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_A2;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_A3;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_A4;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_A5;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_A6;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_AO5;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_AO6;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_A_CY;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_A_XOR;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_B;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_B1;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_B2;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_B3;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_B4;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_B5;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_B6;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_BO5;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_BO6;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_B_CY;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_B_XOR;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_C;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_C1;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_C2;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_C3;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_C4;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_C5;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_C6;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_CO5;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_CO6;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_C_CY;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_C_XOR;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_D;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_D1;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_D2;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_D3;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_D4;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_D5;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_D6;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_DO5;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_DO6;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_D_CY;
  wire [0:0] CLBLM_L_X68Y101_SLICE_X103Y101_D_XOR;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_A;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_A1;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_A2;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_A3;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_A4;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_A5;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_A6;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_AO5;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_AO6;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_AQ;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_A_CY;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_A_XOR;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_B;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_B1;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_B2;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_B3;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_B4;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_B5;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_B6;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_BO5;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_BO6;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_BQ;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_B_CY;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_B_XOR;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_C;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_C1;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_C2;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_C3;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_C4;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_C5;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_C6;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_CLK;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_CO5;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_CO6;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_CQ;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_C_CY;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_C_XOR;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_D;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_D1;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_D2;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_D3;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_D4;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_D5;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_D6;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_DO5;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_DO6;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_DQ;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_D_CY;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_D_XOR;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X102Y102_SR;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_A;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_A1;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_A2;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_A3;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_A4;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_A5;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_A6;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_AO5;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_AO6;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_A_CY;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_A_XOR;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_B;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_B1;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_B2;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_B3;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_B4;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_B5;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_B6;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_BO5;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_BO6;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_B_CY;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_B_XOR;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_C;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_C1;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_C2;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_C3;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_C4;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_C5;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_C6;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_CO5;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_CO6;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_C_CY;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_C_XOR;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_D;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_D1;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_D2;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_D3;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_D4;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_D5;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_D6;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_DO5;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_DO6;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_D_CY;
  wire [0:0] CLBLM_L_X68Y102_SLICE_X103Y102_D_XOR;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_A;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_A1;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_A2;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_A3;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_A4;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_A5;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_A6;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_AO5;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_AO6;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_AQ;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_A_CY;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_A_XOR;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_B;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_B1;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_B2;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_B3;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_B4;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_B5;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_B5Q;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_B6;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_BMUX;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_BO5;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_BO6;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_BQ;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_B_CY;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_B_XOR;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_C;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_C1;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_C2;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_C3;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_C4;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_C5;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_C6;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_CLK;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_CO5;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_CO6;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_CQ;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_C_CY;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_C_XOR;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_D;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_D1;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_D2;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_D3;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_D4;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_D5;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_D6;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_DO5;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_DO6;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_DQ;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_D_CY;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_D_XOR;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X102Y103_SR;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_A;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_A1;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_A2;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_A3;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_A4;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_A5;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_A6;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_AO5;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_AO6;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_A_CY;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_A_XOR;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_B;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_B1;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_B2;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_B3;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_B4;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_B5;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_B6;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_BO5;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_BO6;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_B_CY;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_B_XOR;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_C;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_C1;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_C2;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_C3;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_C4;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_C5;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_C6;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_CO5;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_CO6;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_C_CY;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_C_XOR;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_D;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_D1;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_D2;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_D3;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_D4;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_D5;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_D6;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_DO5;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_DO6;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_D_CY;
  wire [0:0] CLBLM_L_X68Y103_SLICE_X103Y103_D_XOR;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_A;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_A1;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_A2;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_A3;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_A4;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_A5;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_A6;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_AMUX;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_AO5;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_AO6;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_AQ;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_AX;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_A_CY;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_A_XOR;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_B;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_B1;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_B2;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_B3;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_B4;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_B5;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_B6;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_BO5;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_BO6;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_BQ;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_B_CY;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_B_XOR;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_C;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_C1;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_C2;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_C3;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_C4;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_C5;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_C6;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_CLK;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_CO5;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_CO6;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_CQ;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_C_CY;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_C_XOR;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_D;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_D1;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_D2;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_D3;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_D4;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_D5;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_D6;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_DO5;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_DO6;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_D_CY;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_D_XOR;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X102Y105_SR;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_A;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_A1;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_A2;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_A3;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_A4;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_A5;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_A6;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_AO5;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_AO6;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_AQ;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_A_CY;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_A_XOR;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_B;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_B1;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_B2;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_B3;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_B4;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_B5;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_B6;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_BO5;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_BO6;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_BQ;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_B_CY;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_B_XOR;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_C;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_C1;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_C2;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_C3;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_C4;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_C5;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_C6;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_CLK;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_CO5;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_CO6;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_C_CY;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_C_XOR;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_D;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_D1;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_D2;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_D3;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_D4;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_D5;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_D6;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_DO5;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_DO6;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_D_CY;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_D_XOR;
  wire [0:0] CLBLM_L_X68Y105_SLICE_X103Y105_SR;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_A;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_A1;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_A2;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_A3;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_A4;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_A5;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_A6;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_AMUX;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_AO5;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_AO6;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_A_CY;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_A_XOR;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_B;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_B1;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_B2;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_B3;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_B4;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_B5;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_B6;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_BO5;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_BO6;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_B_CY;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_B_XOR;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_C;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_C1;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_C2;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_C3;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_C4;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_C5;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_C6;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_CO5;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_CO6;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_C_CY;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_C_XOR;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_D;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_D1;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_D2;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_D3;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_D4;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_D5;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_D6;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_DO5;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_DO6;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_D_CY;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X102Y106_D_XOR;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_A;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_A1;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_A2;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_A3;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_A4;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_A5;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_A6;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_AMUX;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_AO5;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_AO6;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_A_CY;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_A_XOR;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_B;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_B1;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_B2;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_B3;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_B4;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_B5;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_B5Q;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_B6;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_BMUX;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_BO5;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_BO6;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_BQ;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_B_CY;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_B_XOR;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_C;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_C1;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_C2;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_C3;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_C4;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_C5;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_C6;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_CLK;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_CO5;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_CO6;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_CQ;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_C_CY;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_C_XOR;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_D;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_D1;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_D2;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_D3;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_D4;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_D5;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_D6;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_DO5;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_DO6;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_D_CY;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_D_XOR;
  wire [0:0] CLBLM_L_X68Y106_SLICE_X103Y106_SR;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_A;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_A1;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_A2;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_A3;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_A4;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_A5;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_A6;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_AMUX;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_AO5;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_AO6;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_A_CY;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_A_XOR;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_B;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_B1;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_B2;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_B3;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_B4;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_B5;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_B6;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_BO5;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_BO6;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_B_CY;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_B_XOR;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_C;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_C1;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_C2;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_C3;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_C4;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_C5;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_C6;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_CO5;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_CO6;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_C_CY;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_C_XOR;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_D;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_D1;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_D2;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_D3;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_D4;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_D5;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_D6;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_DO5;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_DO6;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_D_CY;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X102Y107_D_XOR;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_A;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_A1;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_A2;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_A3;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_A4;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_A5;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_A6;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_AO5;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_AO6;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_A_CY;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_A_XOR;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_B;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_B1;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_B2;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_B3;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_B4;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_B5;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_B6;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_BO5;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_BO6;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_B_CY;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_B_XOR;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_C;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_C1;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_C2;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_C3;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_C4;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_C5;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_C6;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_CMUX;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_CO5;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_CO6;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_C_CY;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_C_XOR;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_D;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_D1;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_D2;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_D3;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_D4;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_D5;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_D6;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_DO5;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_DO6;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_D_CY;
  wire [0:0] CLBLM_L_X68Y107_SLICE_X103Y107_D_XOR;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_A;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_A1;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_A2;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_A3;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_A4;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_A5;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_A5Q;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_A6;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_AMUX;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_AO5;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_AO6;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_AQ;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_A_CY;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_A_XOR;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_B;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_B1;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_B2;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_B3;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_B4;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_B5;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_B5Q;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_B6;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_BMUX;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_BO5;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_BO6;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_BQ;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_B_CY;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_B_XOR;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_C;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_C1;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_C2;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_C3;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_C4;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_C5;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_C6;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_CLK;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_CMUX;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_CO5;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_CO6;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_C_CY;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_C_XOR;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_D;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_D1;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_D2;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_D3;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_D4;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_D5;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_D6;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_DO5;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_DO6;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_D_CY;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_D_XOR;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X102Y108_SR;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_A;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_A1;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_A2;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_A3;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_A4;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_A5;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_A5Q;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_A6;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_AMUX;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_AO5;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_AO6;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_AQ;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_A_CY;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_A_XOR;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_B;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_B1;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_B2;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_B3;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_B4;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_B5;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_B6;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_BO5;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_BO6;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_BQ;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_B_CY;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_B_XOR;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_C;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_C1;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_C2;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_C3;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_C4;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_C5;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_C6;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_CLK;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_CO5;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_CO6;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_C_CY;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_C_XOR;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_D;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_D1;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_D2;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_D3;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_D4;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_D5;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_D6;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_DO5;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_DO6;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_D_CY;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_D_XOR;
  wire [0:0] CLBLM_L_X68Y108_SLICE_X103Y108_SR;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_A;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_A1;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_A2;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_A3;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_A4;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_A5;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_A5Q;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_A6;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_AMUX;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_AO5;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_AO6;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_AQ;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_A_CY;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_A_XOR;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_B;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_B1;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_B2;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_B3;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_B4;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_B5;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_B6;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_BMUX;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_BO5;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_BO6;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_B_CY;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_B_XOR;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_C;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_C1;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_C2;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_C3;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_C4;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_C5;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_C6;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_CLK;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_CMUX;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_CO5;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_CO6;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_C_CY;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_C_XOR;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_D;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_D1;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_D2;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_D3;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_D4;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_D5;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_D6;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_DO5;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_DO6;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_D_CY;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_D_XOR;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X102Y109_SR;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_A;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_A1;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_A2;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_A3;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_A4;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_A5;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_A6;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_AO5;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_AO6;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_AQ;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_A_CY;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_A_XOR;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_B;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_B1;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_B2;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_B3;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_B4;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_B5;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_B5Q;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_B6;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_BMUX;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_BO5;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_BO6;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_BQ;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_B_CY;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_B_XOR;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_C;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_C1;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_C2;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_C3;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_C4;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_C5;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_C6;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_CLK;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_CO5;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_CO6;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_C_CY;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_C_XOR;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_D;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_D1;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_D2;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_D3;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_D4;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_D5;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_D6;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_DO5;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_DO6;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_D_CY;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_D_XOR;
  wire [0:0] CLBLM_L_X68Y109_SLICE_X103Y109_SR;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_A;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_A1;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_A2;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_A3;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_A4;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_A5;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_A6;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_AO5;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_AO6;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_A_CY;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_A_XOR;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_B;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_B1;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_B2;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_B3;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_B4;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_B5;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_B6;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_BO5;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_BO6;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_B_CY;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_B_XOR;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_C;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_C1;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_C2;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_C3;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_C4;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_C5;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_C6;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_CO5;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_CO6;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_C_CY;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_C_XOR;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_D;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_D1;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_D2;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_D3;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_D4;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_D5;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_D6;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_DO5;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_DO6;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_D_CY;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X102Y112_D_XOR;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_A;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_A1;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_A2;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_A3;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_A4;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_A5;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_A6;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_AO5;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_AO6;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_AQ;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_AX;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_A_CY;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_A_XOR;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_B;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_B1;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_B2;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_B3;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_B4;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_B5;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_B6;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_BO5;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_BO6;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_BQ;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_BX;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_B_CY;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_B_XOR;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_C;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_C1;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_C2;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_C3;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_C4;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_C5;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_C6;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_CLK;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_CO5;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_CO6;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_C_CY;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_C_XOR;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_D;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_D1;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_D2;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_D3;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_D4;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_D5;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_D6;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_DO5;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_DO6;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_D_CY;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_D_XOR;
  wire [0:0] CLBLM_L_X68Y112_SLICE_X103Y112_SR;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_A;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_A1;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_A2;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_A3;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_A4;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_A5;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_A6;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_AO5;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_AO6;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_AQ;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_AX;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_A_CY;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_A_XOR;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_B;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_B1;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_B2;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_B3;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_B4;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_B5;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_B6;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_BO5;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_BO6;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_B_CY;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_B_XOR;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_C;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_C1;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_C2;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_C3;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_C4;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_C5;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_C6;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_CE;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_CLK;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_CO5;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_CO6;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_C_CY;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_C_XOR;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_D;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_D1;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_D2;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_D3;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_D4;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_D5;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_D6;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_DO5;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_DO6;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_D_CY;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_D_XOR;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X102Y121_SR;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_A;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_A1;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_A2;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_A3;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_A4;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_A5;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_A6;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_AO5;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_AO6;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_A_CY;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_A_XOR;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_B;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_B1;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_B2;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_B3;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_B4;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_B5;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_B6;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_BO5;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_BO6;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_B_CY;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_B_XOR;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_C;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_C1;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_C2;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_C3;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_C4;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_C5;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_C6;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_CO5;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_CO6;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_C_CY;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_C_XOR;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_D;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_D1;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_D2;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_D3;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_D4;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_D5;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_D6;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_DO5;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_DO6;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_D_CY;
  wire [0:0] CLBLM_L_X68Y121_SLICE_X103Y121_D_XOR;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_A;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_A1;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_A2;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_A3;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_A4;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_A5;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_A5Q;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_A6;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_AMUX;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_AO5;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_AO6;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_AQ;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_AX;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_A_CY;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_A_XOR;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_B;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_B1;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_B2;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_B3;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_B4;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_B5;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_B6;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_BO5;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_BO6;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_B_CY;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_B_XOR;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_C;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_C1;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_C2;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_C3;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_C4;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_C5;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_C6;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_CLK;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_CO5;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_CO6;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_C_CY;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_C_XOR;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_D;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_D1;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_D2;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_D3;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_D4;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_D5;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_D6;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_DO5;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_DO6;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_D_CY;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_D_XOR;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X102Y95_SR;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_A;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_A1;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_A2;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_A3;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_A4;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_A5;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_A6;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_AO5;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_AO6;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_A_CY;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_A_XOR;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_B;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_B1;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_B2;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_B3;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_B4;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_B5;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_B6;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_BO5;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_BO6;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_B_CY;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_B_XOR;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_C;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_C1;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_C2;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_C3;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_C4;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_C5;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_C6;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_CO5;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_CO6;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_C_CY;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_C_XOR;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_D;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_D1;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_D2;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_D3;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_D4;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_D5;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_D6;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_DO5;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_DO6;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_D_CY;
  wire [0:0] CLBLM_L_X68Y95_SLICE_X103Y95_D_XOR;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_A;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_A1;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_A2;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_A3;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_A4;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_A5;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_A6;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_AO5;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_AO6;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_AQ;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_A_CY;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_A_XOR;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_B;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_B1;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_B2;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_B3;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_B4;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_B5;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_B6;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_BO5;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_BO6;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_B_CY;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_B_XOR;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_C;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_C1;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_C2;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_C3;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_C4;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_C5;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_C6;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_CLK;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_CMUX;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_CO5;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_CO6;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_C_CY;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_C_XOR;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_D;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_D1;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_D2;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_D3;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_D4;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_D5;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_D6;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_DO5;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_DO6;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_D_CY;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_D_XOR;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X102Y96_SR;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_A;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_A1;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_A2;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_A3;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_A4;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_A5;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_A6;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_AMUX;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_AO5;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_AO6;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_A_CY;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_A_XOR;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_B;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_B1;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_B2;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_B3;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_B4;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_B5;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_B6;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_BO5;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_BO6;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_B_CY;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_B_XOR;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_C;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_C1;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_C2;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_C3;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_C4;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_C5;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_C6;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_CO5;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_CO6;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_C_CY;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_C_XOR;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_D;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_D1;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_D2;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_D3;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_D4;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_D5;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_D6;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_DO5;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_DO6;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_D_CY;
  wire [0:0] CLBLM_L_X68Y96_SLICE_X103Y96_D_XOR;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_A;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_A1;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_A2;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_A3;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_A4;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_A5;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_A6;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_AMUX;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_AO5;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_AO6;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_AQ;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_AX;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_A_CY;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_A_XOR;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_B;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_B1;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_B2;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_B3;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_B4;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_B5;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_B6;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_BO5;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_BO6;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_B_CY;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_B_XOR;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_C;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_C1;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_C2;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_C3;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_C4;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_C5;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_C6;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_CLK;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_CO5;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_CO6;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_C_CY;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_C_XOR;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_D;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_D1;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_D2;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_D3;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_D4;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_D5;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_D6;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_DO5;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_DO6;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_D_CY;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_D_XOR;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X102Y97_SR;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_A;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_A1;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_A2;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_A3;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_A4;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_A5;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_A6;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_AO5;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_AO6;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_AQ;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_AX;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_A_CY;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_A_XOR;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_B;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_B1;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_B2;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_B3;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_B4;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_B5;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_B6;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_BO5;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_BO6;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_B_CY;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_B_XOR;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_C;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_C1;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_C2;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_C3;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_C4;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_C5;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_C6;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_CLK;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_CO5;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_CO6;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_C_CY;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_C_XOR;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_D;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_D1;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_D2;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_D3;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_D4;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_D5;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_D6;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_DO5;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_DO6;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_D_CY;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_D_XOR;
  wire [0:0] CLBLM_L_X68Y97_SLICE_X103Y97_SR;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_A;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_A1;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_A2;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_A3;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_A4;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_A5;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_A6;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_AO5;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_AO6;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_AQ;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_A_CY;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_A_XOR;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_B;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_B1;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_B2;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_B3;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_B4;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_B5;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_B6;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_BO5;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_BO6;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_BQ;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_B_CY;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_B_XOR;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_C;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_C1;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_C2;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_C3;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_C4;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_C5;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_C6;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_CLK;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_CO5;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_CO6;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_CQ;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_C_CY;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_C_XOR;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_D;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_D1;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_D2;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_D3;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_D4;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_D5;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_D6;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_DO5;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_DO6;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_DQ;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_D_CY;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_D_XOR;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X102Y98_SR;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_A;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_A1;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_A2;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_A3;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_A4;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_A5;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_A5Q;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_A6;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_AMUX;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_AO5;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_AO6;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_AQ;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_A_CY;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_A_XOR;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_B;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_B1;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_B2;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_B3;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_B4;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_B5;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_B6;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_BO5;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_BO6;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_BQ;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_B_CY;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_B_XOR;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_C;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_C1;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_C2;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_C3;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_C4;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_C5;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_C6;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_CLK;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_CO5;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_CO6;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_CQ;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_C_CY;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_C_XOR;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_D;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_D1;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_D2;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_D3;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_D4;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_D5;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_D6;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_DO5;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_DO6;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_D_CY;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_D_XOR;
  wire [0:0] CLBLM_L_X68Y98_SLICE_X103Y98_SR;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_A;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_A1;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_A2;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_A3;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_A4;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_A5;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_A6;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_AMUX;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_AO5;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_AO6;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_AQ;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_AX;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_A_CY;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_A_XOR;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_B;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_B1;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_B2;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_B3;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_B4;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_B5;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_B6;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_BMUX;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_BO5;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_BO6;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_B_CY;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_B_XOR;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_C;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_C1;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_C2;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_C3;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_C4;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_C5;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_C6;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_CLK;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_CO5;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_CO6;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_C_CY;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_C_XOR;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_D;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_D1;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_D2;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_D3;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_D4;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_D5;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_D6;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_DMUX;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_DO5;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_DO6;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_D_CY;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_D_XOR;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X102Y99_SR;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_A;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_A1;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_A2;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_A3;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_A4;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_A5;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_A6;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_AO5;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_AO6;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_AQ;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_A_CY;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_A_XOR;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_B;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_B1;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_B2;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_B3;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_B4;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_B5;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_B6;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_BO5;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_BO6;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_BQ;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_B_CY;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_B_XOR;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_C;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_C1;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_C2;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_C3;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_C4;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_C5;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_C5Q;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_C6;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_CLK;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_CMUX;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_CO5;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_CO6;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_CQ;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_C_CY;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_C_XOR;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_D;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_D1;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_D2;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_D3;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_D4;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_D5;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_D5Q;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_D6;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_DMUX;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_DO5;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_DO6;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_DQ;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_D_CY;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_D_XOR;
  wire [0:0] CLBLM_L_X68Y99_SLICE_X103Y99_SR;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_A;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_A1;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_A2;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_A3;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_A4;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_A5;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_A5Q;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_A6;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_AMUX;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_AO5;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_AO6;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_AQ;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_AX;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_A_CY;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_A_XOR;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_B;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_B1;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_B2;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_B3;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_B4;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_B5;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_B6;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_BO5;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_BO6;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_BQ;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_B_CY;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_B_XOR;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_C;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_C1;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_C2;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_C3;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_C4;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_C5;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_C6;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_CLK;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_CO5;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_CO6;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_CQ;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_C_CY;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_C_XOR;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_D;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_D1;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_D2;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_D3;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_D4;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_D5;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_D6;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_DO5;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_DO6;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_D_CY;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_D_XOR;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X104Y100_SR;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_A;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_A1;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_A2;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_A3;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_A4;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_A5;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_A5Q;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_A6;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_AMUX;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_AO5;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_AO6;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_AQ;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_A_CY;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_A_XOR;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_B;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_B1;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_B2;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_B3;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_B4;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_B5;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_B5Q;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_B6;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_BMUX;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_BO5;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_BO6;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_BQ;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_B_CY;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_B_XOR;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_C;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_C1;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_C2;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_C3;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_C4;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_C5;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_C6;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_CLK;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_CO5;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_CO6;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_CQ;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_CX;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_C_CY;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_C_XOR;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_D;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_D1;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_D2;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_D3;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_D4;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_D5;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_D6;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_DO5;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_DO6;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_D_CY;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_D_XOR;
  wire [0:0] CLBLM_L_X70Y100_SLICE_X105Y100_SR;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_A;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_A1;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_A2;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_A3;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_A4;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_A5;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_A6;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_AMUX;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_AO5;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_AO6;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_AQ;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_AX;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_A_CY;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_A_XOR;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_B;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_B1;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_B2;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_B3;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_B4;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_B5;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_B6;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_BO5;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_BO6;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_BQ;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_B_CY;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_B_XOR;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_C;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_C1;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_C2;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_C3;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_C4;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_C5;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_C6;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_CLK;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_CO5;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_CO6;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_CQ;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_C_CY;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_C_XOR;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_D;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_D1;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_D2;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_D3;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_D4;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_D5;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_D6;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_DO5;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_DO6;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_D_CY;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_D_XOR;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X104Y101_SR;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_A;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_A1;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_A2;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_A3;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_A4;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_A5;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_A6;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_AMUX;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_AO5;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_AO6;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_AQ;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_AX;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_A_CY;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_A_XOR;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_B;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_B1;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_B2;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_B3;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_B4;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_B5;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_B6;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_BO5;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_BO6;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_BQ;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_B_CY;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_B_XOR;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_C;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_C1;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_C2;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_C3;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_C4;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_C5;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_C6;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_CLK;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_CO5;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_CO6;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_C_CY;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_C_XOR;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_D;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_D1;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_D2;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_D3;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_D4;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_D5;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_D6;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_DO5;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_DO6;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_D_CY;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_D_XOR;
  wire [0:0] CLBLM_L_X70Y101_SLICE_X105Y101_SR;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_A;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_A1;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_A2;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_A3;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_A4;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_A5;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_A6;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_AO5;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_AO6;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_AQ;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_A_CY;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_A_XOR;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_B;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_B1;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_B2;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_B3;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_B4;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_B5;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_B6;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_BO5;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_BO6;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_B_CY;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_B_XOR;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_C;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_C1;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_C2;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_C3;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_C4;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_C5;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_C6;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_CLK;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_CO5;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_CO6;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_C_CY;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_C_XOR;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_D;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_D1;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_D2;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_D3;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_D4;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_D5;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_D6;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_DO5;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_DO6;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_D_CY;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_D_XOR;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X104Y102_SR;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_A;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_A1;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_A2;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_A3;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_A4;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_A5;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_A6;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_AO5;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_AO6;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_AQ;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_A_CY;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_A_XOR;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_B;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_B1;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_B2;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_B3;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_B4;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_B5;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_B6;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_BO5;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_BO6;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_BQ;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_B_CY;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_B_XOR;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_C;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_C1;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_C2;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_C3;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_C4;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_C5;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_C6;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_CLK;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_CO5;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_CO6;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_CQ;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_C_CY;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_C_XOR;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_D;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_D1;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_D2;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_D3;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_D4;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_D5;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_D6;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_DO5;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_DO6;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_D_CY;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_D_XOR;
  wire [0:0] CLBLM_L_X70Y102_SLICE_X105Y102_SR;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_A;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_A1;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_A2;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_A3;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_A4;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_A5;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_A6;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_AO5;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_AO6;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_AQ;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_A_CY;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_A_XOR;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_B;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_B1;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_B2;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_B3;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_B4;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_B5;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_B5Q;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_B6;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_BMUX;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_BO5;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_BO6;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_BQ;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_B_CY;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_B_XOR;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_C;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_C1;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_C2;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_C3;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_C4;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_C5;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_C5Q;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_C6;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_CLK;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_CMUX;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_CO5;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_CO6;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_CQ;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_C_CY;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_C_XOR;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_D;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_D1;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_D2;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_D3;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_D4;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_D5;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_D6;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_DMUX;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_DO5;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_DO6;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_D_CY;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_D_XOR;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X104Y103_SR;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_A;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_A1;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_A2;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_A3;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_A4;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_A5;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_A6;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_AO5;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_AO6;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_AQ;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_A_CY;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_A_XOR;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_B;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_B1;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_B2;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_B3;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_B4;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_B5;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_B6;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_BO5;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_BO6;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_BQ;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_B_CY;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_B_XOR;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_C;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_C1;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_C2;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_C3;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_C4;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_C5;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_C6;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_CLK;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_CMUX;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_CO5;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_CO6;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_C_CY;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_C_XOR;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_D;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_D1;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_D2;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_D3;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_D4;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_D5;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_D6;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_DMUX;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_DO5;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_DO6;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_D_CY;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_D_XOR;
  wire [0:0] CLBLM_L_X70Y103_SLICE_X105Y103_SR;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_A;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_A1;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_A2;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_A3;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_A4;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_A5;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_A5Q;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_A6;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_AMUX;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_AO5;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_AO6;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_AQ;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_AX;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_A_CY;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_A_XOR;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_B;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_B1;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_B2;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_B3;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_B4;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_B5;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_B6;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_BO5;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_BO6;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_BQ;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_B_CY;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_B_XOR;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_C;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_C1;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_C2;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_C3;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_C4;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_C5;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_C6;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_CLK;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_CMUX;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_CO5;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_CO6;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_C_CY;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_C_XOR;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_D;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_D1;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_D2;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_D3;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_D4;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_D5;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_D6;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_DO5;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_DO6;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_D_CY;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_D_XOR;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X104Y104_SR;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_A;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_A1;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_A2;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_A3;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_A4;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_A5;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_A6;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_AO5;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_AO6;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_AQ;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_A_CY;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_A_XOR;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_B;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_B1;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_B2;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_B3;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_B4;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_B5;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_B6;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_BO5;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_BO6;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_BQ;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_B_CY;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_B_XOR;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_C;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_C1;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_C2;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_C3;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_C4;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_C5;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_C6;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_CLK;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_CO5;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_CO6;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_CQ;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_C_CY;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_C_XOR;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_D;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_D1;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_D2;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_D3;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_D4;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_D5;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_D5Q;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_D6;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_DMUX;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_DO5;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_DO6;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_DQ;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_D_CY;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_D_XOR;
  wire [0:0] CLBLM_L_X70Y104_SLICE_X105Y104_SR;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_A;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_A1;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_A2;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_A3;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_A4;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_A5;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_A6;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_AO5;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_AO6;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_AQ;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_A_CY;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_A_XOR;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_B;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_B1;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_B2;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_B3;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_B4;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_B5;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_B6;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_BO5;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_BO6;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_B_CY;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_B_XOR;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_C;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_C1;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_C2;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_C3;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_C4;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_C5;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_C6;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_CLK;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_CO5;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_CO6;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_C_CY;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_C_XOR;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_D;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_D1;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_D2;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_D3;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_D4;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_D5;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_D6;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_DO5;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_DO6;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_D_CY;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_D_XOR;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X104Y105_SR;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_A;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_A1;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_A2;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_A3;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_A4;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_A5;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_A5Q;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_A6;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_AMUX;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_AO5;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_AO6;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_AQ;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_A_CY;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_A_XOR;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_B;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_B1;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_B2;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_B3;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_B4;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_B5;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_B6;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_BO5;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_BO6;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_BQ;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_B_CY;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_B_XOR;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_C;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_C1;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_C2;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_C3;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_C4;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_C5;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_C6;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_CLK;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_CO5;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_CO6;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_C_CY;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_C_XOR;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_D;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_D1;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_D2;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_D3;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_D4;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_D5;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_D6;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_DO5;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_DO6;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_D_CY;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_D_XOR;
  wire [0:0] CLBLM_L_X70Y105_SLICE_X105Y105_SR;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_A;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_A1;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_A2;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_A3;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_A4;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_A5;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_A5Q;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_A6;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_AMUX;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_AO5;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_AO6;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_AQ;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_AX;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_A_CY;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_A_XOR;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_B;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_B1;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_B2;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_B3;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_B4;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_B5;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_B6;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_BO5;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_BO6;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_BQ;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_BX;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_B_CY;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_B_XOR;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_C;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_C1;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_C2;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_C3;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_C4;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_C5;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_C6;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_CLK;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_CO5;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_CO6;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_C_CY;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_C_XOR;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_D;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_D1;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_D2;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_D3;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_D4;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_D5;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_D6;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_DO5;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_DO6;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_D_CY;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_D_XOR;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X104Y106_SR;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_A;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_A1;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_A2;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_A3;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_A4;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_A5;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_A5Q;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_A6;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_AMUX;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_AO5;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_AO6;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_AQ;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_AX;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_A_CY;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_A_XOR;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_B;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_B1;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_B2;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_B3;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_B4;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_B5;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_B6;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_BO5;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_BO6;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_BQ;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_B_CY;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_B_XOR;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_C;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_C1;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_C2;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_C3;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_C4;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_C5;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_C6;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_CLK;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_CO5;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_CO6;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_C_CY;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_C_XOR;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_D;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_D1;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_D2;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_D3;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_D4;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_D5;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_D6;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_DO5;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_DO6;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_D_CY;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_D_XOR;
  wire [0:0] CLBLM_L_X70Y106_SLICE_X105Y106_SR;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_A;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_A1;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_A2;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_A3;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_A4;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_A5;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_A6;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_AO5;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_AO6;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_AQ;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_A_CY;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_A_XOR;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_B;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_B1;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_B2;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_B3;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_B4;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_B5;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_B6;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_BO5;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_BO6;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_BQ;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_B_CY;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_B_XOR;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_C;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_C1;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_C2;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_C3;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_C4;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_C5;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_C6;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_CLK;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_CO5;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_CO6;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_C_CY;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_C_XOR;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_D;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_D1;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_D2;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_D3;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_D4;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_D5;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_D6;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_DO5;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_DO6;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_D_CY;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_D_XOR;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X104Y107_SR;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_A;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_A1;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_A2;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_A3;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_A4;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_A5;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_A6;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_AO5;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_AO6;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_AQ;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_A_CY;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_A_XOR;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_B;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_B1;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_B2;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_B3;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_B4;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_B5;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_B6;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_BO5;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_BO6;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_BQ;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_B_CY;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_B_XOR;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_C;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_C1;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_C2;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_C3;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_C4;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_C5;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_C6;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_CLK;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_CO5;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_CO6;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_C_CY;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_C_XOR;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_D;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_D1;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_D2;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_D3;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_D4;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_D5;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_D6;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_DO5;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_DO6;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_D_CY;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_D_XOR;
  wire [0:0] CLBLM_L_X70Y107_SLICE_X105Y107_SR;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_A;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_A1;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_A2;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_A3;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_A4;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_A5;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_A6;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_AO5;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_AO6;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_A_CY;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_A_XOR;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_B;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_B1;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_B2;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_B3;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_B4;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_B5;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_B6;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_BO5;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_BO6;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_B_CY;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_B_XOR;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_C;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_C1;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_C2;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_C3;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_C4;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_C5;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_C6;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_CO5;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_CO6;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_C_CY;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_C_XOR;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_D;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_D1;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_D2;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_D3;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_D4;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_D5;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_D6;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_DO5;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_DO6;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_D_CY;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X104Y108_D_XOR;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_A;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_A1;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_A2;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_A3;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_A4;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_A5;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_A6;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_AMUX;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_AO5;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_AO6;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_A_CY;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_A_XOR;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_B;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_B1;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_B2;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_B3;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_B4;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_B5;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_B6;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_BO5;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_BO6;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_B_CY;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_B_XOR;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_C;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_C1;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_C2;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_C3;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_C4;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_C5;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_C6;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_CO5;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_CO6;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_C_CY;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_C_XOR;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_D;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_D1;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_D2;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_D3;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_D4;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_D5;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_D6;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_DO5;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_DO6;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_D_CY;
  wire [0:0] CLBLM_L_X70Y108_SLICE_X105Y108_D_XOR;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_A;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_A1;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_A2;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_A3;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_A4;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_A5;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_A5Q;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_A6;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_AMUX;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_AO5;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_AO6;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_AQ;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_A_CY;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_A_XOR;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_B;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_B1;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_B2;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_B3;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_B4;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_B5;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_B5Q;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_B6;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_BMUX;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_BO5;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_BO6;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_BQ;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_B_CY;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_B_XOR;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_C;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_C1;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_C2;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_C3;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_C4;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_C5;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_C6;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_CLK;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_CO5;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_CO6;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_C_CY;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_C_XOR;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_D;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_D1;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_D2;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_D3;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_D4;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_D5;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_D6;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_DO5;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_DO6;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_D_CY;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_D_XOR;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X104Y109_SR;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_A;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_A1;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_A2;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_A3;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_A4;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_A5;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_A6;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_AO5;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_AO6;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_AQ;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_AX;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_A_CY;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_A_XOR;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_B;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_B1;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_B2;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_B3;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_B4;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_B5;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_B6;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_BO5;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_BO6;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_B_CY;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_B_XOR;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_C;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_C1;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_C2;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_C3;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_C4;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_C5;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_C6;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_CLK;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_CO5;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_CO6;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_C_CY;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_C_XOR;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_D;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_D1;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_D2;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_D3;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_D4;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_D5;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_D6;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_DO5;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_DO6;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_D_CY;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_D_XOR;
  wire [0:0] CLBLM_L_X70Y109_SLICE_X105Y109_SR;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_A;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_A1;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_A2;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_A3;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_A4;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_A5;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_A6;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_AMUX;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_AO5;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_AO6;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_AQ;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_A_CY;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_A_XOR;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_B;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_B1;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_B2;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_B3;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_B4;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_B5;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_B5Q;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_B6;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_BMUX;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_BO5;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_BO6;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_BQ;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_B_CY;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_B_XOR;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_C;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_C1;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_C2;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_C3;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_C4;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_C5;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_C6;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_CLK;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_CO5;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_CO6;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_CQ;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_C_CY;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_C_XOR;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_D;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_D1;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_D2;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_D3;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_D4;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_D5;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_D6;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_DO5;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_DO6;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_D_CY;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_D_XOR;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X104Y110_SR;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_A;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_A1;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_A2;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_A3;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_A4;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_A5;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_A6;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_AO5;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_AO6;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_A_CY;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_A_XOR;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_B;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_B1;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_B2;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_B3;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_B4;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_B5;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_B6;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_BO5;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_BO6;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_B_CY;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_B_XOR;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_C;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_C1;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_C2;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_C3;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_C4;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_C5;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_C6;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_CO5;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_CO6;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_C_CY;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_C_XOR;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_D;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_D1;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_D2;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_D3;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_D4;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_D5;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_D6;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_DO5;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_DO6;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_D_CY;
  wire [0:0] CLBLM_L_X70Y110_SLICE_X105Y110_D_XOR;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_A;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_A1;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_A2;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_A3;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_A4;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_A5;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_A6;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_AMUX;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_AO5;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_AO6;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_AQ;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_AX;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_A_CY;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_A_XOR;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_B;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_B1;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_B2;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_B3;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_B4;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_B5;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_B6;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_BMUX;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_BO5;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_BO6;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_BQ;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_BX;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_B_CY;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_B_XOR;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_C;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_C1;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_C2;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_C3;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_C4;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_C5;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_C6;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_CLK;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_CMUX;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_CO5;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_CO6;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_C_CY;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_C_XOR;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_D;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_D1;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_D2;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_D3;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_D4;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_D5;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_D6;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_DO5;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_DO6;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_D_CY;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_D_XOR;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X104Y111_SR;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_A;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_A1;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_A2;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_A3;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_A4;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_A5;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_A6;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_AO5;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_AO6;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_AQ;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_A_CY;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_A_XOR;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_B;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_B1;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_B2;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_B3;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_B4;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_B5;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_B6;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_BO5;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_BO6;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_BQ;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_B_CY;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_B_XOR;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_C;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_C1;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_C2;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_C3;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_C4;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_C5;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_C6;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_CLK;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_CO5;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_CO6;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_C_CY;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_C_XOR;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_D;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_D1;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_D2;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_D3;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_D4;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_D5;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_D6;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_DO5;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_DO6;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_D_CY;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_D_XOR;
  wire [0:0] CLBLM_L_X70Y111_SLICE_X105Y111_SR;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_A;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_A1;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_A2;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_A3;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_A4;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_A5;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_A5Q;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_A6;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_AMUX;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_AO5;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_AO6;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_AQ;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_AX;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_A_CY;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_A_XOR;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_B;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_B1;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_B2;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_B3;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_B4;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_B5;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_B6;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_BMUX;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_BO5;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_BO6;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_B_CY;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_B_XOR;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_C;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_C1;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_C2;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_C3;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_C4;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_C5;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_C5Q;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_C6;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_CLK;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_CMUX;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_CO5;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_CO6;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_CQ;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_C_CY;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_C_XOR;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_D;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_D1;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_D2;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_D3;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_D4;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_D5;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_D6;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_DO5;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_DO6;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_DQ;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_D_CY;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_D_XOR;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X104Y112_SR;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_A;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_A1;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_A2;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_A3;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_A4;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_A5;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_A5Q;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_A6;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_AMUX;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_AO5;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_AO6;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_AQ;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_A_CY;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_A_XOR;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_B;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_B1;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_B2;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_B3;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_B4;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_B5;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_B5Q;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_B6;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_BMUX;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_BO5;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_BO6;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_BQ;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_B_CY;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_B_XOR;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_C;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_C1;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_C2;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_C3;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_C4;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_C5;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_C5Q;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_C6;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_CLK;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_CMUX;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_CO5;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_CO6;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_CQ;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_C_CY;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_C_XOR;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_D;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_D1;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_D2;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_D3;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_D4;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_D5;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_D5Q;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_D6;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_DMUX;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_DO5;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_DO6;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_DQ;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_D_CY;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_D_XOR;
  wire [0:0] CLBLM_L_X70Y112_SLICE_X105Y112_SR;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_A;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_A1;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_A2;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_A3;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_A4;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_A5;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_A5Q;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_A6;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_AMUX;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_AO5;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_AO6;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_AQ;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_A_CY;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_A_XOR;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_B;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_B1;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_B2;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_B3;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_B4;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_B5;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_B5Q;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_B6;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_BMUX;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_BO5;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_BO6;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_BQ;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_B_CY;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_B_XOR;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_C;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_C1;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_C2;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_C3;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_C4;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_C5;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_C6;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_CLK;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_CO5;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_CO6;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_CQ;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_C_CY;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_C_XOR;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_D;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_D1;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_D2;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_D3;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_D4;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_D5;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_D6;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_DO5;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_DO6;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_D_CY;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_D_XOR;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X104Y113_SR;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_A;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_A1;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_A2;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_A3;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_A4;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_A5;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_A6;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_AO5;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_AO6;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_A_CY;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_A_XOR;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_B;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_B1;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_B2;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_B3;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_B4;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_B5;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_B6;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_BO5;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_BO6;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_B_CY;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_B_XOR;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_C;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_C1;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_C2;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_C3;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_C4;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_C5;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_C6;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_CO5;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_CO6;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_C_CY;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_C_XOR;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_D;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_D1;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_D2;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_D3;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_D4;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_D5;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_D6;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_DO5;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_DO6;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_D_CY;
  wire [0:0] CLBLM_L_X70Y113_SLICE_X105Y113_D_XOR;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_A;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_A1;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_A2;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_A3;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_A4;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_A5;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_A5Q;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_A6;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_AMUX;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_AO5;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_AO6;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_AQ;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_AX;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_A_CY;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_A_XOR;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_B;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_B1;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_B2;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_B3;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_B4;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_B5;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_B6;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_BO5;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_BO6;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_B_CY;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_B_XOR;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_C;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_C1;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_C2;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_C3;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_C4;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_C5;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_C6;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_CLK;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_CO5;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_CO6;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_C_CY;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_C_XOR;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_D;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_D1;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_D2;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_D3;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_D4;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_D5;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_D6;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_DO5;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_DO6;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_D_CY;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_D_XOR;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X104Y114_SR;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_A;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_A1;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_A2;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_A3;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_A4;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_A5;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_A6;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_AO5;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_AO6;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_A_CY;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_A_XOR;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_B;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_B1;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_B2;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_B3;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_B4;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_B5;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_B6;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_BO5;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_BO6;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_B_CY;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_B_XOR;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_C;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_C1;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_C2;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_C3;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_C4;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_C5;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_C6;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_CO5;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_CO6;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_C_CY;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_C_XOR;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_D;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_D1;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_D2;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_D3;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_D4;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_D5;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_D6;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_DO5;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_DO6;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_D_CY;
  wire [0:0] CLBLM_L_X70Y114_SLICE_X105Y114_D_XOR;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_A;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_A1;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_A2;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_A3;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_A4;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_A5;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_A6;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_AO5;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_AO6;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_A_CY;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_A_XOR;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_B;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_B1;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_B2;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_B3;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_B4;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_B5;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_B6;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_BO5;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_BO6;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_B_CY;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_B_XOR;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_C;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_C1;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_C2;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_C3;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_C4;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_C5;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_C6;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_CO5;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_CO6;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_C_CY;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_C_XOR;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_D;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_D1;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_D2;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_D3;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_D4;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_D5;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_D6;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_DO5;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_DO6;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_D_CY;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_D_XOR;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_A;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_A1;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_A2;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_A3;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_A4;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_A5;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_A5Q;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_A6;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_AMUX;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_AO5;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_AO6;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_AQ;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_A_CY;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_A_XOR;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_B;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_B1;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_B2;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_B3;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_B4;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_B5;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_B6;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_BO5;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_BO6;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_B_CY;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_B_XOR;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_C;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_C1;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_C2;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_C3;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_C4;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_C5;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_C6;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_CLK;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_CO5;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_CO6;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_C_CY;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_C_XOR;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_D;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_D1;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_D2;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_D3;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_D4;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_D5;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_D6;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_DO5;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_DO6;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_D_CY;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_D_XOR;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_SR;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_A;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_A1;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_A2;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_A3;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_A4;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_A5;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_A5Q;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_A6;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_AMUX;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_AO5;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_AO6;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_AQ;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_A_CY;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_A_XOR;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_B;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_B1;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_B2;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_B3;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_B4;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_B5;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_B6;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_BO5;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_BO6;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_BQ;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_B_CY;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_B_XOR;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_C;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_C1;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_C2;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_C3;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_C4;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_C5;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_C6;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_CLK;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_CO5;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_CO6;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_C_CY;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_C_XOR;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_D;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_D1;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_D2;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_D3;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_D4;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_D5;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_D6;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_DO5;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_DO6;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_D_CY;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_D_XOR;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_SR;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_A;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_A1;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_A2;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_A3;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_A4;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_A5;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_A6;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_AO5;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_AO6;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_A_CY;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_A_XOR;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_B;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_B1;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_B2;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_B3;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_B4;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_B5;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_B6;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_BO5;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_BO6;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_B_CY;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_B_XOR;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_C;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_C1;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_C2;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_C3;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_C4;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_C5;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_C6;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_CO5;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_CO6;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_C_CY;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_C_XOR;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_D;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_D1;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_D2;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_D3;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_D4;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_D5;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_D6;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_DO5;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_DO6;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_D_CY;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_D_XOR;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_A;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_A1;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_A2;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_A3;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_A4;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_A5;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_A6;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_AO5;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_AO6;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_AQ;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_A_CY;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_A_XOR;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_B;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_B1;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_B2;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_B3;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_B4;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_B5;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_B6;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_BO5;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_BO6;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_BQ;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_B_CY;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_B_XOR;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_C;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_C1;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_C2;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_C3;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_C4;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_C5;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_C6;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_CLK;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_CO5;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_CO6;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_CQ;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_C_CY;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_C_XOR;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_D;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_D1;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_D2;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_D3;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_D4;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_D5;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_D6;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_DO5;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_DO6;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_D_CY;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_D_XOR;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_SR;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_A;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_A1;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_A2;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_A3;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_A4;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_A5;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_A6;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_AO5;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_AO6;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_A_CY;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_A_XOR;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_B;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_B1;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_B2;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_B3;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_B4;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_B5;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_B6;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_BO5;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_BO6;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_B_CY;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_B_XOR;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_C;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_C1;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_C2;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_C3;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_C4;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_C5;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_C6;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_CO5;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_CO6;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_C_CY;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_C_XOR;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_D;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_D1;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_D2;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_D3;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_D4;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_D5;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_D6;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_DO5;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_DO6;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_D_CY;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_D_XOR;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_A;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_A1;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_A2;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_A3;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_A4;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_A5;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_A5Q;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_A6;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_AMUX;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_AO5;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_AO6;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_AQ;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_A_CY;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_A_XOR;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_B;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_B1;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_B2;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_B3;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_B4;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_B5;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_B6;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_BO5;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_BO6;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_BQ;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_B_CY;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_B_XOR;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_C;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_C1;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_C2;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_C3;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_C4;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_C5;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_C6;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_CLK;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_CO5;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_CO6;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_CQ;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_C_CY;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_C_XOR;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_D;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_D1;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_D2;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_D3;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_D4;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_D5;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_D6;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_DO5;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_DO6;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_D_CY;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_D_XOR;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X104Y125_SR;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_A;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_A1;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_A2;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_A3;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_A4;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_A5;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_A6;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_AMUX;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_AO5;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_AO6;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_AQ;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_AX;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_A_CY;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_A_XOR;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_B;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_B1;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_B2;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_B3;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_B4;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_B5;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_B6;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_BMUX;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_BO5;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_BO6;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_BQ;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_BX;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_B_CY;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_B_XOR;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_C;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_C1;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_C2;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_C3;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_C4;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_C5;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_C6;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_CLK;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_CMUX;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_CO5;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_CO6;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_C_CY;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_C_XOR;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_D;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_D1;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_D2;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_D3;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_D4;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_D5;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_D6;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_DO5;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_DO6;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_D_CY;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_D_XOR;
  wire [0:0] CLBLM_L_X70Y125_SLICE_X105Y125_SR;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_A;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_A1;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_A2;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_A3;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_A4;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_A5;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_A6;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_AO5;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_AO6;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_AQ;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_A_CY;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_A_XOR;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_B;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_B1;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_B2;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_B3;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_B4;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_B5;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_B6;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_BO5;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_BO6;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_BQ;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_B_CY;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_B_XOR;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_C;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_C1;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_C2;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_C3;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_C4;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_C5;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_C6;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_CLK;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_CO5;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_CO6;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_CQ;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_C_CY;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_C_XOR;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_D;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_D1;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_D2;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_D3;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_D4;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_D5;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_D6;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_DO5;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_DO6;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_D_CY;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_D_XOR;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X104Y126_SR;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_A;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_A1;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_A2;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_A3;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_A4;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_A5;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_A6;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_AO5;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_AO6;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_AQ;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_A_CY;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_A_XOR;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_B;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_B1;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_B2;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_B3;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_B4;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_B5;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_B6;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_BO5;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_BO6;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_BQ;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_B_CY;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_B_XOR;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_C;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_C1;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_C2;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_C3;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_C4;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_C5;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_C6;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_CLK;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_CO5;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_CO6;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_C_CY;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_C_XOR;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_D;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_D1;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_D2;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_D3;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_D4;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_D5;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_D6;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_DO5;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_DO6;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_D_CY;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_D_XOR;
  wire [0:0] CLBLM_L_X70Y126_SLICE_X105Y126_SR;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_A;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_A1;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_A2;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_A3;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_A4;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_A5;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_A6;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_AMUX;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_AO5;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_AO6;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_AQ;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_AX;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_A_CY;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_A_XOR;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_B;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_B1;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_B2;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_B3;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_B4;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_B5;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_B6;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_BMUX;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_BO5;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_BO6;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_BQ;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_BX;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_B_CY;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_B_XOR;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_C;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_C1;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_C2;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_C3;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_C4;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_C5;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_C6;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_CLK;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_CO5;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_CO6;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_CQ;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_C_CY;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_C_XOR;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_D;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_D1;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_D2;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_D3;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_D4;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_D5;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_D6;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_DO5;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_DO6;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_DQ;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_D_CY;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_D_XOR;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_SR;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_A;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_A1;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_A2;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_A3;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_A4;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_A5;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_A6;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_AO5;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_AO6;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_AQ;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_AX;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_A_CY;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_A_XOR;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_B;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_B1;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_B2;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_B3;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_B4;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_B5;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_B6;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_BMUX;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_BO5;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_BO6;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_B_CY;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_B_XOR;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_C;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_C1;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_C2;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_C3;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_C4;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_C5;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_C6;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_CE;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_CLK;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_CO5;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_CO6;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_C_CY;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_C_XOR;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_D;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_D1;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_D2;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_D3;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_D4;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_D5;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_D6;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_DO5;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_DO6;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_D_CY;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_D_XOR;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_SR;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_A;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_A1;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_A2;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_A3;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_A4;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_A5;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_A6;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_AO5;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_AO6;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_AQ;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_A_CY;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_A_XOR;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_B;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_B1;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_B2;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_B3;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_B4;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_B5;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_B6;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_BO5;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_BO6;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_BQ;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_B_CY;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_B_XOR;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_C;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_C1;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_C2;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_C3;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_C4;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_C5;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_C6;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_CLK;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_CO5;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_CO6;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_CQ;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_C_CY;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_C_XOR;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_D;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_D1;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_D2;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_D3;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_D4;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_D5;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_D6;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_DO5;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_DO6;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_DQ;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_D_CY;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_D_XOR;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_SR;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_A;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_A1;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_A2;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_A3;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_A4;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_A5;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_A6;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_AO5;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_AO6;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_AQ;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_A_CY;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_A_XOR;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_B;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_B1;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_B2;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_B3;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_B4;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_B5;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_B6;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_BO5;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_BO6;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_BQ;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_B_CY;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_B_XOR;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_C;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_C1;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_C2;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_C3;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_C4;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_C5;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_C6;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_CLK;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_CO5;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_CO6;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_CQ;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_C_CY;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_C_XOR;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_D;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_D1;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_D2;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_D3;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_D4;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_D5;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_D6;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_DO5;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_DO6;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_DQ;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_D_CY;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_D_XOR;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_SR;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_A;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_A1;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_A2;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_A3;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_A4;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_A5;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_A6;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_AMUX;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_AO5;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_AO6;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_A_CY;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_A_XOR;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_B;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_B1;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_B2;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_B3;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_B4;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_B5;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_B6;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_BO5;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_BO6;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_BQ;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_B_CY;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_B_XOR;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_C;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_C1;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_C2;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_C3;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_C4;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_C5;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_C6;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_CLK;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_CO5;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_CO6;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_CQ;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_C_CY;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_C_XOR;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_D;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_D1;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_D2;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_D3;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_D4;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_D5;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_D6;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_DO5;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_DO6;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_DQ;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_D_CY;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_D_XOR;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X104Y130_SR;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_A;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_A1;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_A2;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_A3;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_A4;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_A5;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_A5Q;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_A6;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_AMUX;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_AO5;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_AO6;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_AQ;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_A_CY;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_A_XOR;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_B;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_B1;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_B2;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_B3;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_B4;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_B5;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_B6;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_BO5;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_BO6;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_BQ;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_B_CY;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_B_XOR;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_C;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_C1;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_C2;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_C3;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_C4;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_C5;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_C6;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_CLK;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_CO5;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_CO6;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_CQ;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_C_CY;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_C_XOR;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_D;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_D1;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_D2;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_D3;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_D4;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_D5;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_D6;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_DMUX;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_DO5;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_DO6;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_D_CY;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_D_XOR;
  wire [0:0] CLBLM_L_X70Y130_SLICE_X105Y130_SR;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_A;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_A1;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_A2;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_A3;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_A4;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_A5;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_A6;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_AO5;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_AO6;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_AQ;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_A_CY;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_A_XOR;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_B;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_B1;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_B2;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_B3;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_B4;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_B5;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_B6;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_BO5;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_BO6;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_BQ;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_B_CY;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_B_XOR;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_C;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_C1;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_C2;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_C3;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_C4;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_C5;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_C6;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_CLK;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_CO5;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_CO6;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_C_CY;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_C_XOR;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_D;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_D1;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_D2;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_D3;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_D4;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_D5;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_D6;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_DO5;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_DO6;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_D_CY;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_D_XOR;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X104Y131_SR;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_A;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_A1;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_A2;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_A3;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_A4;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_A5;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_A6;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_AO5;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_AO6;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_A_CY;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_A_XOR;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_B;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_B1;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_B2;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_B3;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_B4;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_B5;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_B6;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_BO5;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_BO6;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_B_CY;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_B_XOR;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_C;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_C1;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_C2;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_C3;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_C4;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_C5;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_C6;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_CO5;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_CO6;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_C_CY;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_C_XOR;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_D;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_D1;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_D2;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_D3;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_D4;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_D5;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_D6;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_DO5;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_DO6;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_D_CY;
  wire [0:0] CLBLM_L_X70Y131_SLICE_X105Y131_D_XOR;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_A;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_A1;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_A2;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_A3;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_A4;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_A5;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_A6;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_AO5;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_AO6;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_A_CY;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_A_XOR;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_B;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_B1;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_B2;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_B3;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_B4;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_B5;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_B6;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_BO5;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_BO6;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_B_CY;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_B_XOR;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_C;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_C1;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_C2;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_C3;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_C4;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_C5;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_C6;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_CO5;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_CO6;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_C_CY;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_C_XOR;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_D;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_D1;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_D2;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_D3;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_D4;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_D5;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_D6;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_DO5;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_DO6;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_D_CY;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X104Y132_D_XOR;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_A;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_A1;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_A2;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_A3;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_A4;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_A5;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_A6;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_AO5;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_AO6;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_AQ;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_AX;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_A_CY;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_A_XOR;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_B;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_B1;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_B2;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_B3;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_B4;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_B5;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_B6;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_BO5;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_BO6;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_BQ;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_BX;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_B_CY;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_B_XOR;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_C;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_C1;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_C2;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_C3;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_C4;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_C5;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_C6;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_CE;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_CLK;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_CO5;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_CO6;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_C_CY;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_C_XOR;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_D;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_D1;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_D2;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_D3;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_D4;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_D5;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_D6;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_DO5;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_DO6;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_D_CY;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_D_XOR;
  wire [0:0] CLBLM_L_X70Y132_SLICE_X105Y132_SR;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_A;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_A1;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_A2;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_A3;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_A4;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_A5;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_A5Q;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_A6;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_AMUX;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_AO5;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_AO6;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_AQ;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_AX;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_A_CY;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_A_XOR;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_B;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_B1;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_B2;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_B3;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_B4;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_B5;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_B6;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_BO5;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_BO6;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_BQ;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_B_CY;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_B_XOR;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_C;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_C1;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_C2;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_C3;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_C4;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_C5;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_C6;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_CLK;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_CMUX;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_CO5;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_CO6;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_C_CY;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_C_XOR;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_D;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_D1;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_D2;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_D3;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_D4;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_D5;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_D6;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_DO5;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_DO6;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_D_CY;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_D_XOR;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X104Y133_SR;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_A;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_A1;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_A2;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_A3;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_A4;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_A5;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_A6;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_AO5;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_AO6;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_AQ;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_A_CY;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_A_XOR;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_B;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_B1;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_B2;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_B3;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_B4;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_B5;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_B6;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_BO5;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_BO6;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_BQ;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_B_CY;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_B_XOR;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_C;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_C1;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_C2;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_C3;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_C4;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_C5;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_C6;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_CLK;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_CO5;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_CO6;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_CQ;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_C_CY;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_C_XOR;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_D;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_D1;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_D2;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_D3;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_D4;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_D5;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_D6;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_DO5;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_DO6;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_DQ;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_D_CY;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_D_XOR;
  wire [0:0] CLBLM_L_X70Y133_SLICE_X105Y133_SR;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_A;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_A1;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_A2;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_A3;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_A4;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_A5;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_A6;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_AO5;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_AO6;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_AQ;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_A_CY;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_A_XOR;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_B;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_B1;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_B2;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_B3;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_B4;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_B5;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_B6;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_BO5;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_BO6;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_BQ;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_B_CY;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_B_XOR;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_C;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_C1;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_C2;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_C3;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_C4;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_C5;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_C6;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_CLK;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_CMUX;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_CO5;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_CO6;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_C_CY;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_C_XOR;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_D;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_D1;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_D2;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_D3;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_D4;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_D5;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_D6;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_DO5;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_DO6;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_D_CY;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_D_XOR;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X104Y134_SR;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_A;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_A1;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_A2;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_A3;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_A4;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_A5;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_A6;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_AO5;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_AO6;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_AQ;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_A_CY;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_A_XOR;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_B;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_B1;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_B2;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_B3;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_B4;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_B5;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_B6;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_BO5;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_BO6;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_BQ;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_B_CY;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_B_XOR;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_C;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_C1;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_C2;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_C3;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_C4;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_C5;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_C6;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_CLK;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_CO5;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_CO6;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_CQ;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_C_CY;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_C_XOR;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_D;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_D1;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_D2;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_D3;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_D4;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_D5;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_D6;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_DMUX;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_DO5;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_DO6;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_D_CY;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_D_XOR;
  wire [0:0] CLBLM_L_X70Y134_SLICE_X105Y134_SR;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_A;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_A1;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_A2;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_A3;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_A4;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_A5;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_A6;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_AO5;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_AO6;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_AQ;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_A_CY;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_A_XOR;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_B;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_B1;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_B2;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_B3;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_B4;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_B5;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_B6;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_BO5;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_BO6;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_BQ;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_B_CY;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_B_XOR;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_C;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_C1;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_C2;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_C3;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_C4;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_C5;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_C6;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_CLK;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_CMUX;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_CO5;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_CO6;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_C_CY;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_C_XOR;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_D;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_D1;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_D2;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_D3;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_D4;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_D5;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_D6;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_DO5;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_DO6;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_D_CY;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_D_XOR;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X104Y135_SR;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_A;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_A1;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_A2;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_A3;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_A4;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_A5;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_A5Q;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_A6;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_AMUX;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_AO5;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_AO6;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_AQ;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_A_CY;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_A_XOR;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_B;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_B1;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_B2;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_B3;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_B4;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_B5;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_B6;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_BO5;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_BO6;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_B_CY;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_B_XOR;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_C;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_C1;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_C2;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_C3;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_C4;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_C5;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_C6;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_CLK;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_CO5;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_CO6;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_C_CY;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_C_XOR;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_D;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_D1;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_D2;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_D3;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_D4;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_D5;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_D6;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_DO5;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_DO6;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_D_CY;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_D_XOR;
  wire [0:0] CLBLM_L_X70Y135_SLICE_X105Y135_SR;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_A;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_A1;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_A2;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_A3;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_A4;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_A5;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_A6;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_AO5;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_AO6;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_AQ;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_A_CY;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_A_XOR;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_B;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_B1;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_B2;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_B3;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_B4;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_B5;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_B6;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_BO5;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_BO6;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_BQ;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_B_CY;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_B_XOR;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_C;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_C1;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_C2;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_C3;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_C4;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_C5;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_C6;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_CLK;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_CO5;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_CO6;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_C_CY;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_C_XOR;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_D;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_D1;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_D2;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_D3;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_D4;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_D5;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_D6;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_DO5;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_DO6;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_D_CY;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_D_XOR;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X104Y136_SR;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_A;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_A1;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_A2;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_A3;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_A4;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_A5;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_A5Q;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_A6;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_AMUX;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_AO5;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_AO6;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_AQ;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_A_CY;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_A_XOR;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_B;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_B1;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_B2;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_B3;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_B4;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_B5;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_B6;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_BMUX;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_BO5;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_BO6;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_BQ;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_B_CY;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_B_XOR;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_C;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_C1;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_C2;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_C3;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_C4;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_C5;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_C6;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_CLK;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_CO5;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_CO6;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_C_CY;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_C_XOR;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_D;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_D1;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_D2;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_D3;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_D4;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_D5;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_D6;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_DO5;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_DO6;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_D_CY;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_D_XOR;
  wire [0:0] CLBLM_L_X70Y136_SLICE_X105Y136_SR;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_A;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_A1;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_A2;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_A3;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_A4;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_A5;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_A6;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_AO5;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_AO6;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_AQ;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_AX;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_A_CY;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_A_XOR;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_B;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_B1;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_B2;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_B3;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_B4;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_B5;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_B6;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_BO5;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_BO6;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_B_CY;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_B_XOR;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_C;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_C1;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_C2;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_C3;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_C4;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_C5;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_C6;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_CLK;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_CO5;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_CO6;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_C_CY;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_C_XOR;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_D;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_D1;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_D2;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_D3;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_D4;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_D5;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_D6;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_DO5;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_DO6;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_D_CY;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_D_XOR;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X104Y98_SR;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_A;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_A1;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_A2;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_A3;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_A4;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_A5;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_A6;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_AO5;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_AO6;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_A_CY;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_A_XOR;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_B;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_B1;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_B2;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_B3;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_B4;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_B5;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_B6;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_BO5;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_BO6;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_B_CY;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_B_XOR;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_C;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_C1;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_C2;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_C3;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_C4;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_C5;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_C6;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_CO5;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_CO6;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_C_CY;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_C_XOR;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_D;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_D1;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_D2;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_D3;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_D4;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_D5;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_D6;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_DO5;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_DO6;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_D_CY;
  wire [0:0] CLBLM_L_X70Y98_SLICE_X105Y98_D_XOR;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_A;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_A1;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_A2;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_A3;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_A4;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_A5;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_A6;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_AO5;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_AO6;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_AQ;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_AX;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_A_CY;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_A_XOR;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_B;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_B1;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_B2;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_B3;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_B4;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_B5;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_B6;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_BO5;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_BO6;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_B_CY;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_B_XOR;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_C;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_C1;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_C2;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_C3;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_C4;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_C5;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_C6;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_CLK;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_CO5;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_CO6;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_C_CY;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_C_XOR;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_D;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_D1;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_D2;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_D3;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_D4;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_D5;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_D6;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_DO5;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_DO6;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_D_CY;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_D_XOR;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X104Y99_SR;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_A;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_A1;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_A2;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_A3;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_A4;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_A5;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_A6;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_AMUX;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_AO5;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_AO6;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_A_CY;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_A_XOR;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_B;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_B1;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_B2;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_B3;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_B4;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_B5;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_B6;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_BO5;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_BO6;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_BQ;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_B_CY;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_B_XOR;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_C;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_C1;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_C2;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_C3;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_C4;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_C5;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_C6;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_CLK;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_CO5;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_CO6;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_CQ;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_C_CY;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_C_XOR;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_D;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_D1;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_D2;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_D3;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_D4;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_D5;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_D6;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_DO5;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_DO6;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_D_CY;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_D_XOR;
  wire [0:0] CLBLM_L_X70Y99_SLICE_X105Y99_SR;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_A;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_A1;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_A2;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_A3;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_A4;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_A5;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_A5Q;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_A6;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_AMUX;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_AO5;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_AO6;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_AQ;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_A_CY;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_A_XOR;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_B;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_B1;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_B2;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_B3;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_B4;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_B5;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_B6;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_BMUX;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_BO5;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_BO6;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_B_CY;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_B_XOR;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_C;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_C1;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_C2;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_C3;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_C4;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_C5;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_C6;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_CLK;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_CMUX;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_CO5;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_CO6;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_C_CY;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_C_XOR;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_D;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_D1;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_D2;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_D3;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_D4;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_D5;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_D6;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_DMUX;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_DO5;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_DO6;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_D_CY;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_D_XOR;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X108Y103_SR;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_A;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_A1;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_A2;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_A3;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_A4;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_A5;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_A6;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_AMUX;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_AO5;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_AO6;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_AQ;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_AX;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_A_CY;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_A_XOR;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_B;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_B1;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_B2;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_B3;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_B4;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_B5;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_B6;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_BO5;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_BO6;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_BQ;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_B_CY;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_B_XOR;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_C;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_C1;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_C2;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_C3;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_C4;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_C5;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_C6;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_CLK;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_CO5;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_CO6;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_C_CY;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_C_XOR;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_D;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_D1;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_D2;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_D3;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_D4;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_D5;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_D6;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_DO5;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_DO6;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_D_CY;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_D_XOR;
  wire [0:0] CLBLM_L_X72Y103_SLICE_X109Y103_SR;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_A;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_A1;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_A2;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_A3;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_A4;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_A5;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_A6;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_AO5;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_AO6;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_AQ;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_A_CY;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_A_XOR;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_B;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_B1;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_B2;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_B3;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_B4;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_B5;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_B6;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_BO5;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_BO6;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_BQ;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_B_CY;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_B_XOR;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_C;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_C1;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_C2;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_C3;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_C4;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_C5;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_C6;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_CLK;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_CO5;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_CO6;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_CQ;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_C_CY;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_C_XOR;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_D;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_D1;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_D2;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_D3;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_D4;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_D5;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_D6;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_DO5;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_DO6;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_DQ;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_D_CY;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_D_XOR;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X108Y104_SR;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_A;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_A1;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_A2;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_A3;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_A4;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_A5;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_A5Q;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_A6;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_AMUX;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_AO5;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_AO6;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_AQ;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_A_CY;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_A_XOR;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_B;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_B1;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_B2;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_B3;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_B4;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_B5;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_B5Q;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_B6;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_BMUX;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_BO5;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_BO6;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_BQ;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_B_CY;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_B_XOR;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_C;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_C1;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_C2;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_C3;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_C4;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_C5;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_C5Q;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_C6;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_CLK;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_CMUX;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_CO5;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_CO6;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_CQ;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_C_CY;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_C_XOR;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_D;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_D1;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_D2;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_D3;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_D4;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_D5;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_D6;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_DO5;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_DO6;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_D_CY;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_D_XOR;
  wire [0:0] CLBLM_L_X72Y104_SLICE_X109Y104_SR;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_A;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_A1;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_A2;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_A3;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_A4;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_A5;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_A5Q;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_A6;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_AMUX;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_AO5;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_AO6;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_AQ;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_A_CY;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_A_XOR;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_B;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_B1;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_B2;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_B3;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_B4;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_B5;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_B6;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_BO5;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_BO6;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_BQ;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_B_CY;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_B_XOR;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_C;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_C1;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_C2;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_C3;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_C4;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_C5;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_C6;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_CLK;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_CO5;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_CO6;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_CQ;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_C_CY;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_C_XOR;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_D;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_D1;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_D2;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_D3;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_D4;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_D5;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_D6;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_DO5;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_DO6;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_DQ;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_D_CY;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_D_XOR;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X108Y105_SR;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_A;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_A1;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_A2;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_A3;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_A4;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_A5;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_A6;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_AO5;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_AO6;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_AQ;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_A_CY;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_A_XOR;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_B;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_B1;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_B2;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_B3;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_B4;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_B5;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_B5Q;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_B6;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_BMUX;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_BO5;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_BO6;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_BQ;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_B_CY;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_B_XOR;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_C;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_C1;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_C2;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_C3;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_C4;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_C5;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_C6;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_CLK;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_CO5;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_CO6;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_C_CY;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_C_XOR;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_D;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_D1;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_D2;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_D3;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_D4;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_D5;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_D6;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_DO5;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_DO6;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_D_CY;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_D_XOR;
  wire [0:0] CLBLM_L_X72Y105_SLICE_X109Y105_SR;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_A;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_A1;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_A2;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_A3;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_A4;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_A5;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_A5Q;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_A6;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_AMUX;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_AO5;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_AO6;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_AQ;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_AX;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_A_CY;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_A_XOR;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_B;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_B1;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_B2;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_B3;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_B4;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_B5;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_B6;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_BMUX;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_BO5;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_BO6;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_B_CY;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_B_XOR;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_C;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_C1;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_C2;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_C3;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_C4;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_C5;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_C6;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_CLK;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_CO5;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_CO6;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_C_CY;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_C_XOR;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_D;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_D1;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_D2;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_D3;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_D4;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_D5;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_D6;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_DMUX;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_DO5;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_DO6;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_D_CY;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_D_XOR;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X108Y106_SR;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_A;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_A1;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_A2;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_A3;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_A4;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_A5;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_A6;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_AO5;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_AO6;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_A_CY;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_A_XOR;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_B;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_B1;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_B2;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_B3;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_B4;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_B5;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_B6;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_BO5;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_BO6;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_B_CY;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_B_XOR;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_C;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_C1;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_C2;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_C3;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_C4;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_C5;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_C6;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_CO5;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_CO6;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_C_CY;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_C_XOR;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_D;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_D1;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_D2;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_D3;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_D4;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_D5;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_D6;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_DO5;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_DO6;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_D_CY;
  wire [0:0] CLBLM_L_X72Y106_SLICE_X109Y106_D_XOR;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_A;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_A1;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_A2;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_A3;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_A4;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_A5;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_A5Q;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_A6;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_AMUX;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_AO5;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_AO6;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_AQ;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_AX;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_A_CY;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_A_XOR;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_B;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_B1;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_B2;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_B3;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_B4;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_B5;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_B6;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_BMUX;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_BO5;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_BO6;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_BQ;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_BX;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_B_CY;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_B_XOR;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_C;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_C1;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_C2;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_C3;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_C4;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_C5;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_C6;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_CLK;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_CO5;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_CO6;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_CQ;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_CX;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_C_CY;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_C_XOR;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_D;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_D1;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_D2;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_D3;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_D4;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_D5;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_D6;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_DO5;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_DO6;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_D_CY;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_D_XOR;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X108Y107_SR;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_A;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_A1;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_A2;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_A3;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_A4;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_A5;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_A5Q;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_A6;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_AMUX;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_AO5;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_AO6;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_AQ;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_AX;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_A_CY;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_A_XOR;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_B;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_B1;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_B2;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_B3;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_B4;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_B5;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_B6;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_BMUX;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_BO5;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_BO6;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_BQ;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_BX;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_B_CY;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_B_XOR;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_C;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_C1;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_C2;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_C3;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_C4;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_C5;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_C6;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_CLK;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_CO5;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_CO6;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_C_CY;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_C_XOR;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_D;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_D1;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_D2;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_D3;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_D4;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_D5;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_D6;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_DO5;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_DO6;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_D_CY;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_D_XOR;
  wire [0:0] CLBLM_L_X72Y107_SLICE_X109Y107_SR;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_A;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_A1;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_A2;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_A3;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_A4;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_A5;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_A6;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_AO5;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_AO6;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_AQ;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_A_CY;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_A_XOR;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_B;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_B1;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_B2;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_B3;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_B4;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_B5;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_B6;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_BMUX;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_BO5;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_BO6;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_B_CY;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_B_XOR;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_C;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_C1;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_C2;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_C3;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_C4;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_C5;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_C6;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_CLK;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_CO5;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_CO6;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_CQ;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_C_CY;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_C_XOR;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_D;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_D1;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_D2;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_D3;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_D4;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_D5;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_D6;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_DO5;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_DO6;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_DQ;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_D_CY;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_D_XOR;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X108Y108_SR;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_A;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_A1;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_A2;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_A3;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_A4;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_A5;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_A5Q;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_A6;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_AMUX;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_AO5;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_AO6;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_AQ;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_A_CY;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_A_XOR;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_B;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_B1;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_B2;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_B3;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_B4;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_B5;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_B6;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_BMUX;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_BO5;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_BO6;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_B_CY;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_B_XOR;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_C;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_C1;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_C2;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_C3;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_C4;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_C5;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_C6;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_CLK;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_CMUX;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_CO5;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_CO6;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_C_CY;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_C_XOR;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_D;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_D1;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_D2;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_D3;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_D4;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_D5;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_D6;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_DO5;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_DO6;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_DQ;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_D_CY;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_D_XOR;
  wire [0:0] CLBLM_L_X72Y108_SLICE_X109Y108_SR;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_A;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_A1;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_A2;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_A3;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_A4;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_A5;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_A6;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_AO5;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_AO6;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_AQ;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_AX;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_A_CY;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_A_XOR;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_B;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_B1;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_B2;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_B3;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_B4;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_B5;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_B6;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_BO5;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_BO6;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_B_CY;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_B_XOR;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_C;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_C1;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_C2;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_C3;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_C4;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_C5;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_C6;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_CLK;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_CO5;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_CO6;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_C_CY;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_C_XOR;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_D;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_D1;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_D2;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_D3;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_D4;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_D5;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_D6;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_DO5;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_DO6;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_D_CY;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_D_XOR;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X108Y109_SR;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_A;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_A1;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_A2;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_A3;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_A4;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_A5;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_A5Q;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_A6;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_AMUX;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_AO5;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_AO6;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_AQ;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_A_CY;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_A_XOR;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_B;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_B1;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_B2;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_B3;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_B4;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_B5;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_B5Q;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_B6;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_BMUX;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_BO5;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_BO6;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_BQ;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_B_CY;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_B_XOR;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_C;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_C1;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_C2;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_C3;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_C4;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_C5;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_C5Q;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_C6;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_CLK;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_CMUX;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_CO5;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_CO6;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_CQ;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_C_CY;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_C_XOR;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_D;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_D1;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_D2;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_D3;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_D4;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_D5;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_D6;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_DO5;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_DO6;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_DQ;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_D_CY;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_D_XOR;
  wire [0:0] CLBLM_L_X72Y109_SLICE_X109Y109_SR;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_A;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_A1;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_A2;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_A3;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_A4;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_A5;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_A6;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_AMUX;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_AO5;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_AO6;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_A_CY;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_A_XOR;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_B;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_B1;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_B2;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_B3;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_B4;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_B5;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_B6;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_BO5;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_BO6;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_BQ;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_B_CY;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_B_XOR;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_C;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_C1;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_C2;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_C3;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_C4;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_C5;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_C5Q;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_C6;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_CLK;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_CMUX;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_CO5;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_CO6;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_CQ;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_C_CY;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_C_XOR;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_D;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_D1;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_D2;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_D3;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_D4;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_D5;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_D6;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_DO5;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_DO6;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_DQ;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_D_CY;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_D_XOR;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X108Y111_SR;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_A;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_A1;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_A2;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_A3;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_A4;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_A5;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_A5Q;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_A6;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_AMUX;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_AO5;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_AO6;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_AQ;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_A_CY;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_A_XOR;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_B;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_B1;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_B2;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_B3;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_B4;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_B5;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_B6;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_BO5;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_BO6;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_BQ;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_BX;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_B_CY;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_B_XOR;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_C;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_C1;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_C2;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_C3;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_C4;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_C5;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_C6;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_CLK;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_CO5;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_CO6;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_CQ;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_CX;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_C_CY;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_C_XOR;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_D;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_D1;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_D2;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_D3;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_D4;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_D5;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_D6;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_DO5;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_DO6;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_D_CY;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_D_XOR;
  wire [0:0] CLBLM_L_X72Y111_SLICE_X109Y111_SR;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_A;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_A1;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_A2;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_A3;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_A4;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_A5;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_A6;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_AO5;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_AO6;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_AQ;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_AX;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_A_CY;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_A_XOR;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_B;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_B1;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_B2;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_B3;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_B4;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_B5;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_B6;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_BO5;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_BO6;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_BQ;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_BX;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_B_CY;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_B_XOR;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_C;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_C1;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_C2;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_C3;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_C4;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_C5;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_C6;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_CLK;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_CO5;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_CO6;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_C_CY;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_C_XOR;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_D;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_D1;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_D2;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_D3;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_D4;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_D5;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_D6;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_DO5;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_DO6;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_D_CY;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_D_XOR;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X108Y113_SR;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_A;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_A1;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_A2;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_A3;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_A4;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_A5;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_A6;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_AO5;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_AO6;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_A_CY;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_A_XOR;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_B;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_B1;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_B2;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_B3;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_B4;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_B5;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_B6;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_BO5;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_BO6;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_B_CY;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_B_XOR;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_C;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_C1;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_C2;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_C3;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_C4;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_C5;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_C6;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_CO5;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_CO6;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_C_CY;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_C_XOR;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_D;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_D1;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_D2;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_D3;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_D4;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_D5;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_D6;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_DO5;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_DO6;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_D_CY;
  wire [0:0] CLBLM_L_X72Y113_SLICE_X109Y113_D_XOR;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_A;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_A1;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_A2;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_A3;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_A4;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_A5;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_A6;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_AO5;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_AO6;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_AQ;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_AX;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_A_CY;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_A_XOR;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_B;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_B1;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_B2;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_B3;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_B4;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_B5;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_B6;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_BO5;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_BO6;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_BQ;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_BX;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_B_CY;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_B_XOR;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_C;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_C1;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_C2;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_C3;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_C4;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_C5;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_C6;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_CE;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_CLK;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_CO5;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_CO6;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_C_CY;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_C_XOR;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_D;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_D1;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_D2;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_D3;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_D4;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_D5;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_D6;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_DO5;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_DO6;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_D_CY;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_D_XOR;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_SR;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_A;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_A1;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_A2;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_A3;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_A4;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_A5;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_A6;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_AO5;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_AO6;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_A_CY;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_A_XOR;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_B;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_B1;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_B2;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_B3;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_B4;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_B5;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_B6;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_BO5;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_BO6;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_B_CY;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_B_XOR;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_C;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_C1;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_C2;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_C3;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_C4;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_C5;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_C6;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_CO5;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_CO6;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_C_CY;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_C_XOR;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_D;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_D1;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_D2;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_D3;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_D4;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_D5;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_D6;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_DO5;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_DO6;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_D_CY;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_D_XOR;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_A;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_A1;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_A2;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_A3;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_A4;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_A5;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_A6;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_AO5;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_AO6;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_AQ;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_AX;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_A_CY;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_A_XOR;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_B;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_B1;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_B2;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_B3;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_B4;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_B5;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_B6;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_BO5;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_BO6;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_BQ;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_BX;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_B_CY;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_B_XOR;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_C;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_C1;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_C2;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_C3;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_C4;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_C5;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_C6;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_CE;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_CLK;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_CO5;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_CO6;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_C_CY;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_C_XOR;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_D;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_D1;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_D2;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_D3;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_D4;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_D5;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_D6;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_DO5;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_DO6;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_D_CY;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_D_XOR;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_SR;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_A;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_A1;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_A2;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_A3;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_A4;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_A5;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_A6;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_AO5;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_AO6;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_A_CY;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_A_XOR;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_B;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_B1;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_B2;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_B3;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_B4;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_B5;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_B6;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_BO5;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_BO6;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_B_CY;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_B_XOR;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_C;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_C1;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_C2;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_C3;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_C4;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_C5;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_C6;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_CO5;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_CO6;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_C_CY;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_C_XOR;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_D;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_D1;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_D2;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_D3;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_D4;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_D5;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_D6;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_DO5;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_DO6;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_D_CY;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_D_XOR;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_A;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_A1;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_A2;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_A3;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_A4;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_A5;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_A5Q;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_A6;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_AMUX;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_AO5;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_AO6;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_AQ;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_A_CY;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_A_XOR;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_B;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_B1;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_B2;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_B3;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_B4;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_B5;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_B5Q;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_B6;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_BMUX;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_BO5;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_BO6;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_BQ;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_B_CY;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_B_XOR;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_C;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_C1;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_C2;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_C3;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_C4;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_C5;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_C5Q;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_C6;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_CLK;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_CMUX;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_CO5;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_CO6;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_CQ;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_C_CY;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_C_XOR;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_D;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_D1;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_D2;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_D3;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_D4;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_D5;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_D5Q;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_D6;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_DMUX;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_DO5;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_DO6;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_DQ;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_D_CY;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_D_XOR;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_SR;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_A;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_A1;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_A2;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_A3;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_A4;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_A5;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_A5Q;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_A6;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_AMUX;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_AO5;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_AO6;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_AQ;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_A_CY;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_A_XOR;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_B;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_B1;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_B2;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_B3;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_B4;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_B5;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_B6;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_BO5;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_BO6;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_BQ;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_B_CY;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_B_XOR;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_C;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_C1;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_C2;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_C3;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_C4;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_C5;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_C6;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_CLK;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_CO5;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_CO6;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_C_CY;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_C_XOR;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_D;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_D1;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_D2;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_D3;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_D4;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_D5;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_D6;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_DO5;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_DO6;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_D_CY;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_D_XOR;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_SR;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_A;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_A1;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_A2;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_A3;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_A4;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_A5;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_A5Q;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_A6;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_AMUX;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_AO5;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_AO6;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_AQ;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_A_CY;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_A_XOR;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_B;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_B1;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_B2;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_B3;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_B4;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_B5;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_B6;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_BO5;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_BO6;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_BQ;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_B_CY;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_B_XOR;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_C;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_C1;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_C2;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_C3;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_C4;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_C5;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_C5Q;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_C6;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_CLK;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_CMUX;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_CO5;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_CO6;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_CQ;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_C_CY;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_C_XOR;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_D;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_D1;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_D2;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_D3;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_D4;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_D5;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_D6;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_DO5;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_DO6;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_D_CY;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_D_XOR;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_SR;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_A;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_A1;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_A2;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_A3;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_A4;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_A5;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_A5Q;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_A6;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_AMUX;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_AO5;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_AO6;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_AQ;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_AX;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_A_CY;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_A_XOR;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_B;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_B1;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_B2;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_B3;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_B4;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_B5;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_B5Q;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_B6;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_BMUX;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_BO5;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_BO6;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_BQ;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_BX;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_B_CY;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_B_XOR;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_C;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_C1;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_C2;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_C3;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_C4;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_C5;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_C6;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_CLK;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_CMUX;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_CO5;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_CO6;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_C_CY;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_C_XOR;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_D;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_D1;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_D2;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_D3;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_D4;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_D5;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_D6;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_DMUX;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_DO5;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_DO6;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_D_CY;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_D_XOR;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_SR;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_A;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_A1;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_A2;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_A3;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_A4;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_A5;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_A5Q;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_A6;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_AMUX;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_AO5;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_AO6;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_AQ;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_A_CY;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_A_XOR;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_B;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_B1;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_B2;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_B3;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_B4;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_B5;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_B6;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_BO5;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_BO6;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_BQ;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_B_CY;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_B_XOR;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_C;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_C1;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_C2;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_C3;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_C4;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_C5;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_C6;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_CLK;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_CO5;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_CO6;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_C_CY;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_C_XOR;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_D;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_D1;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_D2;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_D3;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_D4;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_D5;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_D6;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_DO5;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_DO6;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_D_CY;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_D_XOR;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_SR;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_A;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_A1;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_A2;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_A3;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_A4;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_A5;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_A6;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_AO5;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_AO6;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_A_CY;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_A_XOR;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_B;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_B1;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_B2;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_B3;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_B4;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_B5;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_B6;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_BO5;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_BO6;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_B_CY;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_B_XOR;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_C;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_C1;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_C2;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_C3;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_C4;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_C5;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_C6;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_CO5;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_CO6;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_C_CY;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_C_XOR;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_D;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_D1;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_D2;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_D3;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_D4;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_D5;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_D6;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_DO5;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_DO6;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_D_CY;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_D_XOR;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_A;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_A1;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_A2;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_A3;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_A4;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_A5;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_A5Q;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_A6;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_AMUX;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_AO5;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_AO6;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_AQ;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_AX;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_A_CY;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_A_XOR;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_B;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_B1;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_B2;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_B3;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_B4;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_B5;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_B6;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_BO5;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_BO6;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_BQ;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_BX;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_B_CY;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_B_XOR;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_C;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_C1;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_C2;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_C3;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_C4;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_C5;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_C6;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_CE;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_CLK;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_CO5;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_CO6;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_CQ;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_CX;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_C_CY;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_C_XOR;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_D;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_D1;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_D2;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_D3;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_D4;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_D5;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_D6;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_DO5;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_DO6;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_DQ;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_DX;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_D_CY;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_D_XOR;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_SR;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_A;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_A1;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_A2;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_A3;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_A4;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_A5;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_A5Q;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_A6;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_AMUX;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_AO5;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_AO6;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_AQ;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_A_CY;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_A_XOR;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_B;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_B1;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_B2;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_B3;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_B4;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_B5;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_B6;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_BO5;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_BO6;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_B_CY;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_B_XOR;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_C;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_C1;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_C2;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_C3;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_C4;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_C5;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_C6;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_CLK;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_CO5;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_CO6;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_C_CY;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_C_XOR;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_D;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_D1;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_D2;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_D3;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_D4;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_D5;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_D6;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_DO5;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_DO6;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_D_CY;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_D_XOR;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_SR;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_A;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_A1;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_A2;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_A3;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_A4;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_A5;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_A6;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_AO5;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_AO6;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_AQ;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_AX;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_A_CY;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_A_XOR;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_B;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_B1;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_B2;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_B3;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_B4;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_B5;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_B6;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_BO5;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_BO6;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_BQ;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_BX;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_B_CY;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_B_XOR;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_C;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_C1;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_C2;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_C3;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_C4;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_C5;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_C6;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_CE;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_CLK;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_CO5;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_CO6;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_CQ;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_CX;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_C_CY;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_C_XOR;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_D;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_D1;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_D2;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_D3;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_D4;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_D5;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_D6;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_DO5;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_DO6;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_D_CY;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_D_XOR;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_SR;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_A;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_A1;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_A2;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_A3;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_A4;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_A5;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_A5Q;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_A6;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_AMUX;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_AO5;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_AO6;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_AQ;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_AX;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_A_CY;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_A_XOR;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_B;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_B1;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_B2;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_B3;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_B4;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_B5;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_B6;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_BO5;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_BO6;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_BQ;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_B_CY;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_B_XOR;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_C;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_C1;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_C2;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_C3;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_C4;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_C5;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_C6;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_CLK;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_CMUX;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_CO5;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_CO6;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_C_CY;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_C_XOR;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_D;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_D1;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_D2;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_D3;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_D4;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_D5;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_D6;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_DO5;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_DO6;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_D_CY;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_D_XOR;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_SR;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_A;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_A1;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_A2;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_A3;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_A4;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_A5;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_A5Q;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_A6;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_AMUX;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_AO5;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_AO6;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_AQ;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_AX;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_A_CY;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_A_XOR;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_B;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_B1;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_B2;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_B3;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_B4;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_B5;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_B6;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_BMUX;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_BO5;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_BO6;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_BQ;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_BX;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_B_CY;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_B_XOR;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_C;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_C1;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_C2;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_C3;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_C4;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_C5;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_C6;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_CLK;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_CMUX;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_CO5;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_CO6;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_C_CY;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_C_XOR;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_D;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_D1;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_D2;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_D3;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_D4;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_D5;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_D6;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_DO5;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_DO6;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_D_CY;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_D_XOR;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_SR;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_A;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_A1;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_A2;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_A3;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_A4;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_A5;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_A6;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_AO5;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_AO6;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_AQ;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_A_CY;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_A_XOR;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_B;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_B1;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_B2;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_B3;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_B4;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_B5;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_B6;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_BO5;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_BO6;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_BQ;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_B_CY;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_B_XOR;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_C;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_C1;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_C2;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_C3;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_C4;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_C5;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_C6;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_CLK;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_CO5;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_CO6;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_C_CY;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_C_XOR;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_D;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_D1;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_D2;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_D3;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_D4;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_D5;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_D6;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_DO5;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_DO6;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_D_CY;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_D_XOR;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_SR;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_A;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_A1;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_A2;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_A3;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_A4;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_A5;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_A6;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_AO5;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_AO6;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_AQ;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_A_CY;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_A_XOR;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_B;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_B1;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_B2;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_B3;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_B4;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_B5;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_B6;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_BO5;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_BO6;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_B_CY;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_B_XOR;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_C;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_C1;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_C2;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_C3;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_C4;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_C5;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_C6;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_CLK;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_CO5;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_CO6;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_C_CY;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_C_XOR;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_D;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_D1;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_D2;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_D3;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_D4;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_D5;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_D6;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_DO5;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_DO6;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_D_CY;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_D_XOR;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_SR;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_A;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_A1;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_A2;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_A3;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_A4;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_A5;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_A6;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_AO5;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_AO6;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_AQ;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_A_CY;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_A_XOR;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_B;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_B1;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_B2;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_B3;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_B4;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_B5;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_B6;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_BO5;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_BO6;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_B_CY;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_B_XOR;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_C;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_C1;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_C2;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_C3;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_C4;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_C5;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_C6;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_CLK;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_CO5;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_CO6;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_C_CY;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_C_XOR;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_D;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_D1;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_D2;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_D3;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_D4;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_D5;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_D6;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_DO5;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_DO6;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_D_CY;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_D_XOR;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_SR;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_A;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_A1;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_A2;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_A3;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_A4;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_A5;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_A6;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_AO5;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_AO6;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_AQ;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_A_CY;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_A_XOR;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_B;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_B1;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_B2;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_B3;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_B4;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_B5;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_B6;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_BO5;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_BO6;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_BQ;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_B_CY;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_B_XOR;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_C;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_C1;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_C2;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_C3;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_C4;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_C5;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_C6;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_CLK;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_CO5;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_CO6;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_CQ;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_C_CY;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_C_XOR;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_D;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_D1;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_D2;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_D3;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_D4;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_D5;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_D6;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_DO5;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_DO6;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_D_CY;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_D_XOR;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_SR;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_A;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_A1;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_A2;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_A3;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_A4;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_A5;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_A6;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_AO5;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_AO6;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_AQ;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_A_CY;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_A_XOR;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_B;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_B1;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_B2;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_B3;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_B4;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_B5;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_B6;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_BO5;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_BO6;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_BQ;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_B_CY;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_B_XOR;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_C;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_C1;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_C2;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_C3;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_C4;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_C5;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_C6;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_CLK;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_CO5;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_CO6;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_C_CY;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_C_XOR;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_D;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_D1;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_D2;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_D3;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_D4;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_D5;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_D6;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_DO5;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_DO6;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_D_CY;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_D_XOR;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_SR;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_A;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_A1;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_A2;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_A3;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_A4;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_A5;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_A6;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_AO5;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_AO6;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_AQ;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_A_CY;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_A_XOR;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_B;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_B1;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_B2;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_B3;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_B4;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_B5;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_B6;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_BO5;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_BO6;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_BQ;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_B_CY;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_B_XOR;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_C;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_C1;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_C2;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_C3;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_C4;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_C5;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_C6;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_CLK;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_CO5;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_CO6;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_C_CY;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_C_XOR;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_D;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_D1;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_D2;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_D3;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_D4;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_D5;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_D6;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_DO5;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_DO6;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_D_CY;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_D_XOR;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_SR;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_A;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_A1;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_A2;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_A3;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_A4;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_A5;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_A6;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_AO5;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_AO6;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_AQ;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_A_CY;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_A_XOR;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_B;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_B1;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_B2;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_B3;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_B4;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_B5;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_B6;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_BO5;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_BO6;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_BQ;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_B_CY;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_B_XOR;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_C;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_C1;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_C2;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_C3;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_C4;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_C5;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_C6;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_CLK;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_CO5;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_CO6;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_CQ;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_C_CY;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_C_XOR;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_D;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_D1;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_D2;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_D3;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_D4;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_D5;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_D6;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_DO5;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_DO6;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_D_CY;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_D_XOR;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_SR;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_A;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_A1;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_A2;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_A3;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_A4;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_A5;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_A5Q;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_A6;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_AMUX;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_AO5;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_AO6;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_AQ;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_AX;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_A_CY;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_A_XOR;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_B;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_B1;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_B2;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_B3;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_B4;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_B5;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_B6;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_BMUX;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_BO5;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_BO6;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_B_CY;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_B_XOR;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_C;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_C1;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_C2;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_C3;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_C4;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_C5;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_C6;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_CLK;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_CO5;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_CO6;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_CQ;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_C_CY;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_C_XOR;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_D;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_D1;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_D2;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_D3;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_D4;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_D5;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_D6;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_DO5;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_DO6;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_DQ;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_D_CY;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_D_XOR;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_SR;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_A;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_A1;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_A2;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_A3;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_A4;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_A5;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_A6;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_AO5;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_AO6;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_AQ;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_AX;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_A_CY;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_A_XOR;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_B;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_B1;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_B2;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_B3;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_B4;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_B5;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_B6;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_BO5;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_BO6;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_BQ;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_BX;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_B_CY;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_B_XOR;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_C;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_C1;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_C2;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_C3;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_C4;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_C5;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_C6;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_CE;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_CLK;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_CO5;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_CO6;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_C_CY;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_C_XOR;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_D;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_D1;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_D2;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_D3;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_D4;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_D5;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_D6;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_DO5;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_DO6;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_D_CY;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_D_XOR;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_SR;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_A;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_A1;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_A2;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_A3;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_A4;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_A5;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_A5Q;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_A6;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_AMUX;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_AO5;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_AO6;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_AQ;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_AX;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_A_CY;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_A_XOR;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_B;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_B1;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_B2;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_B3;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_B4;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_B5;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_B6;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_BMUX;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_BO5;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_BO6;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_B_CY;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_B_XOR;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_C;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_C1;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_C2;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_C3;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_C4;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_C5;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_C6;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_CLK;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_CO5;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_CO6;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_CQ;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_C_CY;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_C_XOR;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_D;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_D1;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_D2;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_D3;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_D4;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_D5;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_D6;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_DO5;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_DO6;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_DQ;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_D_CY;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_D_XOR;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_SR;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_A;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_A1;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_A2;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_A3;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_A4;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_A5;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_A6;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_AO5;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_AO6;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_AQ;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_A_CY;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_A_XOR;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_B;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_B1;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_B2;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_B3;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_B4;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_B5;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_B6;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_BO5;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_BO6;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_B_CY;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_B_XOR;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_C;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_C1;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_C2;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_C3;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_C4;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_C5;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_C6;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_CLK;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_CO5;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_CO6;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_C_CY;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_C_XOR;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_D;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_D1;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_D2;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_D3;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_D4;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_D5;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_D6;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_DO5;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_DO6;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_D_CY;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_D_XOR;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_SR;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_A;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_A1;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_A2;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_A3;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_A4;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_A5;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_A6;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_AMUX;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_AO5;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_AO6;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_AQ;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_A_CY;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_A_XOR;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_B;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_B1;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_B2;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_B3;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_B4;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_B5;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_B6;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_BO5;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_BO6;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_BQ;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_B_CY;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_B_XOR;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_C;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_C1;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_C2;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_C3;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_C4;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_C5;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_C6;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_CLK;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_CO5;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_CO6;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_C_CY;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_C_XOR;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_D;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_D1;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_D2;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_D3;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_D4;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_D5;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_D6;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_DO5;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_DO6;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_D_CY;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_D_XOR;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_SR;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_A;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_A1;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_A2;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_A3;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_A4;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_A5;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_A6;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_AO5;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_AO6;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_A_CY;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_A_XOR;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_B;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_B1;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_B2;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_B3;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_B4;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_B5;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_B6;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_BO5;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_BO6;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_B_CY;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_B_XOR;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_C;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_C1;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_C2;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_C3;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_C4;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_C5;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_C6;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_CO5;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_CO6;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_C_CY;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_C_XOR;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_D;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_D1;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_D2;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_D3;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_D4;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_D5;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_D6;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_DO5;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_DO6;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_D_CY;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_D_XOR;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_A;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_A1;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_A2;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_A3;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_A4;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_A5;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_A6;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_AO5;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_AO6;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_AQ;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_A_CY;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_A_XOR;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_B;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_B1;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_B2;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_B3;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_B4;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_B5;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_B6;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_BO5;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_BO6;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_BQ;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_B_CY;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_B_XOR;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_C;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_C1;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_C2;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_C3;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_C4;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_C5;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_C6;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_CLK;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_CO5;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_CO6;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_CQ;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_C_CY;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_C_XOR;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_D;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_D1;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_D2;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_D3;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_D4;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_D5;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_D6;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_DO5;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_DO6;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_DQ;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_D_CY;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_D_XOR;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X108Y130_SR;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_A;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_A1;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_A2;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_A3;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_A4;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_A5;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_A6;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_AO5;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_AO6;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_AQ;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_A_CY;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_A_XOR;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_B;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_B1;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_B2;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_B3;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_B4;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_B5;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_B6;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_BO5;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_BO6;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_BQ;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_B_CY;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_B_XOR;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_C;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_C1;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_C2;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_C3;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_C4;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_C5;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_C6;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_CLK;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_CO5;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_CO6;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_CQ;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_C_CY;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_C_XOR;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_D;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_D1;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_D2;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_D3;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_D4;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_D5;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_D6;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_DO5;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_DO6;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_D_CY;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_D_XOR;
  wire [0:0] CLBLM_L_X72Y130_SLICE_X109Y130_SR;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_A;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_A1;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_A2;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_A3;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_A4;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_A5;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_A5Q;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_A6;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_AMUX;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_AO5;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_AO6;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_AQ;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_A_CY;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_A_XOR;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_B;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_B1;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_B2;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_B3;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_B4;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_B5;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_B6;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_BO5;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_BO6;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_BQ;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_B_CY;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_B_XOR;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_C;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_C1;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_C2;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_C3;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_C4;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_C5;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_C6;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_CLK;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_CO5;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_CO6;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_CQ;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_C_CY;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_C_XOR;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_D;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_D1;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_D2;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_D3;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_D4;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_D5;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_D6;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_DMUX;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_DO5;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_DO6;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_D_CY;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_D_XOR;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_SR;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_A;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_A1;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_A2;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_A3;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_A4;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_A5;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_A6;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_AMUX;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_AO5;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_AO6;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_A_CY;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_A_XOR;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_B;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_B1;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_B2;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_B3;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_B4;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_B5;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_B6;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_BO5;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_BO6;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_BQ;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_B_CY;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_B_XOR;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_C;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_C1;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_C2;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_C3;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_C4;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_C5;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_C6;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_CLK;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_CO5;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_CO6;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_CQ;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_C_CY;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_C_XOR;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_D;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_D1;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_D2;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_D3;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_D4;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_D5;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_D6;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_DO5;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_DO6;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_DQ;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_D_CY;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_D_XOR;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_SR;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_A;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_A1;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_A2;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_A3;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_A4;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_A5;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_A6;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_AO5;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_AO6;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_AQ;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_A_CY;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_A_XOR;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_B;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_B1;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_B2;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_B3;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_B4;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_B5;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_B6;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_BO5;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_BO6;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_BQ;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_B_CY;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_B_XOR;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_C;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_C1;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_C2;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_C3;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_C4;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_C5;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_C6;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_CLK;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_CO5;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_CO6;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_CQ;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_C_CY;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_C_XOR;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_D;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_D1;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_D2;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_D3;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_D4;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_D5;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_D6;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_DO5;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_DO6;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_DQ;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_D_CY;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_D_XOR;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X108Y132_SR;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_A;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_A1;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_A2;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_A3;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_A4;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_A5;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_A6;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_AO5;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_AO6;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_AQ;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_AX;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_A_CY;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_A_XOR;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_B;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_B1;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_B2;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_B3;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_B4;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_B5;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_B6;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_BO5;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_BO6;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_B_CY;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_B_XOR;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_C;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_C1;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_C2;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_C3;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_C4;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_C5;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_C6;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_CE;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_CLK;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_CMUX;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_CO5;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_CO6;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_C_CY;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_C_XOR;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_D;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_D1;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_D2;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_D3;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_D4;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_D5;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_D6;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_DO5;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_DO6;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_D_CY;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_D_XOR;
  wire [0:0] CLBLM_L_X72Y132_SLICE_X109Y132_SR;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_A;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_A1;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_A2;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_A3;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_A4;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_A5;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_A5Q;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_A6;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_AMUX;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_AO5;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_AO6;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_AQ;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_A_CY;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_A_XOR;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_B;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_B1;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_B2;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_B3;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_B4;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_B5;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_B6;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_BMUX;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_BO5;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_BO6;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_B_CY;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_B_XOR;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_C;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_C1;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_C2;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_C3;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_C4;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_C5;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_C6;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_CLK;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_CO5;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_CO6;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_CQ;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_C_CY;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_C_XOR;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_D;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_D1;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_D2;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_D3;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_D4;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_D5;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_D6;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_DMUX;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_DO5;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_DO6;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_D_CY;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_D_XOR;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X108Y133_SR;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_A;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_A1;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_A2;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_A3;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_A4;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_A5;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_A6;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_AMUX;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_AO5;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_AO6;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_A_CY;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_A_XOR;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_B;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_B1;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_B2;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_B3;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_B4;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_B5;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_B6;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_BO5;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_BO6;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_BQ;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_B_CY;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_B_XOR;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_C;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_C1;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_C2;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_C3;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_C4;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_C5;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_C6;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_CLK;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_CO5;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_CO6;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_C_CY;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_C_XOR;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_D;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_D1;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_D2;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_D3;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_D4;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_D5;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_D6;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_DO5;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_DO6;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_D_CY;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_D_XOR;
  wire [0:0] CLBLM_L_X72Y133_SLICE_X109Y133_SR;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_A;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_A1;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_A2;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_A3;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_A4;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_A5;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_A6;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_AO5;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_AO6;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_AQ;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_A_CY;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_A_XOR;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_B;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_B1;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_B2;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_B3;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_B4;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_B5;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_B6;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_BO5;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_BO6;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_B_CY;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_B_XOR;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_C;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_C1;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_C2;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_C3;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_C4;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_C5;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_C6;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_CLK;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_CO5;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_CO6;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_C_CY;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_C_XOR;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_D;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_D1;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_D2;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_D3;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_D4;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_D5;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_D6;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_DO5;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_DO6;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_D_CY;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_D_XOR;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X108Y134_SR;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_A;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_A1;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_A2;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_A3;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_A4;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_A5;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_A6;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_AMUX;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_AO5;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_AO6;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_A_CY;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_A_XOR;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_B;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_B1;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_B2;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_B3;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_B4;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_B5;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_B6;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_BMUX;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_BO5;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_BO6;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_B_CY;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_B_XOR;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_C;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_C1;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_C2;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_C3;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_C4;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_C5;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_C6;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_CO5;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_CO6;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_C_CY;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_C_XOR;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_D;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_D1;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_D2;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_D3;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_D4;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_D5;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_D6;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_DO5;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_DO6;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_D_CY;
  wire [0:0] CLBLM_L_X72Y134_SLICE_X109Y134_D_XOR;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_A;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_A1;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_A2;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_A3;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_A4;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_A5;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_A5Q;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_A6;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_AMUX;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_AO5;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_AO6;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_AQ;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_AX;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_A_CY;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_A_XOR;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_B;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_B1;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_B2;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_B3;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_B4;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_B5;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_B5Q;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_B6;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_BMUX;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_BO5;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_BO6;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_BQ;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_BX;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_B_CY;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_B_XOR;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_C;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_C1;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_C2;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_C3;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_C4;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_C5;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_C6;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_CLK;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_CO5;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_CO6;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_C_CY;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_C_XOR;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_D;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_D1;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_D2;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_D3;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_D4;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_D5;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_D6;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_DO5;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_DO6;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_D_CY;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_D_XOR;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X108Y98_SR;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_A;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_A1;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_A2;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_A3;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_A4;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_A5;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_A6;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_AO5;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_AO6;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_A_CY;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_A_XOR;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_B;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_B1;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_B2;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_B3;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_B4;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_B5;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_B6;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_BO5;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_BO6;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_B_CY;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_B_XOR;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_C;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_C1;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_C2;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_C3;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_C4;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_C5;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_C6;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_CO5;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_CO6;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_C_CY;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_C_XOR;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_D;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_D1;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_D2;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_D3;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_D4;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_D5;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_D6;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_DO5;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_DO6;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_D_CY;
  wire [0:0] CLBLM_L_X72Y98_SLICE_X109Y98_D_XOR;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_A;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_A1;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_A2;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_A3;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_A4;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_A5;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_A6;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_AO5;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_AO6;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_AQ;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_A_CY;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_A_XOR;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_B;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_B1;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_B2;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_B3;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_B4;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_B5;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_B6;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_BO5;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_BO6;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_B_CY;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_B_XOR;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_C;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_C1;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_C2;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_C3;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_C4;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_C5;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_C6;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_CLK;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_CO5;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_CO6;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_C_CY;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_C_XOR;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_D;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_D1;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_D2;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_D3;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_D4;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_D5;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_D6;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_DO5;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_DO6;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_D_CY;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_D_XOR;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X112Y102_SR;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_A;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_A1;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_A2;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_A3;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_A4;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_A5;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_A6;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_AO5;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_AO6;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_A_CY;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_A_XOR;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_B;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_B1;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_B2;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_B3;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_B4;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_B5;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_B6;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_BO5;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_BO6;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_B_CY;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_B_XOR;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_C;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_C1;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_C2;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_C3;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_C4;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_C5;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_C6;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_CO5;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_CO6;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_C_CY;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_C_XOR;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_D;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_D1;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_D2;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_D3;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_D4;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_D5;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_D6;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_DO5;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_DO6;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_D_CY;
  wire [0:0] CLBLM_L_X74Y102_SLICE_X113Y102_D_XOR;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_A;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_A1;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_A2;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_A3;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_A4;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_A5;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_A6;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_AO5;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_AO6;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_AQ;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_A_CY;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_A_XOR;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_B;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_B1;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_B2;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_B3;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_B4;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_B5;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_B6;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_BO5;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_BO6;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_BQ;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_B_CY;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_B_XOR;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_C;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_C1;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_C2;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_C3;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_C4;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_C5;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_C6;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_CLK;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_CO5;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_CO6;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_C_CY;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_C_XOR;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_D;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_D1;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_D2;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_D3;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_D4;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_D5;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_D6;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_DMUX;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_DO5;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_DO6;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_D_CY;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_D_XOR;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X112Y103_SR;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_A;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_A1;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_A2;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_A3;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_A4;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_A5;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_A6;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_AO5;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_AO6;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_AQ;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_A_CY;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_A_XOR;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_B;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_B1;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_B2;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_B3;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_B4;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_B5;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_B6;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_BO5;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_BO6;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_BQ;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_B_CY;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_B_XOR;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_C;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_C1;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_C2;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_C3;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_C4;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_C5;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_C6;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_CLK;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_CO5;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_CO6;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_C_CY;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_C_XOR;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_D;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_D1;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_D2;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_D3;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_D4;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_D5;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_D6;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_DO5;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_DO6;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_D_CY;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_D_XOR;
  wire [0:0] CLBLM_L_X74Y103_SLICE_X113Y103_SR;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_A;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_A1;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_A2;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_A3;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_A4;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_A5;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_A6;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_AO5;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_AO6;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_AQ;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_A_CY;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_A_XOR;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_B;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_B1;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_B2;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_B3;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_B4;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_B5;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_B6;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_BO5;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_BO6;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_BQ;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_B_CY;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_B_XOR;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_C;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_C1;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_C2;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_C3;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_C4;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_C5;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_C6;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_CLK;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_CO5;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_CO6;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_CQ;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_C_CY;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_C_XOR;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_D;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_D1;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_D2;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_D3;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_D4;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_D5;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_D6;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_DO5;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_DO6;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_D_CY;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_D_XOR;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X112Y104_SR;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_A;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_A1;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_A2;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_A3;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_A4;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_A5;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_A6;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_AO5;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_AO6;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_A_CY;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_A_XOR;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_B;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_B1;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_B2;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_B3;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_B4;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_B5;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_B6;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_BO5;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_BO6;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_B_CY;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_B_XOR;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_C;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_C1;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_C2;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_C3;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_C4;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_C5;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_C6;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_CO5;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_CO6;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_C_CY;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_C_XOR;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_D;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_D1;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_D2;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_D3;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_D4;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_D5;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_D6;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_DO5;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_DO6;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_D_CY;
  wire [0:0] CLBLM_L_X74Y104_SLICE_X113Y104_D_XOR;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_A;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_A1;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_A2;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_A3;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_A4;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_A5;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_A6;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_AO5;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_AO6;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_AQ;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_A_CY;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_A_XOR;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_B;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_B1;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_B2;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_B3;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_B4;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_B5;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_B6;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_BO5;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_BO6;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_BQ;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_B_CY;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_B_XOR;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_C;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_C1;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_C2;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_C3;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_C4;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_C5;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_C6;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_CLK;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_CO5;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_CO6;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_CQ;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_C_CY;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_C_XOR;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_D;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_D1;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_D2;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_D3;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_D4;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_D5;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_D6;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_DO5;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_DO6;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_DQ;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_D_CY;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_D_XOR;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X112Y107_SR;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_A;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_A1;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_A2;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_A3;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_A4;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_A5;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_A6;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_AO5;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_AO6;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_AQ;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_A_CY;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_A_XOR;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_B;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_B1;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_B2;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_B3;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_B4;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_B5;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_B6;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_BO5;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_BO6;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_B_CY;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_B_XOR;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_C;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_C1;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_C2;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_C3;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_C4;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_C5;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_C6;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_CLK;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_CO5;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_CO6;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_C_CY;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_C_XOR;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_D;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_D1;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_D2;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_D3;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_D4;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_D5;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_D6;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_DO5;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_DO6;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_D_CY;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_D_XOR;
  wire [0:0] CLBLM_L_X74Y107_SLICE_X113Y107_SR;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_A;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_A1;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_A2;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_A3;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_A4;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_A5;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_A6;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_AO5;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_AO6;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_A_CY;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_A_XOR;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_B;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_B1;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_B2;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_B3;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_B4;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_B5;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_B6;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_BO5;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_BO6;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_B_CY;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_B_XOR;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_C;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_C1;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_C2;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_C3;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_C4;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_C5;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_C6;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_CO5;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_CO6;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_C_CY;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_C_XOR;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_D;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_D1;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_D2;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_D3;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_D4;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_D5;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_D6;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_DO5;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_DO6;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_D_CY;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X112Y109_D_XOR;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_A;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_A1;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_A2;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_A3;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_A4;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_A5;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_A5Q;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_A6;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_AMUX;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_AO5;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_AO6;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_AQ;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_A_CY;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_A_XOR;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_B;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_B1;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_B2;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_B3;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_B4;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_B5;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_B6;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_BO5;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_BO6;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_B_CY;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_B_XOR;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_C;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_C1;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_C2;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_C3;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_C4;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_C5;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_C6;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_CLK;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_CO5;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_CO6;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_C_CY;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_C_XOR;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_D;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_D1;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_D2;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_D3;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_D4;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_D5;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_D6;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_DO5;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_DO6;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_D_CY;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_D_XOR;
  wire [0:0] CLBLM_L_X74Y109_SLICE_X113Y109_SR;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_A;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_A1;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_A2;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_A3;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_A4;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_A5;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_A6;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_AO5;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_AO6;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_AQ;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_AX;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_A_CY;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_A_XOR;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_B;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_B1;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_B2;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_B3;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_B4;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_B5;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_B6;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_BO5;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_BO6;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_BQ;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_BX;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_B_CY;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_B_XOR;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_C;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_C1;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_C2;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_C3;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_C4;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_C5;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_C6;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_CE;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_CLK;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_CO5;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_CO6;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_C_CY;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_C_XOR;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_D;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_D1;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_D2;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_D3;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_D4;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_D5;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_D6;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_DO5;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_DO6;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_D_CY;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_D_XOR;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_SR;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_A;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_A1;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_A2;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_A3;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_A4;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_A5;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_A6;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_AO5;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_AO6;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_A_CY;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_A_XOR;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_B;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_B1;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_B2;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_B3;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_B4;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_B5;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_B6;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_BO5;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_BO6;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_B_CY;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_B_XOR;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_C;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_C1;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_C2;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_C3;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_C4;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_C5;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_C6;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_CO5;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_CO6;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_C_CY;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_C_XOR;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_D;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_D1;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_D2;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_D3;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_D4;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_D5;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_D6;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_DO5;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_DO6;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_D_CY;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_D_XOR;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_A;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_A1;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_A2;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_A3;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_A4;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_A5;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_A6;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_AO5;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_AO6;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_AQ;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_A_CY;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_A_XOR;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_B;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_B1;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_B2;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_B3;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_B4;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_B5;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_B6;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_BMUX;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_BO5;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_BO6;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_B_CY;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_B_XOR;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_C;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_C1;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_C2;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_C3;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_C4;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_C5;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_C6;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_CLK;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_CO5;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_CO6;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_CQ;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_C_CY;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_C_XOR;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_D;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_D1;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_D2;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_D3;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_D4;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_D5;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_D6;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_DO5;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_DO6;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_D_CY;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_D_XOR;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_SR;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_A;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_A1;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_A2;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_A3;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_A4;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_A5;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_A6;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_AO5;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_AO6;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_A_CY;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_A_XOR;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_B;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_B1;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_B2;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_B3;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_B4;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_B5;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_B6;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_BO5;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_BO6;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_B_CY;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_B_XOR;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_C;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_C1;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_C2;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_C3;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_C4;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_C5;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_C6;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_CO5;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_CO6;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_C_CY;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_C_XOR;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_D;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_D1;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_D2;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_D3;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_D4;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_D5;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_D6;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_DO5;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_DO6;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_D_CY;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_D_XOR;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_A;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_A1;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_A2;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_A3;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_A4;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_A5;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_A6;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_AO5;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_AO6;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_AQ;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_A_CY;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_A_XOR;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_B;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_B1;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_B2;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_B3;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_B4;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_B5;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_B6;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_BMUX;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_BO5;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_BO6;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_B_CY;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_B_XOR;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_C;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_C1;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_C2;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_C3;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_C4;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_C5;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_C6;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_CLK;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_CO5;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_CO6;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_CQ;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_C_CY;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_C_XOR;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_D;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_D1;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_D2;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_D3;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_D4;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_D5;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_D6;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_DO5;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_DO6;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_DQ;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_D_CY;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_D_XOR;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_SR;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_A;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_A1;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_A2;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_A3;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_A4;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_A5;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_A6;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_AMUX;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_AO5;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_AO6;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_A_CY;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_A_XOR;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_B;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_B1;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_B2;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_B3;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_B4;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_B5;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_B6;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_BO5;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_BO6;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_B_CY;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_B_XOR;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_C;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_C1;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_C2;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_C3;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_C4;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_C5;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_C6;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_CO5;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_CO6;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_C_CY;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_C_XOR;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_D;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_D1;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_D2;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_D3;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_D4;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_D5;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_D6;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_DO5;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_DO6;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_D_CY;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_D_XOR;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_A;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_A1;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_A2;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_A3;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_A4;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_A5;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_A6;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_AO5;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_AO6;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_A_CY;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_A_XOR;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_B;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_B1;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_B2;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_B3;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_B4;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_B5;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_B6;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_BO5;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_BO6;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_B_CY;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_B_XOR;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_C;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_C1;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_C2;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_C3;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_C4;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_C5;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_C6;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_CO5;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_CO6;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_C_CY;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_C_XOR;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_D;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_D1;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_D2;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_D3;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_D4;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_D5;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_D6;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_DO5;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_DO6;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_D_CY;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_D_XOR;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_A;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_A1;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_A2;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_A3;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_A4;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_A5;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_A6;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_AO5;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_AO6;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_A_CY;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_A_XOR;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_B;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_B1;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_B2;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_B3;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_B4;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_B5;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_B6;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_BO5;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_BO6;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_B_CY;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_B_XOR;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_C;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_C1;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_C2;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_C3;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_C4;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_C5;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_C6;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_CO5;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_CO6;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_C_CY;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_C_XOR;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_D;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_D1;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_D2;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_D3;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_D4;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_D5;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_D6;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_DO5;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_DO6;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_D_CY;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_D_XOR;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_A;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_A1;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_A2;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_A3;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_A4;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_A5;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_A6;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_AO5;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_AO6;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_A_CY;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_A_XOR;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_B;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_B1;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_B2;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_B3;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_B4;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_B5;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_B6;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_BO5;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_BO6;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_B_CY;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_B_XOR;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_C;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_C1;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_C2;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_C3;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_C4;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_C5;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_C6;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_CO5;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_CO6;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_C_CY;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_C_XOR;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_D;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_D1;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_D2;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_D3;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_D4;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_D5;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_D6;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_DO5;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_DO6;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_D_CY;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_D_XOR;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_A;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_A1;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_A2;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_A3;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_A4;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_A5;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_A5Q;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_A6;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_AMUX;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_AO5;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_AO6;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_AQ;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_A_CY;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_A_XOR;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_B;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_B1;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_B2;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_B3;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_B4;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_B5;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_B5Q;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_B6;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_BMUX;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_BO5;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_BO6;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_BQ;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_B_CY;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_B_XOR;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_C;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_C1;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_C2;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_C3;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_C4;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_C5;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_C6;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_CLK;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_CO5;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_CO6;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_C_CY;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_C_XOR;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_D;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_D1;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_D2;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_D3;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_D4;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_D5;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_D6;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_DO5;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_DO6;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_D_CY;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_D_XOR;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_SR;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_A;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_A1;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_A2;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_A3;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_A4;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_A5;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_A5Q;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_A6;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_AMUX;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_AO5;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_AO6;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_AQ;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_A_CY;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_A_XOR;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_B;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_B1;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_B2;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_B3;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_B4;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_B5;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_B6;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_BO5;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_BO6;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_BQ;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_B_CY;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_B_XOR;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_C;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_C1;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_C2;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_C3;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_C4;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_C5;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_C6;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_CLK;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_CO5;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_CO6;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_C_CY;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_C_XOR;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_D;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_D1;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_D2;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_D3;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_D4;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_D5;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_D6;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_DO5;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_DO6;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_D_CY;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_D_XOR;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X112Y122_SR;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_A;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_A1;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_A2;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_A3;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_A4;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_A5;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_A6;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_AO5;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_AO6;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_AQ;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_A_CY;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_A_XOR;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_B;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_B1;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_B2;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_B3;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_B4;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_B5;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_B6;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_BO5;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_BO6;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_B_CY;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_B_XOR;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_C;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_C1;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_C2;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_C3;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_C4;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_C5;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_C6;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_CLK;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_CO5;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_CO6;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_C_CY;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_C_XOR;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_D;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_D1;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_D2;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_D3;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_D4;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_D5;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_D6;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_DO5;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_DO6;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_D_CY;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_D_XOR;
  wire [0:0] CLBLM_L_X74Y122_SLICE_X113Y122_SR;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_A;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_A1;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_A2;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_A3;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_A4;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_A5;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_A6;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_AO5;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_AO6;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_AQ;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_A_CY;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_A_XOR;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_B;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_B1;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_B2;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_B3;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_B4;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_B5;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_B5Q;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_B6;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_BMUX;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_BO5;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_BO6;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_BQ;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_B_CY;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_B_XOR;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_C;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_C1;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_C2;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_C3;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_C4;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_C5;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_C6;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_CLK;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_CO5;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_CO6;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_C_CY;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_C_XOR;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_D;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_D1;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_D2;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_D3;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_D4;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_D5;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_D6;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_DO5;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_DO6;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_D_CY;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_D_XOR;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_SR;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_A;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_A1;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_A2;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_A3;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_A4;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_A5;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_A5Q;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_A6;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_AMUX;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_AO5;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_AO6;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_AQ;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_AX;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_A_CY;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_A_XOR;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_B;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_B1;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_B2;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_B3;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_B4;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_B5;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_B6;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_BO5;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_BO6;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_BQ;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_B_CY;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_B_XOR;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_C;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_C1;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_C2;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_C3;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_C4;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_C5;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_C6;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_CLK;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_CMUX;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_CO5;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_CO6;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_C_CY;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_C_XOR;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_D;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_D1;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_D2;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_D3;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_D4;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_D5;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_D6;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_DO5;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_DO6;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_DQ;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_D_CY;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_D_XOR;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_SR;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_A;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_A1;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_A2;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_A3;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_A4;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_A5;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_A6;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_AO5;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_AO6;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_AQ;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_AX;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_A_CY;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_A_XOR;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_B;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_B1;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_B2;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_B3;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_B4;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_B5;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_B6;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_BO5;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_BO6;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_B_CY;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_B_XOR;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_C;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_C1;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_C2;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_C3;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_C4;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_C5;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_C6;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_CE;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_CLK;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_CO5;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_CO6;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_C_CY;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_C_XOR;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_D;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_D1;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_D2;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_D3;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_D4;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_D5;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_D6;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_DO5;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_DO6;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_D_CY;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_D_XOR;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_SR;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_A;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_A1;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_A2;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_A3;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_A4;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_A5;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_A6;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_AO5;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_AO6;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_A_CY;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_A_XOR;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_B;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_B1;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_B2;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_B3;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_B4;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_B5;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_B6;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_BO5;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_BO6;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_B_CY;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_B_XOR;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_C;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_C1;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_C2;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_C3;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_C4;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_C5;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_C6;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_CO5;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_CO6;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_C_CY;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_C_XOR;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_D;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_D1;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_D2;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_D3;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_D4;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_D5;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_D6;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_DO5;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_DO6;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_D_CY;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_D_XOR;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_A;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_A1;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_A2;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_A3;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_A4;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_A5;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_A5Q;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_A6;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_AMUX;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_AO5;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_AO6;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_AQ;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_AX;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_A_CY;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_A_XOR;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_B;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_B1;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_B2;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_B3;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_B4;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_B5;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_B6;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_BMUX;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_BO5;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_BO6;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_B_CY;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_B_XOR;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_C;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_C1;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_C2;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_C3;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_C4;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_C5;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_C6;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_CLK;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_CMUX;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_CO5;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_CO6;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_C_CY;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_C_XOR;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_D;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_D1;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_D2;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_D3;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_D4;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_D5;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_D6;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_DO5;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_DO6;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_DQ;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_D_CY;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_D_XOR;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_SR;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_A;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_A1;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_A2;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_A3;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_A4;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_A5;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_A5Q;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_A6;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_AMUX;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_AO5;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_AO6;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_AQ;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_A_CY;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_A_XOR;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_B;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_B1;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_B2;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_B3;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_B4;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_B5;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_B6;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_BO5;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_BO6;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_BQ;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_B_CY;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_B_XOR;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_C;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_C1;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_C2;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_C3;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_C4;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_C5;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_C6;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_CLK;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_CO5;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_CO6;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_CQ;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_C_CY;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_C_XOR;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_D;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_D1;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_D2;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_D3;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_D4;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_D5;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_D6;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_DO5;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_DO6;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_D_CY;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_D_XOR;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_SR;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_A;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_A1;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_A2;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_A3;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_A4;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_A5;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_A6;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_AMUX;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_AO5;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_AO6;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_AQ;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_AX;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_A_CY;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_A_XOR;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_B;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_B1;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_B2;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_B3;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_B4;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_B5;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_B6;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_BO5;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_BO6;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_BQ;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_BX;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_B_CY;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_B_XOR;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_C;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_C1;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_C2;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_C3;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_C4;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_C5;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_C6;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_CE;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_CLK;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_CMUX;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_CO5;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_CO6;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_C_CY;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_C_XOR;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_D;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_D1;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_D2;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_D3;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_D4;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_D5;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_D6;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_DO5;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_DO6;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_D_CY;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_D_XOR;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_SR;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_A;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_A1;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_A2;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_A3;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_A4;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_A5;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_A5Q;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_A6;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_AMUX;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_AO5;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_AO6;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_AQ;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_AX;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_A_CY;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_A_XOR;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_B;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_B1;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_B2;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_B3;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_B4;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_B5;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_B6;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_BMUX;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_BO5;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_BO6;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_B_CY;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_B_XOR;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_C;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_C1;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_C2;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_C3;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_C4;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_C5;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_C6;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_CLK;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_CO5;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_CO6;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_CQ;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_C_CY;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_C_XOR;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_D;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_D1;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_D2;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_D3;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_D4;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_D5;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_D6;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_DO5;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_DO6;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_D_CY;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_D_XOR;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_SR;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_A;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_A1;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_A2;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_A3;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_A4;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_A5;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_A6;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_AO5;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_AO6;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_AQ;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_A_CY;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_A_XOR;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_B;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_B1;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_B2;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_B3;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_B4;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_B5;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_B6;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_BO5;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_BO6;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_BQ;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_B_CY;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_B_XOR;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_C;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_C1;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_C2;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_C3;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_C4;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_C5;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_C6;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_CLK;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_CO5;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_CO6;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_CQ;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_C_CY;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_C_XOR;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_D;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_D1;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_D2;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_D3;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_D4;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_D5;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_D6;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_DO5;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_DO6;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_DQ;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_D_CY;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_D_XOR;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_SR;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_A;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_A1;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_A2;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_A3;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_A4;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_A5;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_A6;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_AMUX;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_AO5;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_AO6;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_A_CY;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_A_XOR;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_B;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_B1;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_B2;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_B3;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_B4;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_B5;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_B6;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_BMUX;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_BO5;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_BO6;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_B_CY;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_B_XOR;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_C;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_C1;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_C2;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_C3;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_C4;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_C5;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_C6;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_CLK;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_CO5;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_CO6;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_CQ;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_C_CY;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_C_XOR;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_D;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_D1;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_D2;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_D3;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_D4;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_D5;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_D6;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_DO5;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_DO6;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_D_CY;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_D_XOR;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_SR;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_A;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_A1;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_A2;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_A3;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_A4;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_A5;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_A5Q;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_A6;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_AMUX;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_AO5;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_AO6;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_AQ;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_A_CY;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_A_XOR;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_B;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_B1;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_B2;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_B3;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_B4;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_B5;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_B6;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_BO5;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_BO6;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_BQ;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_BX;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_B_CY;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_B_XOR;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_C;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_C1;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_C2;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_C3;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_C4;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_C5;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_C6;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_CLK;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_CO5;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_CO6;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_C_CY;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_C_XOR;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_D;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_D1;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_D2;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_D3;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_D4;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_D5;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_D6;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_DO5;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_DO6;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_D_CY;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_D_XOR;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_SR;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_A;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_A1;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_A2;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_A3;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_A4;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_A5;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_A6;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_AO5;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_AO6;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_AQ;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_A_CY;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_A_XOR;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_B;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_B1;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_B2;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_B3;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_B4;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_B5;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_B6;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_BMUX;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_BO5;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_BO6;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_B_CY;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_B_XOR;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_C;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_C1;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_C2;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_C3;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_C4;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_C5;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_C6;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_CLK;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_CO5;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_CO6;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_C_CY;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_C_XOR;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_D;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_D1;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_D2;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_D3;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_D4;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_D5;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_D6;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_DO5;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_DO6;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_D_CY;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_D_XOR;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_SR;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_A;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_A1;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_A2;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_A3;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_A4;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_A5;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_A6;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_AO5;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_AO6;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_AQ;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_AX;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_A_CY;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_A_XOR;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_B;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_B1;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_B2;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_B3;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_B4;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_B5;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_B6;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_BO5;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_BO6;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_B_CY;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_B_XOR;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_C;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_C1;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_C2;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_C3;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_C4;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_C5;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_C6;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_CLK;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_CO5;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_CO6;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_C_CY;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_C_XOR;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_D;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_D1;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_D2;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_D3;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_D4;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_D5;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_D6;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_DO5;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_DO6;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_D_CY;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_D_XOR;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X112Y131_SR;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_A;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_A1;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_A2;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_A3;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_A4;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_A5;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_A6;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_AO5;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_AO6;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_A_CY;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_A_XOR;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_B;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_B1;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_B2;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_B3;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_B4;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_B5;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_B6;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_BO5;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_BO6;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_B_CY;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_B_XOR;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_C;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_C1;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_C2;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_C3;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_C4;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_C5;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_C6;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_CO5;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_CO6;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_C_CY;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_C_XOR;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_D;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_D1;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_D2;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_D3;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_D4;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_D5;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_D6;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_DO5;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_DO6;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_D_CY;
  wire [0:0] CLBLM_L_X74Y131_SLICE_X113Y131_D_XOR;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_A;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_A1;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_A2;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_A3;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_A4;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_A5;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_A5Q;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_A6;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_AMUX;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_AO5;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_AO6;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_AQ;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_AX;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_A_CY;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_A_XOR;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_B;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_B1;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_B2;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_B3;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_B4;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_B5;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_B6;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_BMUX;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_BO5;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_BO6;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_B_CY;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_B_XOR;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_C;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_C1;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_C2;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_C3;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_C4;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_C5;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_C5Q;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_C6;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_CLK;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_CMUX;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_CO5;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_CO6;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_CQ;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_C_CY;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_C_XOR;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_D;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_D1;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_D2;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_D3;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_D4;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_D5;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_D6;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_DO5;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_DO6;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_D_CY;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_D_XOR;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X112Y132_SR;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_A;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_A1;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_A2;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_A3;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_A4;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_A5;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_A6;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_AO5;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_AO6;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_AQ;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_A_CY;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_A_XOR;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_B;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_B1;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_B2;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_B3;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_B4;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_B5;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_B6;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_BO5;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_BO6;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_BQ;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_B_CY;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_B_XOR;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_C;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_C1;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_C2;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_C3;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_C4;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_C5;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_C6;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_CLK;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_CO5;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_CO6;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_C_CY;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_C_XOR;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_D;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_D1;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_D2;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_D3;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_D4;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_D5;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_D6;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_DO5;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_DO6;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_D_CY;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_D_XOR;
  wire [0:0] CLBLM_L_X74Y132_SLICE_X113Y132_SR;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_A;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_A1;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_A2;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_A3;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_A4;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_A5;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_A6;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_AO5;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_AO6;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_AQ;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_A_CY;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_A_XOR;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_B;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_B1;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_B2;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_B3;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_B4;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_B5;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_B6;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_BO5;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_BO6;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_BQ;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_B_CY;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_B_XOR;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_C;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_C1;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_C2;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_C3;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_C4;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_C5;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_C6;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_CLK;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_CO5;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_CO6;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_CQ;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_C_CY;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_C_XOR;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_D;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_D1;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_D2;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_D3;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_D4;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_D5;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_D6;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_DMUX;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_DO5;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_DO6;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_D_CY;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_D_XOR;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X112Y133_SR;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_A;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_A1;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_A2;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_A3;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_A4;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_A5;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_A6;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_AMUX;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_AO5;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_AO6;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_A_CY;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_A_XOR;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_B;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_B1;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_B2;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_B3;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_B4;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_B5;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_B6;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_BO5;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_BO6;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_B_CY;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_B_XOR;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_C;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_C1;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_C2;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_C3;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_C4;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_C5;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_C6;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_CO5;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_CO6;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_C_CY;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_C_XOR;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_D;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_D1;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_D2;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_D3;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_D4;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_D5;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_D6;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_DO5;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_DO6;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_D_CY;
  wire [0:0] CLBLM_L_X74Y133_SLICE_X113Y133_D_XOR;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_A;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_A1;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_A2;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_A3;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_A4;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_A5;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_A6;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_AMUX;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_AO5;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_AO6;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_A_CY;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_A_XOR;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_B;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_B1;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_B2;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_B3;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_B4;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_B5;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_B6;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_BO5;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_BO6;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_BQ;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_B_CY;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_B_XOR;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_C;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_C1;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_C2;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_C3;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_C4;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_C5;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_C6;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_CLK;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_CO5;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_CO6;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_CQ;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_C_CY;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_C_XOR;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_D;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_D1;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_D2;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_D3;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_D4;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_D5;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_D6;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_DO5;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_DO6;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_DQ;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_D_CY;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_D_XOR;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X112Y134_SR;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_A;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_A1;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_A2;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_A3;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_A4;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_A5;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_A5Q;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_A6;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_AMUX;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_AO5;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_AO6;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_AQ;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_AX;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_A_CY;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_A_XOR;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_B;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_B1;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_B2;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_B3;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_B4;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_B5;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_B6;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_BO5;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_BO6;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_BQ;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_B_CY;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_B_XOR;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_C;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_C1;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_C2;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_C3;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_C4;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_C5;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_C6;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_CLK;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_CO5;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_CO6;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_CQ;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_C_CY;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_C_XOR;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_D;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_D1;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_D2;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_D3;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_D4;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_D5;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_D6;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_DMUX;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_DO5;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_DO6;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_D_CY;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_D_XOR;
  wire [0:0] CLBLM_L_X74Y134_SLICE_X113Y134_SR;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_A;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_A1;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_A2;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_A3;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_A4;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_A5;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_A6;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_AO5;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_AO6;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_AQ;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_A_CY;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_A_XOR;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_B;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_B1;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_B2;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_B3;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_B4;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_B5;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_B6;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_BO5;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_BO6;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_B_CY;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_B_XOR;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_C;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_C1;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_C2;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_C3;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_C4;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_C5;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_C6;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_CLK;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_CO5;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_CO6;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_C_CY;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_C_XOR;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_D;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_D1;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_D2;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_D3;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_D4;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_D5;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_D6;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_DO5;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_DO6;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_D_CY;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_D_XOR;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X112Y135_SR;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_A;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_A1;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_A2;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_A3;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_A4;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_A5;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_A6;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_AO5;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_AO6;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_AQ;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_A_CY;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_A_XOR;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_B;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_B1;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_B2;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_B3;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_B4;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_B5;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_B6;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_BO5;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_BO6;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_BQ;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_B_CY;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_B_XOR;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_C;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_C1;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_C2;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_C3;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_C4;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_C5;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_C6;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_CLK;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_CO5;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_CO6;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_C_CY;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_C_XOR;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_D;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_D1;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_D2;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_D3;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_D4;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_D5;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_D6;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_DO5;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_DO6;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_D_CY;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_D_XOR;
  wire [0:0] CLBLM_L_X74Y135_SLICE_X113Y135_SR;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_A;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_A1;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_A2;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_A3;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_A4;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_A5;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_A6;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_AO5;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_AO6;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_A_CY;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_A_XOR;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_B;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_B1;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_B2;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_B3;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_B4;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_B5;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_B6;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_BO5;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_BO6;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_B_CY;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_B_XOR;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_C;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_C1;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_C2;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_C3;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_C4;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_C5;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_C6;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_CO5;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_CO6;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_C_CY;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_C_XOR;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_D;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_D1;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_D2;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_D3;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_D4;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_D5;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_D6;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_DO5;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_DO6;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_D_CY;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X116Y109_D_XOR;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_A;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_A1;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_A2;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_A3;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_A4;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_A5;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_A6;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_AO5;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_AO6;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_A_CY;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_A_XOR;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_B;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_B1;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_B2;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_B3;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_B4;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_B5;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_B6;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_BO5;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_BO6;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_B_CY;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_B_XOR;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_C;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_C1;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_C2;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_C3;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_C4;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_C5;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_C6;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_CO5;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_CO6;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_C_CY;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_C_XOR;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_D;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_D1;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_D2;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_D3;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_D4;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_D5;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_D6;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_DO5;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_DO6;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_D_CY;
  wire [0:0] CLBLM_L_X76Y109_SLICE_X117Y109_D_XOR;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_A;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_A1;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_A2;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_A3;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_A4;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_A5;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_A6;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_AO5;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_AO6;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_AQ;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_AX;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_A_CY;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_A_XOR;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_B;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_B1;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_B2;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_B3;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_B4;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_B5;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_B6;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_BO5;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_BO6;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_BQ;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_BX;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_B_CY;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_B_XOR;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_C;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_C1;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_C2;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_C3;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_C4;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_C5;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_C6;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_CLK;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_CO5;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_CO6;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_C_CY;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_C_XOR;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_D;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_D1;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_D2;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_D3;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_D4;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_D5;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_D6;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_DO5;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_DO6;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_D_CY;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_D_XOR;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X116Y111_SR;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_A;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_A1;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_A2;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_A3;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_A4;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_A5;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_A6;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_AO5;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_AO6;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_A_CY;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_A_XOR;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_B;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_B1;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_B2;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_B3;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_B4;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_B5;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_B6;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_BO5;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_BO6;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_B_CY;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_B_XOR;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_C;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_C1;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_C2;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_C3;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_C4;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_C5;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_C6;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_CO5;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_CO6;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_C_CY;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_C_XOR;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_D;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_D1;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_D2;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_D3;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_D4;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_D5;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_D6;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_DO5;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_DO6;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_D_CY;
  wire [0:0] CLBLM_L_X76Y111_SLICE_X117Y111_D_XOR;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_A;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_A1;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_A2;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_A3;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_A4;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_A5;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_A5Q;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_A6;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_AMUX;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_AO5;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_AO6;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_AQ;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_AX;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_A_CY;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_A_XOR;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_B;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_B1;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_B2;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_B3;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_B4;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_B5;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_B6;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_BO5;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_BO6;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_BQ;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_BX;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_B_CY;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_B_XOR;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_C;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_C1;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_C2;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_C3;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_C4;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_C5;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_C6;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_CE;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_CLK;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_CO5;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_CO6;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_CQ;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_CX;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_C_CY;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_C_XOR;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_D;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_D1;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_D2;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_D3;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_D4;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_D5;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_D6;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_DO5;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_DO6;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_DQ;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_DX;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_D_CY;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_D_XOR;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X116Y118_SR;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_A;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_A1;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_A2;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_A3;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_A4;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_A5;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_A6;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_AO5;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_AO6;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_AQ;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_A_CY;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_A_XOR;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_B;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_B1;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_B2;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_B3;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_B4;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_B5;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_B6;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_BO5;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_BO6;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_BQ;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_B_CY;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_B_XOR;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_C;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_C1;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_C2;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_C3;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_C4;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_C5;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_C6;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_CLK;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_CO5;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_CO6;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_CQ;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_C_CY;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_C_XOR;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_D;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_D1;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_D2;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_D3;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_D4;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_D5;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_D6;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_DO5;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_DO6;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_D_CY;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_D_XOR;
  wire [0:0] CLBLM_L_X76Y118_SLICE_X117Y118_SR;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_A;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_A1;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_A2;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_A3;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_A4;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_A5;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_A5Q;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_A6;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_AMUX;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_AO5;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_AO6;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_AQ;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_A_CY;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_A_XOR;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_B;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_B1;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_B2;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_B3;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_B4;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_B5;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_B6;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_BO5;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_BO6;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_B_CY;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_B_XOR;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_C;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_C1;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_C2;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_C3;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_C4;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_C5;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_C6;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_CLK;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_CO5;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_CO6;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_C_CY;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_C_XOR;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_D;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_D1;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_D2;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_D3;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_D4;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_D5;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_D6;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_DO5;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_DO6;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_D_CY;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_D_XOR;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X116Y119_SR;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_A;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_A1;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_A2;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_A3;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_A4;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_A5;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_A6;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_AO5;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_AO6;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_A_CY;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_A_XOR;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_B;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_B1;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_B2;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_B3;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_B4;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_B5;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_B6;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_BO5;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_BO6;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_B_CY;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_B_XOR;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_C;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_C1;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_C2;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_C3;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_C4;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_C5;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_C6;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_CO5;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_CO6;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_C_CY;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_C_XOR;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_D;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_D1;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_D2;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_D3;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_D4;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_D5;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_D6;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_DO5;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_DO6;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_D_CY;
  wire [0:0] CLBLM_L_X76Y119_SLICE_X117Y119_D_XOR;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_A;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_A1;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_A2;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_A3;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_A4;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_A5;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_A5Q;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_A6;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_AMUX;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_AO5;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_AO6;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_AQ;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_A_CY;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_A_XOR;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_B;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_B1;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_B2;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_B3;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_B4;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_B5;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_B6;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_BO5;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_BO6;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_BQ;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_B_CY;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_B_XOR;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_C;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_C1;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_C2;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_C3;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_C4;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_C5;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_C5Q;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_C6;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_CLK;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_CMUX;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_CO5;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_CO6;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_CQ;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_C_CY;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_C_XOR;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_D;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_D1;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_D2;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_D3;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_D4;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_D5;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_D6;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_DO5;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_DO6;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_D_CY;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_D_XOR;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X116Y122_SR;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_A;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_A1;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_A2;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_A3;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_A4;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_A5;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_A6;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_AO5;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_AO6;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_AQ;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_AX;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_A_CY;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_A_XOR;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_B;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_B1;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_B2;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_B3;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_B4;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_B5;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_B6;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_BO5;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_BO6;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_B_CY;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_B_XOR;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_C;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_C1;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_C2;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_C3;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_C4;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_C5;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_C6;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_CLK;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_CO5;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_CO6;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_C_CY;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_C_XOR;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_D;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_D1;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_D2;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_D3;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_D4;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_D5;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_D6;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_DO5;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_DO6;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_D_CY;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_D_XOR;
  wire [0:0] CLBLM_L_X76Y122_SLICE_X117Y122_SR;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_A;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_A1;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_A2;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_A3;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_A4;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_A5;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_A5Q;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_A6;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_AMUX;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_AO5;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_AO6;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_AQ;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_AX;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_A_CY;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_A_XOR;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_B;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_B1;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_B2;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_B3;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_B4;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_B5;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_B6;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_BO5;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_BO6;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_BQ;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_B_CY;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_B_XOR;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_C;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_C1;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_C2;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_C3;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_C4;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_C5;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_C6;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_CLK;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_CO5;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_CO6;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_CQ;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_C_CY;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_C_XOR;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_D;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_D1;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_D2;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_D3;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_D4;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_D5;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_D6;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_DO5;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_DO6;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_D_CY;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_D_XOR;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X116Y123_SR;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_A;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_A1;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_A2;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_A3;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_A4;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_A5;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_A6;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_AMUX;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_AO5;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_AO6;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_AQ;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_A_CY;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_A_XOR;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_B;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_B1;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_B2;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_B3;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_B4;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_B5;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_B5Q;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_B6;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_BMUX;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_BO5;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_BO6;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_BQ;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_B_CY;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_B_XOR;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_C;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_C1;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_C2;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_C3;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_C4;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_C5;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_C6;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_CLK;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_CO5;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_CO6;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_CQ;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_C_CY;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_C_XOR;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_D;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_D1;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_D2;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_D3;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_D4;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_D5;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_D6;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_DO5;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_DO6;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_D_CY;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_D_XOR;
  wire [0:0] CLBLM_L_X76Y123_SLICE_X117Y123_SR;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_A;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_A1;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_A2;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_A3;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_A4;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_A5;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_A5Q;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_A6;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_AMUX;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_AO5;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_AO6;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_AQ;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_AX;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_A_CY;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_A_XOR;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_B;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_B1;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_B2;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_B3;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_B4;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_B5;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_B5Q;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_B6;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_BMUX;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_BO5;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_BO6;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_BQ;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_BX;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_B_CY;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_B_XOR;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_C;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_C1;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_C2;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_C3;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_C4;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_C5;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_C6;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_CE;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_CLK;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_CO5;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_CO6;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_CQ;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_CX;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_C_CY;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_C_XOR;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_D;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_D1;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_D2;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_D3;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_D4;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_D5;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_D6;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_DO5;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_DO6;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_DQ;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_DX;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_D_CY;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_D_XOR;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_SR;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_A;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_A1;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_A2;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_A3;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_A4;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_A5;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_A6;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_AO5;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_AO6;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_AQ;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_A_CY;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_A_XOR;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_B;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_B1;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_B2;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_B3;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_B4;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_B5;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_B6;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_BO5;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_BO6;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_BQ;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_B_CY;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_B_XOR;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_C;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_C1;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_C2;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_C3;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_C4;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_C5;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_C6;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_CLK;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_CO5;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_CO6;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_C_CY;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_C_XOR;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_D;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_D1;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_D2;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_D3;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_D4;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_D5;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_D6;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_DO5;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_DO6;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_D_CY;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_D_XOR;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_SR;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_A;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_A1;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_A2;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_A3;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_A4;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_A5;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_A5Q;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_A6;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_AMUX;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_AO5;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_AO6;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_AQ;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_A_CY;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_A_XOR;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_B;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_B1;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_B2;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_B3;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_B4;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_B5;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_B6;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_BO5;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_BO6;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_BQ;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_B_CY;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_B_XOR;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_C;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_C1;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_C2;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_C3;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_C4;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_C5;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_C5Q;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_C6;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_CLK;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_CMUX;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_CO5;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_CO6;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_CQ;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_C_CY;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_C_XOR;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_D;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_D1;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_D2;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_D3;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_D4;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_D5;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_D6;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_DO5;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_DO6;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_D_CY;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_D_XOR;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_SR;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_A;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_A1;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_A2;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_A3;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_A4;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_A5;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_A6;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_AO5;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_AO6;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_AQ;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_A_CY;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_A_XOR;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_B;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_B1;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_B2;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_B3;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_B4;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_B5;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_B6;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_BO5;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_BO6;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_BQ;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_B_CY;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_B_XOR;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_C;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_C1;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_C2;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_C3;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_C4;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_C5;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_C6;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_CLK;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_CO5;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_CO6;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_C_CY;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_C_XOR;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_D;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_D1;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_D2;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_D3;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_D4;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_D5;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_D6;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_DO5;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_DO6;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_D_CY;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_D_XOR;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_SR;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_A;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_A1;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_A2;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_A3;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_A4;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_A5;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_A6;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_AMUX;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_AO5;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_AO6;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_A_CY;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_A_XOR;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_B;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_B1;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_B2;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_B3;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_B4;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_B5;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_B5Q;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_B6;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_BMUX;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_BO5;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_BO6;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_BQ;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_B_CY;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_B_XOR;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_C;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_C1;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_C2;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_C3;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_C4;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_C5;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_C6;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_CLK;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_CO5;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_CO6;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_CQ;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_C_CY;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_C_XOR;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_D;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_D1;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_D2;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_D3;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_D4;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_D5;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_D6;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_DO5;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_DO6;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_DQ;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_D_CY;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_D_XOR;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X116Y126_SR;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_A;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_A1;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_A2;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_A3;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_A4;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_A5;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_A6;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_AO5;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_AO6;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_AQ;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_A_CY;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_A_XOR;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_B;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_B1;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_B2;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_B3;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_B4;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_B5;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_B6;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_BO5;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_BO6;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_B_CY;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_B_XOR;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_C;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_C1;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_C2;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_C3;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_C4;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_C5;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_C6;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_CLK;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_CO5;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_CO6;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_C_CY;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_C_XOR;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_D;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_D1;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_D2;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_D3;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_D4;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_D5;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_D6;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_DO5;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_DO6;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_D_CY;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_D_XOR;
  wire [0:0] CLBLM_L_X76Y126_SLICE_X117Y126_SR;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_A;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_A1;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_A2;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_A3;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_A4;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_A5;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_A6;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_AO5;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_AO6;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_AQ;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_AX;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_A_CY;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_A_XOR;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_B;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_B1;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_B2;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_B3;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_B4;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_B5;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_B6;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_BO5;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_BO6;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_B_CY;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_B_XOR;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_C;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_C1;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_C2;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_C3;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_C4;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_C5;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_C6;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_CLK;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_CO5;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_C_CY;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_C_XOR;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_D;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_D1;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_D2;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_D3;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_D4;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_D5;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_D6;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_DO5;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_DO6;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_D_CY;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_D_XOR;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_SR;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_A;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_A1;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_A2;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_A3;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_A4;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_A5;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_A6;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_AO5;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_AO6;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_A_CY;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_A_XOR;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_B;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_B1;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_B2;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_B3;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_B4;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_B5;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_B6;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_BO5;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_BO6;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_B_CY;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_B_XOR;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_C;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_C1;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_C2;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_C3;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_C4;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_C5;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_C6;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_CO5;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_CO6;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_C_CY;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_C_XOR;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_D;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_D1;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_D2;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_D3;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_D4;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_D5;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_D6;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_DO5;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_DO6;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_D_CY;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_D_XOR;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_A;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_A1;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_A2;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_A3;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_A4;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_A5;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_A5Q;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_A6;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_AMUX;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_AO5;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_AO6;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_AQ;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_AX;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_A_CY;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_A_XOR;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_B;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_B1;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_B2;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_B3;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_B4;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_B5;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_B6;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_BO5;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_BO6;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_BQ;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_B_CY;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_B_XOR;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_C;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_C1;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_C2;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_C3;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_C4;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_C5;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_C5Q;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_C6;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_CLK;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_CMUX;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_CO5;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_CO6;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_CQ;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_C_CY;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_C_XOR;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_D;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_D1;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_D2;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_D3;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_D4;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_D5;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_D6;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_DO5;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_DO6;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_D_CY;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_D_XOR;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_SR;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_A;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_A1;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_A2;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_A3;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_A4;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_A5;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_A5Q;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_A6;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_AMUX;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_AO5;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_AO6;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_AQ;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_AX;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_A_CY;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_A_XOR;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_B;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_B1;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_B2;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_B3;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_B4;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_B5;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_B5Q;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_B6;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_BMUX;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_BO5;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_BO6;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_BQ;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_B_CY;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_B_XOR;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_C;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_C1;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_C2;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_C3;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_C4;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_C5;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_C6;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_CLK;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_CMUX;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_CO5;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_CO6;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_C_CY;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_C_XOR;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_D;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_D1;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_D2;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_D3;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_D4;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_D5;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_D6;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_DO5;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_DO6;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_D_CY;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_D_XOR;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_SR;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_A;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_A1;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_A2;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_A3;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_A4;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_A5;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_A6;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_AMUX;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_AO5;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_AO6;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_AQ;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_AX;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_A_CY;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_A_XOR;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_B;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_B1;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_B2;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_B3;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_B4;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_B5;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_B5Q;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_B6;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_BMUX;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_BO5;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_BO6;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_BQ;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_BX;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_B_CY;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_B_XOR;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_C;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_C1;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_C2;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_C3;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_C4;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_C5;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_C6;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_CLK;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_CO5;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_CO6;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_CQ;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_C_CY;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_C_XOR;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_D;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_D1;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_D2;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_D3;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_D4;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_D5;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_D6;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_DMUX;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_DO5;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_DO6;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_D_CY;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_D_XOR;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X116Y129_SR;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_A;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_A1;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_A2;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_A3;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_A4;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_A5;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_A6;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_AO5;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_AO6;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_A_CY;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_A_XOR;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_B;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_B1;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_B2;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_B3;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_B4;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_B5;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_B6;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_BO5;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_BO6;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_B_CY;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_B_XOR;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_C;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_C1;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_C2;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_C3;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_C4;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_C5;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_C6;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_CO5;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_CO6;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_C_CY;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_C_XOR;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_D;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_D1;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_D2;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_D3;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_D4;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_D5;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_D6;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_DO5;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_DO6;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_D_CY;
  wire [0:0] CLBLM_L_X76Y129_SLICE_X117Y129_D_XOR;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_A;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_A1;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_A2;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_A3;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_A4;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_A5;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_A5Q;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_A6;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_AMUX;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_AO5;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_AO6;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_AQ;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_AX;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_A_CY;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_A_XOR;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_B;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_B1;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_B2;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_B3;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_B4;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_B5;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_B6;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_BO5;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_BO6;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_BQ;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_B_CY;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_B_XOR;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_C;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_C1;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_C2;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_C3;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_C4;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_C5;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_C6;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_CLK;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_CMUX;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_CO5;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_CO6;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_C_CY;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_C_XOR;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_D;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_D1;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_D2;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_D3;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_D4;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_D5;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_D6;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_DO5;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_DO6;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_DQ;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_D_CY;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_D_XOR;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X116Y130_SR;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_A;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_A1;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_A2;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_A3;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_A4;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_A5;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_A6;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_AO5;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_AO6;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_A_CY;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_A_XOR;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_B;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_B1;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_B2;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_B3;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_B4;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_B5;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_B6;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_BO5;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_BO6;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_B_CY;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_B_XOR;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_C;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_C1;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_C2;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_C3;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_C4;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_C5;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_C6;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_CO5;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_CO6;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_C_CY;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_C_XOR;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_D;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_D1;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_D2;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_D3;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_D4;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_D5;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_D6;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_DO5;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_DO6;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_D_CY;
  wire [0:0] CLBLM_L_X76Y130_SLICE_X117Y130_D_XOR;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_A;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_A1;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_A2;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_A3;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_A4;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_A5;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_A6;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_AO5;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_AO6;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_AQ;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_A_CY;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_A_XOR;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_B;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_B1;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_B2;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_B3;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_B4;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_B5;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_B6;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_BO5;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_BO6;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_BQ;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_B_CY;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_B_XOR;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_C;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_C1;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_C2;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_C3;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_C4;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_C5;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_C6;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_CLK;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_CO5;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_CO6;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_C_CY;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_C_XOR;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_D;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_D1;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_D2;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_D3;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_D4;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_D5;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_D6;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_DO5;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_DO6;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_D_CY;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_D_XOR;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_SR;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_A;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_A1;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_A2;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_A3;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_A4;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_A5;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_A6;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_AO5;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_AO6;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_A_CY;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_A_XOR;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_B;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_B1;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_B2;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_B3;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_B4;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_B5;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_B6;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_BO5;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_BO6;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_B_CY;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_B_XOR;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_C;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_C1;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_C2;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_C3;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_C4;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_C5;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_C6;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_CO5;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_CO6;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_C_CY;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_C_XOR;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_D;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_D1;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_D2;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_D3;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_D4;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_D5;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_D6;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_DO5;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_DO6;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_D_CY;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_D_XOR;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_A;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_A1;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_A2;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_A3;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_A4;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_A5;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_A6;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_AO5;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_AO6;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_AQ;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_A_CY;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_A_XOR;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_B;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_B1;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_B2;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_B3;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_B4;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_B5;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_B6;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_BO5;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_BO6;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_BQ;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_B_CY;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_B_XOR;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_C;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_C1;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_C2;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_C3;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_C4;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_C5;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_C6;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_CLK;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_CO5;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_CO6;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_C_CY;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_C_XOR;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_D;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_D1;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_D2;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_D3;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_D4;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_D5;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_D6;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_DO5;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_DO6;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_D_CY;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_D_XOR;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X116Y134_SR;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_A;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_A1;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_A2;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_A3;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_A4;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_A5;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_A6;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_AO5;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_AO6;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_AQ;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_A_CY;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_A_XOR;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_B;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_B1;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_B2;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_B3;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_B4;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_B5;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_B6;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_BO5;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_BO6;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_BQ;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_B_CY;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_B_XOR;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_C;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_C1;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_C2;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_C3;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_C4;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_C5;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_C6;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_CLK;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_CMUX;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_CO5;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_CO6;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_C_CY;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_C_XOR;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_D;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_D1;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_D2;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_D3;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_D4;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_D5;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_D6;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_DO5;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_DO6;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_D_CY;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_D_XOR;
  wire [0:0] CLBLM_L_X76Y134_SLICE_X117Y134_SR;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_A;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_A1;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_A2;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_A3;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_A4;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_A5;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_A5Q;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_A6;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_AMUX;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_AO5;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_AO6;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_AQ;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_A_CY;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_A_XOR;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_B;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_B1;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_B2;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_B3;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_B4;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_B5;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_B6;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_BO5;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_BO6;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_BQ;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_BX;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_B_CY;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_B_XOR;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_C;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_C1;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_C2;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_C3;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_C4;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_C5;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_C6;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_CLK;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_CO5;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_CO6;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_C_CY;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_C_XOR;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_D;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_D1;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_D2;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_D3;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_D4;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_D5;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_D6;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_DO5;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_DO6;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_D_CY;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_D_XOR;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X120Y104_SR;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_A;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_A1;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_A2;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_A3;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_A4;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_A5;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_A6;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_AO5;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_AO6;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_A_CY;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_A_XOR;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_B;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_B1;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_B2;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_B3;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_B4;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_B5;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_B6;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_BO5;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_BO6;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_B_CY;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_B_XOR;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_C;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_C1;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_C2;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_C3;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_C4;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_C5;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_C6;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_CO5;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_CO6;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_C_CY;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_C_XOR;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_D;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_D1;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_D2;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_D3;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_D4;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_D5;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_D6;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_DO5;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_DO6;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_D_CY;
  wire [0:0] CLBLM_L_X78Y104_SLICE_X121Y104_D_XOR;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_A;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_A1;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_A2;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_A3;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_A4;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_A5;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_A6;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_AO5;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_AO6;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_AQ;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_AX;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_A_CY;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_A_XOR;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_B;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_B1;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_B2;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_B3;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_B4;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_B5;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_B6;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_BO5;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_BO6;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_B_CY;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_B_XOR;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_C;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_C1;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_C2;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_C3;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_C4;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_C5;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_C6;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_CLK;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_CO5;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_CO6;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_C_CY;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_C_XOR;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_D;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_D1;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_D2;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_D3;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_D4;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_D5;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_D6;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_DO5;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_DO6;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_D_CY;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_D_XOR;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X120Y106_SR;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_A;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_A1;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_A2;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_A3;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_A4;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_A5;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_A6;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_AO5;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_AO6;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_A_CY;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_A_XOR;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_B;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_B1;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_B2;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_B3;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_B4;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_B5;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_B6;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_BO5;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_BO6;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_B_CY;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_B_XOR;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_C;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_C1;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_C2;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_C3;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_C4;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_C5;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_C6;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_CO5;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_CO6;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_C_CY;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_C_XOR;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_D;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_D1;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_D2;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_D3;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_D4;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_D5;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_D6;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_DO5;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_DO6;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_D_CY;
  wire [0:0] CLBLM_L_X78Y106_SLICE_X121Y106_D_XOR;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_A;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_A1;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_A2;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_A3;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_A4;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_A5;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_A6;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_AO5;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_AO6;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_AQ;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_A_CY;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_A_XOR;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_B;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_B1;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_B2;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_B3;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_B4;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_B5;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_B6;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_BO5;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_BO6;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_B_CY;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_B_XOR;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_C;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_C1;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_C2;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_C3;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_C4;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_C5;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_C6;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_CLK;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_CO5;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_CO6;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_C_CY;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_C_XOR;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_D;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_D1;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_D2;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_D3;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_D4;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_D5;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_D6;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_DO5;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_DO6;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_D_CY;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_D_XOR;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_SR;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_A;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_A1;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_A2;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_A3;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_A4;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_A5;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_A6;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_AO5;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_AO6;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_A_CY;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_A_XOR;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_B;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_B1;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_B2;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_B3;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_B4;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_B5;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_B6;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_BO5;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_BO6;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_B_CY;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_B_XOR;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_C;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_C1;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_C2;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_C3;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_C4;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_C5;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_C6;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_CO5;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_CO6;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_C_CY;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_C_XOR;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_D;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_D1;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_D2;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_D3;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_D4;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_D5;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_D6;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_DO5;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_DO6;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_D_CY;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_D_XOR;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_A;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_A1;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_A2;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_A3;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_A4;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_A5;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_A6;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_AO5;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_AO6;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_AQ;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_A_CY;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_A_XOR;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_B;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_B1;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_B2;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_B3;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_B4;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_B5;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_B6;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_BO5;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_BO6;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_BQ;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_B_CY;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_B_XOR;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_C;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_C1;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_C2;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_C3;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_C4;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_C5;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_C6;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_CLK;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_CMUX;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_CO5;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_CO6;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_C_CY;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_C_XOR;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_D;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_D1;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_D2;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_D3;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_D4;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_D5;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_D6;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_DO5;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_DO6;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_D_CY;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_D_XOR;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_SR;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_A;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_A1;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_A2;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_A3;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_A4;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_A5;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_A6;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_AO5;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_AO6;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_A_CY;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_A_XOR;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_B;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_B1;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_B2;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_B3;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_B4;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_B5;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_B6;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_BO5;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_BO6;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_B_CY;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_B_XOR;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_C;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_C1;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_C2;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_C3;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_C4;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_C5;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_C6;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_CO5;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_CO6;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_C_CY;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_C_XOR;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_D;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_D1;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_D2;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_D3;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_D4;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_D5;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_D6;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_DO5;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_DO6;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_D_CY;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_D_XOR;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_A;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_A1;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_A2;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_A3;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_A4;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_A5;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_A6;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_AMUX;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_AO5;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_AO6;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_A_CY;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_A_XOR;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_B;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_B1;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_B2;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_B3;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_B4;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_B5;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_B6;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_BO5;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_BO6;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_B_CY;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_B_XOR;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_C;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_C1;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_C2;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_C3;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_C4;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_C5;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_C6;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_CO5;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_CO6;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_C_CY;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_C_XOR;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_D;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_D1;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_D2;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_D3;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_D4;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_D5;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_D6;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_DO5;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_DO6;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_D_CY;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_D_XOR;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_A;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_A1;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_A2;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_A3;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_A4;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_A5;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_A6;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_AO5;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_AO6;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_AQ;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_A_CY;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_A_XOR;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_B;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_B1;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_B2;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_B3;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_B4;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_B5;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_B6;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_BO5;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_BO6;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_BQ;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_B_CY;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_B_XOR;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_C;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_C1;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_C2;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_C3;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_C4;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_C5;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_C6;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_CLK;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_CO5;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_CO6;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_C_CY;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_C_XOR;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_D;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_D1;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_D2;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_D3;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_D4;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_D5;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_D6;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_DO5;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_DO6;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_D_CY;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_D_XOR;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_SR;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_A;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_A1;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_A2;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_A3;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_A4;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_A5;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_A6;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_AMUX;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_AO5;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_AO6;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_A_CY;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_A_XOR;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_B;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_B1;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_B2;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_B3;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_B4;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_B5;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_B6;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_BO5;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_BO6;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_B_CY;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_B_XOR;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_C;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_C1;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_C2;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_C3;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_C4;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_C5;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_C6;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_CO5;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_CO6;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_C_CY;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_C_XOR;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_D;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_D1;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_D2;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_D3;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_D4;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_D5;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_D6;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_DO5;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_DO6;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_D_CY;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_D_XOR;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_A;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_A1;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_A2;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_A3;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_A4;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_A5;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_A5Q;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_A6;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_AMUX;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_AO5;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_AO6;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_AQ;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_A_CY;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_A_XOR;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_B;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_B1;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_B2;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_B3;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_B4;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_B5;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_B6;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_BO5;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_BO6;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_BQ;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_B_CY;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_B_XOR;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_C;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_C1;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_C2;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_C3;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_C4;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_C5;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_C6;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_CLK;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_CMUX;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_CO5;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_CO6;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_C_CY;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_C_XOR;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_D;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_D1;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_D2;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_D3;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_D4;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_D5;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_D6;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_DO5;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_DO6;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_D_CY;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_D_XOR;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_SR;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_A;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_A1;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_A2;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_A3;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_A4;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_A5;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_A6;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_AO5;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_AO6;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_AQ;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_A_CY;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_A_XOR;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_B;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_B1;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_B2;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_B3;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_B4;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_B5;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_B6;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_BO5;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_BO6;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_BQ;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_B_CY;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_B_XOR;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_C;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_C1;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_C2;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_C3;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_C4;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_C5;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_C6;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_CLK;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_CO5;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_CO6;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_CQ;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_C_CY;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_C_XOR;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_D;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_D1;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_D2;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_D3;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_D4;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_D5;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_D6;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_DO5;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_DO6;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_D_CY;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_D_XOR;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_SR;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_A;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_A1;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_A2;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_A3;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_A4;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_A5;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_A6;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_AO5;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_AO6;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_A_CY;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_A_XOR;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_B;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_B1;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_B2;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_B3;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_B4;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_B5;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_B6;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_BO5;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_BO6;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_B_CY;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_B_XOR;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_C;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_C1;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_C2;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_C3;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_C4;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_C5;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_C6;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_CO5;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_CO6;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_C_CY;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_C_XOR;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_D;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_D1;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_D2;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_D3;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_D4;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_D5;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_D6;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_DO5;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_DO6;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_D_CY;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_D_XOR;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_A;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_A1;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_A2;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_A3;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_A4;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_A5;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_A6;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_AO5;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_AO6;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_A_CY;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_A_XOR;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_B;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_B1;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_B2;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_B3;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_B4;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_B5;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_B6;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_BO5;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_BO6;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_B_CY;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_B_XOR;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_C;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_C1;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_C2;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_C3;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_C4;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_C5;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_C6;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_CO5;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_CO6;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_C_CY;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_C_XOR;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_D;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_D1;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_D2;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_D3;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_D4;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_D5;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_D6;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_DO5;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_DO6;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_D_CY;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X120Y127_D_XOR;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_A;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_A1;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_A2;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_A3;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_A4;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_A5;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_A6;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_AMUX;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_AO5;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_AO6;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_A_CY;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_A_XOR;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_B;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_B1;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_B2;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_B3;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_B4;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_B5;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_B6;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_BO5;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_BO6;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_B_CY;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_B_XOR;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_C;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_C1;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_C2;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_C3;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_C4;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_C5;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_C6;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_CO5;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_CO6;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_C_CY;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_C_XOR;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_D;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_D1;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_D2;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_D3;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_D4;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_D5;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_D6;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_DO5;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_DO6;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_D_CY;
  wire [0:0] CLBLM_L_X78Y127_SLICE_X121Y127_D_XOR;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_A;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_A1;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_A2;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_A3;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_A4;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_A5;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_A6;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_AO5;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_AO6;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_AQ;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_A_CY;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_A_XOR;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_B;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_B1;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_B2;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_B3;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_B4;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_B5;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_B6;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_BO5;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_BO6;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_B_CY;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_B_XOR;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_C;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_C1;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_C2;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_C3;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_C4;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_C5;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_C6;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_CLK;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_CO5;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_CO6;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_C_CY;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_C_XOR;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_D;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_D1;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_D2;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_D3;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_D4;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_D5;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_D6;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_DO5;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_DO6;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_D_CY;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_D_XOR;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X120Y128_SR;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_A;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_A1;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_A2;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_A3;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_A4;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_A5;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_A6;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_AO5;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_AO6;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_A_CY;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_A_XOR;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_B;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_B1;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_B2;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_B3;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_B4;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_B5;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_B6;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_BO5;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_BO6;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_B_CY;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_B_XOR;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_C;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_C1;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_C2;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_C3;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_C4;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_C5;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_C6;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_CO5;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_CO6;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_C_CY;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_C_XOR;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_D;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_D1;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_D2;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_D3;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_D4;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_D5;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_D6;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_DO5;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_DO6;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_D_CY;
  wire [0:0] CLBLM_L_X78Y128_SLICE_X121Y128_D_XOR;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_A;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_A1;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_A2;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_A3;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_A4;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_A5;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_A6;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_AO5;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_AO6;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_A_CY;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_A_XOR;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_B;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_B1;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_B2;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_B3;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_B4;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_B5;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_B6;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_BO5;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_BO6;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_B_CY;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_B_XOR;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_C;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_C1;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_C2;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_C3;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_C4;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_C5;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_C6;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_CO5;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_CO6;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_C_CY;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_C_XOR;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_D;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_D1;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_D2;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_D3;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_D4;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_D5;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_D6;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_DO5;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_DO6;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_D_CY;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_D_XOR;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_A;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_A1;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_A2;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_A3;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_A4;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_A5;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_A6;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_AO5;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_AO6;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_A_CY;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_A_XOR;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_B;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_B1;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_B2;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_B3;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_B4;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_B5;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_B6;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_BO5;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_BO6;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_B_CY;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_B_XOR;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_C;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_C1;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_C2;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_C3;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_C4;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_C5;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_C6;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_CO5;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_CO6;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_C_CY;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_C_XOR;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_D;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_D1;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_D2;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_D3;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_D4;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_D5;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_D6;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_DO5;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_DO6;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_D_CY;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_D_XOR;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_A;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_A1;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_A2;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_A3;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_A4;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_A5;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_A6;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_AO5;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_AO6;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_AQ;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_A_CY;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_A_XOR;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_B;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_B1;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_B2;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_B3;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_B4;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_B5;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_B6;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_BO5;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_BO6;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_BQ;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_B_CY;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_B_XOR;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_C;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_C1;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_C2;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_C3;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_C4;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_C5;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_C6;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_CLK;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_CO5;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_CO6;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_C_CY;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_C_XOR;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_D;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_D1;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_D2;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_D3;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_D4;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_D5;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_D6;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_DO5;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_DO6;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_D_CY;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_D_XOR;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X120Y130_SR;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_A;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_A1;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_A2;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_A3;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_A4;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_A5;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_A6;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_AO5;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_AO6;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_A_CY;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_A_XOR;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_B;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_B1;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_B2;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_B3;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_B4;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_B5;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_B6;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_BO5;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_BO6;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_B_CY;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_B_XOR;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_C;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_C1;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_C2;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_C3;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_C4;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_C5;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_C6;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_CO5;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_CO6;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_C_CY;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_C_XOR;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_D;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_D1;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_D2;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_D3;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_D4;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_D5;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_D6;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_DO5;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_DO6;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_D_CY;
  wire [0:0] CLBLM_L_X78Y130_SLICE_X121Y130_D_XOR;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_A;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_A1;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_A2;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_A3;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_A4;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_A5;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_A6;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_AO5;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_AO6;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_AQ;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_A_CY;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_A_XOR;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_B;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_B1;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_B2;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_B3;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_B4;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_B5;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_B6;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_BO5;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_BO6;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_B_CY;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_B_XOR;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_C;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_C1;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_C2;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_C3;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_C4;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_C5;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_C6;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_CLK;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_CO5;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_CO6;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_C_CY;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_C_XOR;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_D;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_D1;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_D2;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_D3;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_D4;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_D5;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_D6;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_DO5;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_DO6;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_D_CY;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_D_XOR;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X120Y131_SR;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_A;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_A1;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_A2;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_A3;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_A4;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_A5;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_A6;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_AO5;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_AO6;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_A_CY;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_A_XOR;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_B;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_B1;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_B2;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_B3;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_B4;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_B5;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_B6;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_BO5;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_BO6;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_B_CY;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_B_XOR;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_C;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_C1;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_C2;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_C3;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_C4;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_C5;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_C6;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_CO5;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_CO6;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_C_CY;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_C_XOR;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_D;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_D1;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_D2;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_D3;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_D4;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_D5;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_D6;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_DO5;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_DO6;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_D_CY;
  wire [0:0] CLBLM_L_X78Y131_SLICE_X121Y131_D_XOR;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_A;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_A1;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_A2;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_A3;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_A4;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_A5;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_A6;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_AO5;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_AO6;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_AQ;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_AX;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_A_CY;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_A_XOR;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_B;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_B1;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_B2;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_B3;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_B4;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_B5;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_B6;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_BO5;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_BO6;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_B_CY;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_B_XOR;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_C;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_C1;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_C2;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_C3;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_C4;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_C5;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_C6;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_CLK;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_CO5;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_CO6;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_C_CY;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_C_XOR;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_D;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_D1;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_D2;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_D3;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_D4;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_D5;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_D6;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_DO5;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_DO6;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_D_CY;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_D_XOR;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X124Y132_SR;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_A;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_A1;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_A2;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_A3;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_A4;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_A5;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_A6;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_AO5;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_AO6;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_A_CY;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_A_XOR;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_B;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_B1;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_B2;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_B3;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_B4;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_B5;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_B6;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_BO5;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_BO6;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_B_CY;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_B_XOR;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_C;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_C1;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_C2;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_C3;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_C4;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_C5;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_C6;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_CO5;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_CO6;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_C_CY;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_C_XOR;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_D;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_D1;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_D2;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_D3;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_D4;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_D5;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_D6;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_DO5;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_DO6;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_D_CY;
  wire [0:0] CLBLM_L_X80Y132_SLICE_X125Y132_D_XOR;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_A;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_A1;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_A2;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_A3;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_A4;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_A5;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_A6;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_AO5;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_AO6;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_AQ;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_AX;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_A_CY;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_A_XOR;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_B;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_B1;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_B2;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_B3;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_B4;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_B5;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_B6;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_BO5;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_BO6;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_B_CY;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_B_XOR;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_C;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_C1;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_C2;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_C3;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_C4;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_C5;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_C6;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_CLK;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_CO5;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_CO6;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_C_CY;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_C_XOR;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_D;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_D1;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_D2;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_D3;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_D4;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_D5;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_D6;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_DO5;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_DO6;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_D_CY;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_D_XOR;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X128Y130_SR;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_A;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_A1;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_A2;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_A3;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_A4;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_A5;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_A6;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_AO5;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_AO6;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_A_CY;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_A_XOR;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_B;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_B1;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_B2;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_B3;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_B4;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_B5;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_B6;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_BO5;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_BO6;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_B_CY;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_B_XOR;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_C;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_C1;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_C2;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_C3;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_C4;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_C5;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_C6;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_CO5;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_CO6;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_C_CY;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_C_XOR;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_D;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_D1;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_D2;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_D3;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_D4;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_D5;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_D6;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_DO5;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_DO6;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_D_CY;
  wire [0:0] CLBLM_L_X82Y130_SLICE_X129Y130_D_XOR;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_A;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_A1;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_A2;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_A3;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_A4;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_A5;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_A5Q;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_A6;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_AMUX;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_AO5;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_AO6;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_AQ;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_A_CY;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_A_XOR;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_B;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_B1;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_B2;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_B3;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_B4;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_B5;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_B6;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_BO5;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_BO6;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_BQ;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_BX;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_B_CY;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_B_XOR;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_C;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_C1;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_C2;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_C3;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_C4;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_C5;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_C6;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_CLK;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_CO5;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_CO6;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_C_CY;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_C_XOR;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_D;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_D1;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_D2;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_D3;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_D4;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_D5;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_D6;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_DO5;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_DO6;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_D_CY;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_D_XOR;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X128Y98_SR;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_A;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_A1;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_A2;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_A3;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_A4;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_A5;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_A6;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_AO5;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_AO6;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_A_CY;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_A_XOR;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_B;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_B1;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_B2;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_B3;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_B4;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_B5;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_B6;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_BO5;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_BO6;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_B_CY;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_B_XOR;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_C;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_C1;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_C2;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_C3;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_C4;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_C5;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_C6;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_CO5;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_CO6;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_C_CY;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_C_XOR;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_D;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_D1;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_D2;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_D3;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_D4;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_D5;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_D6;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_DO5;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_DO6;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_D_CY;
  wire [0:0] CLBLM_L_X82Y98_SLICE_X129Y98_D_XOR;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_A;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_A1;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_A2;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_A3;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_A4;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_A5;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_A6;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_AO5;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_AO6;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_AQ;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_AX;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_A_CY;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_A_XOR;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_B;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_B1;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_B2;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_B3;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_B4;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_B5;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_B6;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_BO5;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_BO6;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_BQ;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_BX;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_B_CY;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_B_XOR;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_C;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_C1;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_C2;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_C3;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_C4;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_C5;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_C6;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_CLK;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_CO5;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_CO6;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_CQ;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_CX;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_C_CY;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_C_XOR;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_D;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_D1;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_D2;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_D3;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_D4;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_D5;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_D6;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_DO5;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_DO6;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_D_CY;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_D_XOR;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X162Y67_SR;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_A;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_A1;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_A2;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_A3;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_A4;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_A5;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_A6;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_AO5;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_AO6;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_AQ;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_AX;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_A_CY;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_A_XOR;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_B;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_B1;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_B2;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_B3;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_B4;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_B5;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_B6;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_BO5;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_BO6;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_BQ;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_BX;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_B_CY;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_B_XOR;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_C;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_C1;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_C2;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_C3;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_C4;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_C5;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_C6;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_CLK;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_CO5;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_CO6;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_CQ;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_CX;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_C_CY;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_C_XOR;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_D;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_D1;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_D2;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_D3;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_D4;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_D5;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_D6;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_DO5;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_DO6;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_D_CY;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_D_XOR;
  wire [0:0] CLBLM_R_X103Y67_SLICE_X163Y67_SR;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_A;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_A1;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_A2;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_A3;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_A4;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_A5;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_A5Q;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_A6;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_AMUX;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_AO5;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_AO6;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_AQ;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_AX;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_A_CY;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_A_XOR;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_B;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_B1;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_B2;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_B3;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_B4;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_B5;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_B6;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_BO5;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_BO6;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_B_CY;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_B_XOR;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_C;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_C1;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_C2;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_C3;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_C4;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_C5;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_C6;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_CLK;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_CO5;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_CO6;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_C_CY;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_C_XOR;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_D;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_D1;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_D2;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_D3;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_D4;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_D5;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_D6;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_DO5;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_DO6;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_D_CY;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_D_XOR;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X162Y69_SR;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_A;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_A1;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_A2;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_A3;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_A4;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_A5;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_A6;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_AO5;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_AO6;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_AQ;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_AX;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_A_CY;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_A_XOR;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_B;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_B1;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_B2;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_B3;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_B4;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_B5;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_B6;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_BO5;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_BO6;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_B_CY;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_B_XOR;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_C;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_C1;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_C2;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_C3;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_C4;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_C5;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_C6;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_CLK;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_CO5;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_CO6;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_C_CY;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_C_XOR;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_D;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_D1;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_D2;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_D3;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_D4;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_D5;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_D6;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_DO5;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_DO6;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_D_CY;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_D_XOR;
  wire [0:0] CLBLM_R_X103Y69_SLICE_X163Y69_SR;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_A;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_A1;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_A2;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_A3;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_A4;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_A5;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_A6;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_AO5;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_AO6;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_AQ;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_AX;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_A_CY;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_A_XOR;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_B;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_B1;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_B2;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_B3;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_B4;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_B5;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_B6;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_BO5;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_BO6;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_BQ;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_BX;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_B_CY;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_B_XOR;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_C;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_C1;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_C2;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_C3;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_C4;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_C5;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_C6;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_CLK;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_CO5;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_CO6;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_CQ;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_CX;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_C_CY;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_C_XOR;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_D;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_D1;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_D2;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_D3;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_D4;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_D5;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_D6;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_DO5;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_DO6;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_D_CY;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_D_XOR;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X162Y75_SR;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_A;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_A1;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_A2;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_A3;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_A4;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_A5;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_A6;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_AO5;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_AO6;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_AQ;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_AX;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_A_CY;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_A_XOR;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_B;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_B1;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_B2;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_B3;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_B4;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_B5;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_B6;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_BO5;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_BO6;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_BQ;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_BX;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_B_CY;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_B_XOR;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_C;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_C1;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_C2;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_C3;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_C4;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_C5;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_C6;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_CLK;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_CO5;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_CO6;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_C_CY;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_C_XOR;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_D;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_D1;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_D2;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_D3;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_D4;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_D5;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_D6;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_DO5;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_DO6;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_D_CY;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_D_XOR;
  wire [0:0] CLBLM_R_X103Y75_SLICE_X163Y75_SR;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_A;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_A1;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_A2;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_A3;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_A4;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_A5;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_A6;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_AO5;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_AO6;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_AQ;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_AX;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_A_CY;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_A_XOR;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_B;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_B1;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_B2;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_B3;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_B4;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_B5;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_B6;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_BO5;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_BO6;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_BQ;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_BX;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_B_CY;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_B_XOR;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_C;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_C1;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_C2;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_C3;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_C4;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_C5;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_C6;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_CLK;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_CO5;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_CO6;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_C_CY;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_C_XOR;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_D;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_D1;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_D2;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_D3;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_D4;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_D5;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_D6;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_DO5;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_DO6;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_D_CY;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_D_XOR;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X162Y76_SR;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_A;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_A1;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_A2;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_A3;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_A4;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_A5;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_A6;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_AO5;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_AO6;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_AQ;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_AX;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_A_CY;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_A_XOR;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_B;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_B1;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_B2;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_B3;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_B4;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_B5;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_B6;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_BO5;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_BO6;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_B_CY;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_B_XOR;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_C;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_C1;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_C2;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_C3;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_C4;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_C5;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_C6;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_CLK;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_CO5;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_CO6;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_C_CY;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_C_XOR;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_D;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_D1;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_D2;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_D3;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_D4;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_D5;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_D6;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_DO5;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_DO6;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_D_CY;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_D_XOR;
  wire [0:0] CLBLM_R_X103Y76_SLICE_X163Y76_SR;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_A;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_A1;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_A2;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_A3;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_A4;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_A5;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_A6;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_AO5;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_AO6;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_AQ;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_AX;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_A_CY;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_A_XOR;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_B;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_B1;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_B2;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_B3;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_B4;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_B5;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_B6;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_BO5;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_BO6;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_B_CY;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_B_XOR;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_C;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_C1;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_C2;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_C3;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_C4;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_C5;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_C6;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_CE;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_CLK;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_CO5;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_CO6;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_C_CY;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_C_XOR;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_D;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_D1;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_D2;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_D3;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_D4;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_D5;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_D6;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_DO5;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_DO6;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_D_CY;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_D_XOR;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X80Y122_SR;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_A;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_A1;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_A2;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_A3;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_A4;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_A5;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_A6;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_AO5;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_AO6;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_A_CY;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_A_XOR;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_B;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_B1;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_B2;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_B3;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_B4;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_B5;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_B6;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_BO5;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_BO6;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_B_CY;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_B_XOR;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_C;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_C1;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_C2;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_C3;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_C4;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_C5;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_C6;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_CO5;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_CO6;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_C_CY;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_C_XOR;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_D;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_D1;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_D2;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_D3;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_D4;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_D5;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_D6;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_DO5;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_DO6;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_D_CY;
  wire [0:0] CLBLM_R_X53Y122_SLICE_X81Y122_D_XOR;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_A;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_A1;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_A2;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_A3;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_A4;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_A5;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_A6;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_AMUX;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_AO5;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_AO6;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_AQ;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_AX;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_A_CY;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_A_XOR;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_B;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_B1;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_B2;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_B3;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_B4;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_B5;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_B6;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_BMUX;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_BO5;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_BO6;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_BQ;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_BX;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_B_CY;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_B_XOR;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_C;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_C1;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_C2;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_C3;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_C4;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_C5;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_C6;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_CLK;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_CO5;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_CO6;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_C_CY;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_C_XOR;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_D;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_D1;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_D2;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_D3;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_D4;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_D5;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_D6;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_DO5;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_DO6;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_D_CY;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_D_XOR;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_SR;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_A;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_A1;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_A2;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_A3;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_A4;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_A5;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_A6;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_AO5;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_AO6;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_A_CY;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_A_XOR;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_B;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_B1;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_B2;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_B3;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_B4;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_B5;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_B6;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_BO5;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_BO6;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_B_CY;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_B_XOR;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_C;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_C1;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_C2;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_C3;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_C4;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_C5;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_C6;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_CO5;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_CO6;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_C_CY;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_C_XOR;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_D;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_D1;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_D2;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_D3;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_D4;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_D5;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_D6;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_DO5;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_DO6;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_D_CY;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_D_XOR;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_A;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_A1;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_A2;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_A3;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_A4;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_A5;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_A6;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_AO5;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_AO6;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_AQ;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_A_CY;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_A_XOR;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_B;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_B1;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_B2;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_B3;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_B4;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_B5;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_B6;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_BO5;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_BO6;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_BQ;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_B_CY;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_B_XOR;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_C;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_C1;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_C2;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_C3;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_C4;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_C5;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_C6;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_CLK;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_CO5;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_CO6;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_C_CY;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_C_XOR;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_D;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_D1;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_D2;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_D3;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_D4;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_D5;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_D6;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_DMUX;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_DO5;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_DO6;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_D_CY;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_D_XOR;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_SR;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_A;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_A1;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_A2;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_A3;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_A4;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_A5;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_A6;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_AMUX;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_AO5;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_AO6;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_AQ;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_A_CY;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_A_XOR;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_B;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_B1;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_B2;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_B3;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_B4;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_B5;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_B6;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_BO5;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_BO6;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_BQ;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_B_CY;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_B_XOR;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_C;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_C1;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_C2;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_C3;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_C4;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_C5;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_C6;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_CLK;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_CO5;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_CO6;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_CQ;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_C_CY;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_C_XOR;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_D;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_D1;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_D2;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_D3;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_D4;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_D5;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_D6;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_DO5;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_DO6;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_DQ;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_D_CY;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_D_XOR;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_SR;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_A;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_A1;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_A2;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_A3;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_A4;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_A5;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_A6;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_AMUX;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_AO5;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_AO6;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_AQ;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_AX;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_A_CY;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_A_XOR;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_B;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_B1;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_B2;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_B3;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_B4;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_B5;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_B6;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_BO5;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_BO6;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_B_CY;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_B_XOR;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_C;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_C1;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_C2;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_C3;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_C4;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_C5;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_C6;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_CLK;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_CO5;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_CO6;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_C_CY;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_C_XOR;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_D;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_D1;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_D2;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_D3;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_D4;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_D5;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_D6;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_DO5;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_DO6;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_D_CY;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_D_XOR;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_SR;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_A;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_A1;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_A2;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_A3;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_A4;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_A5;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_A6;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_AO5;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_AO6;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_AQ;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_A_CY;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_A_XOR;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_B;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_B1;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_B2;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_B3;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_B4;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_B5;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_B6;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_BMUX;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_BO5;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_BO6;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_B_CY;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_B_XOR;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_C;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_C1;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_C2;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_C3;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_C4;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_C5;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_C6;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_CLK;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_CO5;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_CO6;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_C_CY;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_C_XOR;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_D;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_D1;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_D2;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_D3;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_D4;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_D5;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_D6;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_DO5;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_DO6;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_D_CY;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_D_XOR;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_SR;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_A;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_A1;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_A2;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_A3;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_A4;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_A5;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_A6;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_AO5;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_AO6;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_AQ;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_A_CY;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_A_XOR;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_B;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_B1;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_B2;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_B3;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_B4;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_B5;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_B6;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_BO5;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_BO6;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_BQ;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_B_CY;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_B_XOR;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_C;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_C1;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_C2;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_C3;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_C4;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_C5;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_C5Q;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_C6;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_CLK;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_CMUX;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_CO5;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_CO6;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_CQ;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_C_CY;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_C_XOR;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_D;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_D1;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_D2;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_D3;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_D4;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_D5;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_D6;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_DO5;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_DO6;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_D_CY;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_D_XOR;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_SR;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_A;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_A1;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_A2;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_A3;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_A4;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_A5;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_A5Q;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_A6;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_AMUX;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_AO5;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_AO6;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_AQ;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_A_CY;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_A_XOR;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_B;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_B1;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_B2;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_B3;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_B4;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_B5;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_B6;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_BO5;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_BO6;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_BQ;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_B_CY;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_B_XOR;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_C;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_C1;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_C2;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_C3;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_C4;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_C5;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_C5Q;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_C6;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_CLK;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_CMUX;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_CO5;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_CO6;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_CQ;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_C_CY;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_C_XOR;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_D;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_D1;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_D2;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_D3;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_D4;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_D5;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_D6;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_DO5;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_DO6;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_D_CY;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_D_XOR;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_SR;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_A;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_A1;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_A2;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_A3;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_A4;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_A5;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_A6;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_AMUX;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_AO5;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_AO6;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_A_CY;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_A_XOR;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_B;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_B1;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_B2;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_B3;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_B4;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_B5;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_B6;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_BO5;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_BO6;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_BQ;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_B_CY;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_B_XOR;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_C;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_C1;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_C2;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_C3;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_C4;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_C5;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_C6;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_CLK;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_CO5;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_CO6;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_C_CY;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_C_XOR;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_D;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_D1;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_D2;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_D3;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_D4;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_D5;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_D6;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_DO5;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_DO6;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_D_CY;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_D_XOR;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_SR;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_A;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_A1;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_A2;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_A3;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_A4;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_A5;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_A6;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_AO5;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_AO6;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_AQ;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_A_CY;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_A_XOR;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_B;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_B1;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_B2;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_B3;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_B4;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_B5;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_B6;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_BO5;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_BO6;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_BQ;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_B_CY;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_B_XOR;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_C;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_C1;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_C2;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_C3;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_C4;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_C5;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_C6;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_CLK;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_CO5;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_CO6;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_CQ;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_C_CY;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_C_XOR;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_D;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_D1;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_D2;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_D3;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_D4;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_D5;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_D6;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_DMUX;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_DO5;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_DO6;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_D_CY;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_D_XOR;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_SR;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_A;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_A1;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_A2;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_A3;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_A4;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_A5;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_A6;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_AO5;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_AO6;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_AQ;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_A_CY;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_A_XOR;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_B;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_B1;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_B2;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_B3;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_B4;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_B5;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_B6;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_BO5;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_BO6;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_BQ;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_B_CY;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_B_XOR;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_C;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_C1;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_C2;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_C3;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_C4;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_C5;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_C6;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_CLK;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_CMUX;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_CO5;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_CO6;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_C_CY;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_C_XOR;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_D;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_D1;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_D2;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_D3;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_D4;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_D5;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_D6;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_DO5;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_DO6;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_D_CY;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_D_XOR;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_SR;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_A;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_A1;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_A2;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_A3;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_A4;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_A5;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_A6;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_AO5;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_AO6;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_AQ;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_A_CY;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_A_XOR;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_B;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_B1;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_B2;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_B3;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_B4;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_B5;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_B6;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_BO5;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_BO6;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_BQ;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_B_CY;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_B_XOR;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_C;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_C1;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_C2;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_C3;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_C4;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_C5;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_C6;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_CLK;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_CO5;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_CO6;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_CQ;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_C_CY;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_C_XOR;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_D;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_D1;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_D2;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_D3;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_D4;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_D5;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_D6;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_DO5;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_DO6;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_DQ;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_D_CY;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_D_XOR;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_SR;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_A;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_A1;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_A2;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_A3;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_A4;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_A5;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_A6;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_AO5;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_AO6;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_A_CY;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_A_XOR;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_B;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_B1;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_B2;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_B3;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_B4;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_B5;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_B6;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_BO5;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_BO6;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_B_CY;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_B_XOR;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_C;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_C1;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_C2;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_C3;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_C4;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_C5;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_C6;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_CO5;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_CO6;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_C_CY;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_C_XOR;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_D;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_D1;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_D2;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_D3;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_D4;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_D5;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_D6;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_DO5;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_DO6;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_D_CY;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X94Y122_D_XOR;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_A;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_A1;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_A2;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_A3;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_A4;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_A5;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_A6;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_AO5;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_AO6;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_AQ;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_AX;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_A_CY;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_A_XOR;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_B;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_B1;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_B2;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_B3;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_B4;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_B5;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_B6;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_BO5;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_BO6;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_B_CY;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_B_XOR;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_C;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_C1;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_C2;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_C3;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_C4;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_C5;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_C6;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_CE;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_CLK;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_CO5;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_CO6;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_CQ;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_CX;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_C_CY;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_C_XOR;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_D;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_D1;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_D2;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_D3;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_D4;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_D5;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_D6;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_DO5;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_DO6;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_D_CY;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_D_XOR;
  wire [0:0] CLBLM_R_X63Y122_SLICE_X95Y122_SR;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_A;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_A1;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_A2;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_A3;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_A4;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_A5;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_A6;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_AO5;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_AO6;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_AQ;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_A_CY;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_A_XOR;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_B;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_B1;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_B2;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_B3;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_B4;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_B5;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_B6;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_BO5;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_BO6;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_BQ;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_B_CY;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_B_XOR;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_C;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_C1;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_C2;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_C3;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_C4;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_C5;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_C6;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_CLK;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_CO5;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_CO6;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_C_CY;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_C_XOR;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_D;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_D1;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_D2;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_D3;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_D4;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_D5;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_D6;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_DO5;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_DO6;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_D_CY;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_D_XOR;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_SR;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_A;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_A1;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_A2;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_A3;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_A4;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_A5;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_A6;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_AO5;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_AO6;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_AQ;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_A_CY;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_A_XOR;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_B;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_B1;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_B2;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_B3;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_B4;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_B5;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_B6;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_BO5;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_BO6;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_BQ;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_B_CY;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_B_XOR;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_C;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_C1;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_C2;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_C3;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_C4;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_C5;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_C6;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_CLK;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_CO5;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_CO6;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_CQ;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_C_CY;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_C_XOR;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_D;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_D1;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_D2;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_D3;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_D4;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_D5;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_D6;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_DO5;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_DO6;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_DQ;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_D_CY;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_D_XOR;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_SR;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_A;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_A1;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_A2;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_A3;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_A4;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_A5;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_A6;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_AMUX;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_AO5;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_AO6;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_AQ;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_AX;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_A_CY;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_A_XOR;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_B;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_B1;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_B2;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_B3;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_B4;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_B5;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_B5Q;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_B6;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_BMUX;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_BO5;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_BO6;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_BQ;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_BX;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_B_CY;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_B_XOR;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_C;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_C1;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_C2;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_C3;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_C4;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_C5;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_C6;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_CLK;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_CO5;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_CO6;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_CQ;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_CX;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_C_CY;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_C_XOR;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_D;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_D1;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_D2;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_D3;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_D4;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_D5;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_D6;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_DO5;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_DO6;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_D_CY;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_D_XOR;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_SR;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_A;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_A1;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_A2;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_A3;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_A4;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_A5;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_A6;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_AO5;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_AO6;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_AQ;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_AX;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_A_CY;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_A_XOR;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_B;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_B1;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_B2;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_B3;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_B4;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_B5;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_B6;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_BMUX;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_BO5;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_BO6;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_B_CY;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_B_XOR;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_C;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_C1;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_C2;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_C3;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_C4;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_C5;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_C6;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_CLK;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_CO5;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_CO6;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_C_CY;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_C_XOR;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_D;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_D1;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_D2;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_D3;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_D4;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_D5;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_D6;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_DO5;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_DO6;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_D_CY;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_D_XOR;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_SR;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_A;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_A1;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_A2;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_A3;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_A4;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_A5;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_A6;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_AMUX;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_AO5;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_AO6;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_AQ;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_AX;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_A_CY;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_A_XOR;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_B;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_B1;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_B2;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_B3;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_B4;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_B5;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_B6;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_BMUX;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_BO5;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_BO6;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_BQ;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_BX;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_B_CY;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_B_XOR;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_C;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_C1;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_C2;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_C3;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_C4;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_C5;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_C6;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_CLK;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_CMUX;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_CO5;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_CO6;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_C_CY;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_C_XOR;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_D;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_D1;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_D2;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_D3;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_D4;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_D5;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_D6;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_DMUX;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_DO5;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_DO6;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_D_CY;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_D_XOR;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_SR;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_A;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_A1;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_A2;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_A3;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_A4;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_A5;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_A6;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_AO5;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_AO6;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_A_CY;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_A_XOR;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_B;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_B1;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_B2;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_B3;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_B4;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_B5;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_B6;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_BO5;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_BO6;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_B_CY;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_B_XOR;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_C;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_C1;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_C2;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_C3;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_C4;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_C5;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_C6;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_CO5;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_CO6;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_C_CY;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_C_XOR;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_D;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_D1;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_D2;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_D3;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_D4;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_D5;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_D6;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_DO5;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_DO6;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_D_CY;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_D_XOR;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_A;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_A1;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_A2;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_A3;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_A4;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_A5;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_A5Q;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_A6;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_AMUX;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_AO5;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_AO6;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_AQ;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_A_CY;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_A_XOR;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_B;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_B1;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_B2;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_B3;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_B4;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_B5;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_B6;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_BMUX;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_BO5;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_BO6;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_B_CY;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_B_XOR;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_C;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_C1;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_C2;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_C3;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_C4;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_C5;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_C6;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_CLK;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_CMUX;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_CO5;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_CO6;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_C_CY;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_C_XOR;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_D;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_D1;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_D2;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_D3;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_D4;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_D5;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_D5Q;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_D6;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_DMUX;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_DO5;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_DO6;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_DQ;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_D_CY;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_D_XOR;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_SR;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_A;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_A1;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_A2;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_A3;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_A4;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_A5;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_A6;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_AMUX;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_AO5;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_AO6;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_A_CY;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_A_XOR;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_B;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_B1;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_B2;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_B3;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_B4;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_B5;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_B5Q;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_B6;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_BMUX;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_BO5;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_BO6;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_BQ;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_B_CY;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_B_XOR;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_C;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_C1;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_C2;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_C3;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_C4;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_C5;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_C6;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_CLK;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_CMUX;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_CO5;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_CO6;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_C_CY;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_C_XOR;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_D;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_D1;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_D2;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_D3;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_D4;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_D5;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_D6;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_DO5;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_DO6;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_D_CY;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_D_XOR;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_SR;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_A;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_A1;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_A2;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_A3;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_A4;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_A5;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_A6;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_AO5;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_AO6;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_AQ;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_A_CY;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_A_XOR;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_B;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_B1;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_B2;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_B3;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_B4;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_B5;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_B6;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_BO5;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_BO6;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_BQ;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_B_CY;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_B_XOR;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_C;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_C1;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_C2;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_C3;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_C4;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_C5;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_C6;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_CLK;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_CO5;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_CO6;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_C_CY;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_C_XOR;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_D;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_D1;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_D2;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_D3;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_D4;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_D5;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_D6;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_DO5;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_DO6;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_D_CY;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_D_XOR;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_SR;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_A;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_A1;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_A2;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_A3;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_A4;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_A5;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_A5Q;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_A6;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_AMUX;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_AO5;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_AO6;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_AQ;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_A_CY;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_A_XOR;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_B;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_B1;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_B2;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_B3;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_B4;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_B5;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_B6;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_BO5;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_BO6;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_BQ;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_B_CY;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_B_XOR;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_C;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_C1;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_C2;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_C3;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_C4;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_C5;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_C6;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_CLK;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_CO5;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_CO6;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_CQ;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_C_CY;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_C_XOR;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_D;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_D1;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_D2;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_D3;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_D4;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_D5;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_D6;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_DO5;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_DO6;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_D_CY;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_D_XOR;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_SR;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_A;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_A1;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_A2;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_A3;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_A4;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_A5;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_A6;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_AO5;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_AO6;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_A_CY;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_A_XOR;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_B;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_B1;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_B2;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_B3;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_B4;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_B5;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_B6;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_BO5;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_BO6;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_B_CY;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_B_XOR;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_C;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_C1;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_C2;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_C3;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_C4;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_C5;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_C6;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_CO5;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_CO6;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_C_CY;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_C_XOR;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_D;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_D1;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_D2;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_D3;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_D4;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_D5;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_D6;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_DO5;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_DO6;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_D_CY;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_D_XOR;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_A;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_A1;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_A2;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_A3;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_A4;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_A5;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_A6;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_AO5;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_AO6;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_AQ;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_A_CY;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_A_XOR;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_B;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_B1;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_B2;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_B3;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_B4;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_B5;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_B6;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_BO5;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_BO6;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_B_CY;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_B_XOR;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_C;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_C1;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_C2;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_C3;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_C4;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_C5;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_C6;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_CLK;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_CO5;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_CO6;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_C_CY;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_C_XOR;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_D;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_D1;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_D2;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_D3;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_D4;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_D5;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_D6;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_DO5;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_DO6;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_D_CY;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_D_XOR;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_SR;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_A;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_A1;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_A2;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_A3;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_A4;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_A5;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_A6;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_AO5;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_AO6;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_A_CY;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_A_XOR;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_B;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_B1;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_B2;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_B3;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_B4;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_B5;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_B6;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_BO5;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_BO6;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_B_CY;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_B_XOR;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_C;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_C1;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_C2;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_C3;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_C4;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_C5;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_C6;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_CO5;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_CO6;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_C_CY;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_C_XOR;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_D;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_D1;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_D2;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_D3;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_D4;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_D5;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_D6;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_DO5;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_DO6;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_D_CY;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_D_XOR;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_A;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_A1;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_A2;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_A3;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_A4;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_A5;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_A6;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_AO5;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_AO6;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_AQ;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_A_CY;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_A_XOR;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_B;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_B1;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_B2;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_B3;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_B4;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_B5;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_B6;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_BO5;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_BO6;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_B_CY;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_B_XOR;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_C;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_C1;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_C2;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_C3;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_C4;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_C5;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_C6;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_CLK;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_CO5;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_CO6;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_C_CY;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_C_XOR;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_D;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_D1;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_D2;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_D3;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_D4;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_D5;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_D6;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_DO5;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_DO6;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_D_CY;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_D_XOR;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_SR;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_A;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_A1;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_A2;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_A3;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_A4;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_A5;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_A5Q;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_A6;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_AMUX;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_AO5;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_AO6;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_AQ;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_AX;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_A_CY;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_A_XOR;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_B;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_B1;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_B2;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_B3;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_B4;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_B5;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_B6;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_BO5;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_BO6;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_BQ;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_B_CY;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_B_XOR;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_C;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_C1;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_C2;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_C3;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_C4;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_C5;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_C6;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_CLK;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_CO5;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_CO6;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_C_CY;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_C_XOR;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_D;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_D1;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_D2;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_D3;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_D4;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_D5;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_D6;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_DO5;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_DO6;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_D_CY;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_D_XOR;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_SR;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_A;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_A1;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_A2;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_A3;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_A4;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_A5;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_A6;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_AO5;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_AO6;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_AQ;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_A_CY;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_A_XOR;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_B;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_B1;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_B2;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_B3;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_B4;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_B5;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_B6;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_BO5;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_BO6;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_BQ;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_B_CY;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_B_XOR;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_C;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_C1;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_C2;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_C3;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_C4;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_C5;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_C6;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_CLK;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_CO5;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_CO6;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_C_CY;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_C_XOR;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_D;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_D1;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_D2;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_D3;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_D4;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_D5;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_D6;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_DMUX;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_DO5;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_DO6;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_D_CY;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_D_XOR;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_SR;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_A;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_A1;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_A2;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_A3;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_A4;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_A5;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_A6;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_AMUX;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_AO5;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_AO6;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_A_CY;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_A_XOR;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_B;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_B1;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_B2;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_B3;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_B4;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_B5;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_B5Q;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_B6;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_BMUX;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_BO5;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_BO6;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_BQ;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_B_CY;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_B_XOR;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_C;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_C1;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_C2;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_C3;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_C4;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_C5;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_C5Q;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_C6;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_CLK;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_CMUX;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_CO5;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_CO6;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_CQ;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_C_CY;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_C_XOR;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_D;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_D1;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_D2;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_D3;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_D4;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_D5;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_D6;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_DO5;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_DO6;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_D_CY;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_D_XOR;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_SR;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_A;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_A1;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_A2;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_A3;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_A4;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_A5;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_A5Q;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_A6;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_AMUX;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_AO5;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_AO6;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_AQ;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_A_CY;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_A_XOR;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_B;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_B1;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_B2;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_B3;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_B4;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_B5;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_B5Q;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_B6;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_BMUX;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_BO5;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_BO6;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_BQ;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_BX;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_B_CY;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_B_XOR;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_C;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_C1;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_C2;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_C3;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_C4;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_C5;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_C6;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_CLK;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_CO5;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_CO6;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_C_CY;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_C_XOR;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_D;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_D1;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_D2;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_D3;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_D4;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_D5;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_D6;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_DO5;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_DO6;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_D_CY;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_D_XOR;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_SR;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_A;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_A1;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_A2;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_A3;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_A4;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_A5;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_A6;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_AO5;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_AO6;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_AQ;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_A_CY;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_A_XOR;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_B;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_B1;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_B2;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_B3;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_B4;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_B5;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_B5Q;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_B6;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_BMUX;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_BO5;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_BO6;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_BQ;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_BX;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_B_CY;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_B_XOR;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_C;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_C1;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_C2;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_C3;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_C4;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_C5;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_C6;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_CLK;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_CO5;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_CO6;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_CQ;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_C_CY;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_C_XOR;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_D;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_D1;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_D2;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_D3;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_D4;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_D5;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_D6;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_DO5;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_DO6;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_D_CY;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_D_XOR;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_SR;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_A;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_A1;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_A2;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_A3;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_A4;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_A5;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_A6;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_AO5;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_AO6;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_AQ;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_A_CY;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_A_XOR;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_B;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_B1;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_B2;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_B3;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_B4;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_B5;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_B6;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_BMUX;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_BO5;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_BO6;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_B_CY;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_B_XOR;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_C;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_C1;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_C2;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_C3;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_C4;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_C5;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_C5Q;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_C6;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_CLK;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_CMUX;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_CO5;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_CO6;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_CQ;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_C_CY;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_C_XOR;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_D;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_D1;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_D2;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_D3;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_D4;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_D5;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_D5Q;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_D6;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_DMUX;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_DO5;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_DO6;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_DQ;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_D_CY;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_D_XOR;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_SR;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_A;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_A1;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_A2;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_A3;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_A4;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_A5;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_A6;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_AO5;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_AO6;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_AQ;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_A_CY;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_A_XOR;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_B;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_B1;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_B2;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_B3;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_B4;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_B5;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_B6;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_BO5;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_BO6;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_BQ;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_B_CY;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_B_XOR;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_C;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_C1;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_C2;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_C3;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_C4;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_C5;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_C6;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_CLK;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_CO5;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_CO6;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_CQ;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_C_CY;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_C_XOR;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_D;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_D1;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_D2;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_D3;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_D4;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_D5;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_D6;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_DO5;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_DO6;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_DQ;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_D_CY;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_D_XOR;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_SR;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_A;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_A1;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_A2;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_A3;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_A4;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_A5;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_A6;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_AO5;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_AO6;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_AQ;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_A_CY;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_A_XOR;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_B;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_B1;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_B2;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_B3;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_B4;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_B5;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_B6;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_BO5;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_BO6;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_BQ;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_B_CY;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_B_XOR;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_C;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_C1;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_C2;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_C3;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_C4;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_C5;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_C5Q;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_C6;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_CLK;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_CMUX;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_CO5;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_CO6;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_CQ;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_C_CY;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_C_XOR;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_D;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_D1;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_D2;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_D3;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_D4;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_D5;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_D6;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_DO5;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_DO6;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_DQ;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_D_CY;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_D_XOR;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_SR;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_A;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_A1;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_A2;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_A3;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_A4;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_A5;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_A6;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_AO5;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_AO6;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_A_CY;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_A_XOR;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_B;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_B1;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_B2;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_B3;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_B4;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_B5;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_B6;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_BO5;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_BO6;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_B_CY;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_B_XOR;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_C;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_C1;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_C2;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_C3;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_C4;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_C5;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_C6;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_CO5;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_CO6;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_C_CY;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_C_XOR;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_D;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_D1;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_D2;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_D3;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_D4;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_D5;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_D6;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_DO5;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_DO6;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_D_CY;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X98Y108_D_XOR;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_A;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_A1;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_A2;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_A3;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_A4;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_A5;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_A6;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_AO5;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_AO6;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_A_CY;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_A_XOR;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_B;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_B1;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_B2;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_B3;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_B4;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_B5;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_B6;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_BO5;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_BO6;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_B_CY;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_B_XOR;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_C;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_C1;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_C2;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_C3;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_C4;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_C5;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_C6;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_CMUX;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_CO5;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_CO6;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_C_CY;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_C_XOR;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_D;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_D1;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_D2;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_D3;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_D4;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_D5;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_D6;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_DO5;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_DO6;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_D_CY;
  wire [0:0] CLBLM_R_X65Y108_SLICE_X99Y108_D_XOR;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_A;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_A1;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_A2;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_A3;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_A4;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_A5;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_A5Q;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_A6;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_AMUX;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_AO5;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_AO6;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_AQ;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_AX;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_A_CY;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_A_XOR;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_B;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_B1;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_B2;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_B3;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_B4;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_B5;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_B6;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_BO5;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_BO6;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_BQ;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_B_CY;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_B_XOR;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_C;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_C1;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_C2;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_C3;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_C4;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_C5;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_C6;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_CLK;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_CO5;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_CO6;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_CQ;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_C_CY;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_C_XOR;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_D;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_D1;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_D2;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_D3;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_D4;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_D5;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_D6;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_DO5;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_DO6;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_D_CY;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_D_XOR;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X98Y109_SR;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_A;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_A1;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_A2;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_A3;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_A4;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_A5;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_A5Q;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_A6;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_AMUX;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_AO5;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_AO6;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_AQ;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_AX;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_A_CY;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_A_XOR;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_B;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_B1;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_B2;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_B3;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_B4;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_B5;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_B6;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_BO5;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_BO6;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_BQ;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_B_CY;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_B_XOR;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_C;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_C1;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_C2;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_C3;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_C4;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_C5;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_C6;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_CLK;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_CO5;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_CO6;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_CQ;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_C_CY;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_C_XOR;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_D;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_D1;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_D2;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_D3;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_D4;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_D5;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_D6;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_DMUX;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_DO5;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_DO6;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_D_CY;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_D_XOR;
  wire [0:0] CLBLM_R_X65Y109_SLICE_X99Y109_SR;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_A;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_A1;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_A2;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_A3;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_A4;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_A5;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_A5Q;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_A6;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_AMUX;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_AO5;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_AO6;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_AQ;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_AX;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_A_CY;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_A_XOR;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_B;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_B1;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_B2;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_B3;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_B4;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_B5;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_B6;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_BO5;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_BO6;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_BQ;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_B_CY;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_B_XOR;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_C;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_C1;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_C2;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_C3;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_C4;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_C5;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_C6;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_CLK;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_CO5;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_CO6;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_CQ;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_C_CY;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_C_XOR;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_D;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_D1;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_D2;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_D3;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_D4;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_D5;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_D6;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_DO5;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_DO6;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_DQ;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_D_CY;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_D_XOR;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X98Y110_SR;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_A;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_A1;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_A2;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_A3;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_A4;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_A5;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_A6;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_AMUX;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_AO5;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_AO6;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_AQ;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_AX;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_A_CY;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_A_XOR;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_B;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_B1;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_B2;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_B3;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_B4;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_B5;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_B5Q;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_B6;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_BMUX;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_BO5;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_BO6;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_BQ;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_BX;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_B_CY;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_B_XOR;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_C;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_C1;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_C2;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_C3;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_C4;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_C5;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_C6;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_CLK;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_CO5;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_CO6;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_CQ;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_CX;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_C_CY;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_C_XOR;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_D;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_D1;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_D2;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_D3;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_D4;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_D5;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_D6;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_DO5;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_DO6;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_D_CY;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_D_XOR;
  wire [0:0] CLBLM_R_X65Y110_SLICE_X99Y110_SR;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_A;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_A1;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_A2;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_A3;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_A4;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_A5;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_A6;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_AO5;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_AO6;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_AQ;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_A_CY;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_A_XOR;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_B;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_B1;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_B2;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_B3;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_B4;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_B5;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_B6;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_BO5;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_BO6;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_B_CY;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_B_XOR;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_C;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_C1;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_C2;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_C3;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_C4;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_C5;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_C6;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_CLK;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_CO5;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_CO6;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_C_CY;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_C_XOR;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_D;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_D1;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_D2;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_D3;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_D4;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_D5;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_D6;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_DO5;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_DO6;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_D_CY;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_D_XOR;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X98Y111_SR;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_A;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_A1;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_A2;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_A3;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_A4;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_A5;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_A6;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_AMUX;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_AO5;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_AO6;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_A_CY;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_A_XOR;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_B;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_B1;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_B2;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_B3;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_B4;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_B5;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_B6;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_BO5;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_BO6;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_B_CY;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_B_XOR;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_C;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_C1;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_C2;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_C3;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_C4;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_C5;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_C6;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_CO5;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_CO6;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_C_CY;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_C_XOR;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_D;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_D1;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_D2;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_D3;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_D4;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_D5;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_D6;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_DO5;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_DO6;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_D_CY;
  wire [0:0] CLBLM_R_X65Y111_SLICE_X99Y111_D_XOR;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_A;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_A1;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_A2;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_A3;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_A4;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_A5;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_A6;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_AO5;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_AO6;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_AQ;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_A_CY;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_A_XOR;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_B;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_B1;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_B2;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_B3;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_B4;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_B5;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_B6;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_BO5;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_BO6;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_BQ;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_B_CY;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_B_XOR;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_C;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_C1;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_C2;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_C3;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_C4;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_C5;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_C6;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_CLK;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_CO5;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_CO6;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_CQ;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_C_CY;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_C_XOR;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_D;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_D1;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_D2;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_D3;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_D4;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_D5;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_D6;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_DO5;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_DO6;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_D_CY;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_D_XOR;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_SR;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_A;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_A1;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_A2;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_A3;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_A4;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_A5;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_A6;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_AO5;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_AO6;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_AQ;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_A_CY;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_A_XOR;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_B;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_B1;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_B2;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_B3;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_B4;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_B5;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_B6;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_BO5;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_BO6;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_BQ;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_B_CY;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_B_XOR;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_C;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_C1;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_C2;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_C3;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_C4;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_C5;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_C5Q;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_C6;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_CLK;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_CMUX;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_CO5;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_CO6;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_CQ;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_C_CY;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_C_XOR;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_D;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_D1;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_D2;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_D3;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_D4;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_D5;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_D6;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_DO5;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_DO6;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_DQ;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_D_CY;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_D_XOR;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_SR;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_A;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_A1;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_A2;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_A3;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_A4;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_A5;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_A5Q;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_A6;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_AMUX;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_AO5;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_AO6;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_AQ;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_AX;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_A_CY;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_A_XOR;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_B;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_B1;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_B2;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_B3;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_B4;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_B5;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_B6;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_BO5;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_BO6;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_BQ;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_B_CY;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_B_XOR;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_C;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_C1;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_C2;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_C3;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_C4;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_C5;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_C6;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_CLK;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_CO5;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_CO6;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_CQ;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_C_CY;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_C_XOR;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_D;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_D1;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_D2;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_D3;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_D4;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_D5;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_D6;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_DO5;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_DO6;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_D_CY;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_D_XOR;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X100Y100_SR;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_A;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_A1;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_A2;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_A3;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_A4;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_A5;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_A6;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_AO5;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_AO6;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_A_CY;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_A_XOR;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_B;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_B1;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_B2;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_B3;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_B4;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_B5;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_B6;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_BO5;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_BO6;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_B_CY;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_B_XOR;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_C;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_C1;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_C2;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_C3;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_C4;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_C5;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_C6;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_CO5;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_CO6;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_C_CY;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_C_XOR;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_D;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_D1;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_D2;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_D3;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_D4;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_D5;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_D6;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_DO5;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_DO6;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_D_CY;
  wire [0:0] CLBLM_R_X67Y100_SLICE_X101Y100_D_XOR;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_A;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_A1;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_A2;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_A3;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_A4;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_A5;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_A6;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_AO5;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_AO6;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_AQ;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_A_CY;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_A_XOR;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_B;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_B1;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_B2;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_B3;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_B4;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_B5;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_B6;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_BMUX;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_BO5;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_BO6;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_B_CY;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_B_XOR;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_C;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_C1;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_C2;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_C3;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_C4;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_C5;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_C6;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_CLK;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_CO5;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_CO6;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_CQ;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_C_CY;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_C_XOR;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_D;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_D1;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_D2;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_D3;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_D4;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_D5;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_D6;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_DO5;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_DO6;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_D_CY;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_D_XOR;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X100Y101_SR;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_A;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_A1;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_A2;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_A3;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_A4;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_A5;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_A6;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_AO5;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_AO6;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_AQ;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_A_CY;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_A_XOR;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_B;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_B1;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_B2;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_B3;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_B4;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_B5;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_B6;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_BO5;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_BO6;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_BQ;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_B_CY;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_B_XOR;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_C;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_C1;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_C2;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_C3;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_C4;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_C5;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_C6;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_CLK;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_CMUX;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_CO5;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_CO6;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_C_CY;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_C_XOR;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_D;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_D1;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_D2;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_D3;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_D4;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_D5;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_D6;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_DO5;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_DO6;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_D_CY;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_D_XOR;
  wire [0:0] CLBLM_R_X67Y101_SLICE_X101Y101_SR;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_A;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_A1;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_A2;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_A3;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_A4;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_A5;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_A6;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_AMUX;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_AO5;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_AO6;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_AQ;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_AX;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_A_CY;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_A_XOR;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_B;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_B1;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_B2;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_B3;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_B4;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_B5;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_B5Q;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_B6;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_BMUX;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_BO5;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_BO6;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_BQ;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_BX;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_B_CY;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_B_XOR;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_C;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_C1;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_C2;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_C3;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_C4;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_C5;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_C6;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_CLK;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_CO5;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_CO6;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_C_CY;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_C_XOR;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_D;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_D1;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_D2;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_D3;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_D4;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_D5;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_D6;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_DO5;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_DO6;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_D_CY;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_D_XOR;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X100Y103_SR;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_A;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_A1;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_A2;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_A3;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_A4;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_A5;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_A6;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_AO5;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_AO6;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_AQ;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_A_CY;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_A_XOR;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_B;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_B1;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_B2;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_B3;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_B4;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_B5;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_B6;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_BO5;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_BO6;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_B_CY;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_B_XOR;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_C;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_C1;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_C2;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_C3;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_C4;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_C5;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_C6;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_CLK;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_CO5;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_CO6;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_C_CY;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_C_XOR;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_D;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_D1;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_D2;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_D3;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_D4;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_D5;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_D6;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_DO5;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_DO6;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_D_CY;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_D_XOR;
  wire [0:0] CLBLM_R_X67Y103_SLICE_X101Y103_SR;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_A;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_A1;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_A2;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_A3;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_A4;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_A5;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_A6;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_AMUX;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_AO5;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_AO6;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_A_CY;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_A_XOR;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_B;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_B1;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_B2;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_B3;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_B4;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_B5;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_B6;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_BO5;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_BO6;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_B_CY;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_B_XOR;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_C;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_C1;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_C2;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_C3;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_C4;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_C5;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_C6;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_CMUX;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_CO5;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_CO6;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_C_CY;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_C_XOR;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_D;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_D1;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_D2;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_D3;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_D4;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_D5;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_D6;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_DMUX;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_DO5;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_DO6;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_D_CY;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X100Y105_D_XOR;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_A;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_A1;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_A2;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_A3;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_A4;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_A5;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_A6;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_AO5;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_AO6;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_A_CY;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_A_XOR;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_B;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_B1;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_B2;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_B3;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_B4;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_B5;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_B6;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_BO5;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_BO6;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_B_CY;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_B_XOR;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_C;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_C1;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_C2;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_C3;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_C4;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_C5;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_C6;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_CO5;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_CO6;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_C_CY;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_C_XOR;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_D;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_D1;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_D2;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_D3;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_D4;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_D5;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_D6;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_DMUX;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_DO5;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_DO6;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_D_CY;
  wire [0:0] CLBLM_R_X67Y105_SLICE_X101Y105_D_XOR;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_A;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_A1;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_A2;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_A3;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_A4;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_A5;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_A6;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_AO5;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_AO6;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_AQ;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_A_CY;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_A_XOR;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_B;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_B1;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_B2;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_B3;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_B4;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_B5;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_B6;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_BMUX;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_BO5;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_BO6;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_B_CY;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_B_XOR;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_C;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_C1;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_C2;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_C3;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_C4;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_C5;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_C5Q;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_C6;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_CLK;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_CMUX;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_CO5;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_CO6;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_CQ;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_C_CY;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_C_XOR;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_D;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_D1;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_D2;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_D3;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_D4;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_D5;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_D6;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_DO5;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_DO6;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_DQ;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_D_CY;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_D_XOR;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X100Y108_SR;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_A;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_A1;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_A2;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_A3;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_A4;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_A5;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_A6;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_AMUX;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_AO5;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_AO6;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_A_CY;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_A_XOR;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_B;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_B1;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_B2;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_B3;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_B4;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_B5;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_B6;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_BO5;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_BO6;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_BQ;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_B_CY;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_B_XOR;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_C;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_C1;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_C2;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_C3;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_C4;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_C5;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_C6;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_CLK;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_CO5;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_CO6;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_C_CY;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_C_XOR;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_D;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_D1;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_D2;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_D3;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_D4;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_D5;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_D6;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_DO5;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_DO6;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_D_CY;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_D_XOR;
  wire [0:0] CLBLM_R_X67Y108_SLICE_X101Y108_SR;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_A;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_A1;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_A2;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_A3;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_A4;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_A5;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_A6;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_AO5;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_AO6;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_AQ;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_A_CY;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_A_XOR;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_B;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_B1;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_B2;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_B3;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_B4;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_B5;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_B6;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_BO5;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_BO6;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_BQ;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_B_CY;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_B_XOR;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_C;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_C1;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_C2;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_C3;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_C4;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_C5;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_C6;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_CLK;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_CO5;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_CO6;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_CQ;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_C_CY;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_C_XOR;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_D;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_D1;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_D2;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_D3;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_D4;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_D5;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_D6;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_DMUX;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_DO5;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_DO6;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_D_CY;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_D_XOR;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X100Y109_SR;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_A;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_A1;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_A2;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_A3;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_A4;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_A5;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_A6;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_AO5;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_AO6;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_AQ;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_A_CY;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_A_XOR;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_B;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_B1;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_B2;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_B3;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_B4;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_B5;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_B6;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_BO5;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_BO6;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_BQ;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_B_CY;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_B_XOR;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_C;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_C1;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_C2;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_C3;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_C4;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_C5;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_C6;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_CLK;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_CO5;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_CO6;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_C_CY;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_C_XOR;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_D;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_D1;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_D2;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_D3;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_D4;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_D5;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_D6;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_DO5;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_DO6;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_D_CY;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_D_XOR;
  wire [0:0] CLBLM_R_X67Y109_SLICE_X101Y109_SR;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_A;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_A1;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_A2;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_A3;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_A4;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_A5;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_A6;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_AO5;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_AO6;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_AQ;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_A_CY;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_A_XOR;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_B;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_B1;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_B2;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_B3;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_B4;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_B5;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_B6;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_BO5;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_BO6;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_BQ;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_B_CY;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_B_XOR;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_C;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_C1;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_C2;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_C3;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_C4;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_C5;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_C6;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_CLK;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_CO5;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_CO6;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_CQ;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_C_CY;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_C_XOR;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_D;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_D1;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_D2;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_D3;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_D4;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_D5;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_D6;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_DO5;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_DO6;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_D_CY;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_D_XOR;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X100Y110_SR;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_A;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_A1;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_A2;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_A3;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_A4;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_A5;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_A6;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_AO5;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_AO6;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_AQ;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_A_CY;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_A_XOR;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_B;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_B1;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_B2;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_B3;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_B4;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_B5;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_B6;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_BO5;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_BO6;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_BQ;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_B_CY;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_B_XOR;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_C;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_C1;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_C2;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_C3;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_C4;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_C5;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_C6;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_CLK;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_CO5;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_CO6;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_CQ;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_C_CY;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_C_XOR;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_D;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_D1;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_D2;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_D3;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_D4;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_D5;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_D6;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_DO5;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_DO6;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_DQ;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_D_CY;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_D_XOR;
  wire [0:0] CLBLM_R_X67Y110_SLICE_X101Y110_SR;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_A;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_A1;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_A2;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_A3;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_A4;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_A5;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_A5Q;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_A6;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_AMUX;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_AO5;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_AO6;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_AQ;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_AX;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_A_CY;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_A_XOR;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_B;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_B1;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_B2;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_B3;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_B4;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_B5;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_B6;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_BO5;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_BO6;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_BQ;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_B_CY;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_B_XOR;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_C;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_C1;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_C2;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_C3;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_C4;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_C5;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_C6;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_CLK;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_CMUX;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_CO5;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_CO6;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_C_CY;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_C_XOR;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_D;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_D1;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_D2;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_D3;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_D4;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_D5;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_D6;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_DO5;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_DO6;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_D_CY;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_D_XOR;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X100Y111_SR;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_A;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_A1;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_A2;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_A3;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_A4;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_A5;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_A5Q;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_A6;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_AMUX;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_AO5;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_AO6;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_AQ;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_A_CY;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_A_XOR;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_B;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_B1;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_B2;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_B3;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_B4;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_B5;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_B5Q;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_B6;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_BMUX;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_BO5;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_BO6;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_BQ;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_B_CY;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_B_XOR;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_C;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_C1;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_C2;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_C3;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_C4;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_C5;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_C6;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_CLK;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_CMUX;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_CO5;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_CO6;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_C_CY;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_C_XOR;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_D;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_D1;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_D2;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_D3;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_D4;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_D5;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_D6;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_DMUX;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_DO5;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_DO6;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_D_CY;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_D_XOR;
  wire [0:0] CLBLM_R_X67Y111_SLICE_X101Y111_SR;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_A;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_A1;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_A2;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_A3;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_A4;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_A5;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_A5Q;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_A6;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_AMUX;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_AO5;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_AO6;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_AQ;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_A_CY;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_A_XOR;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_B;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_B1;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_B2;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_B3;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_B4;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_B5;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_B6;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_BO5;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_BO6;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_B_CY;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_B_XOR;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_C;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_C1;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_C2;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_C3;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_C4;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_C5;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_C6;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_CLK;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_CO5;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_CO6;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_C_CY;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_C_XOR;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_D;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_D1;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_D2;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_D3;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_D4;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_D5;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_D6;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_DO5;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_DO6;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_D_CY;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_D_XOR;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X100Y115_SR;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_A;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_A1;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_A2;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_A3;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_A4;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_A5;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_A6;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_AO5;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_AO6;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_A_CY;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_A_XOR;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_B;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_B1;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_B2;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_B3;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_B4;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_B5;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_B6;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_BO5;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_BO6;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_B_CY;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_B_XOR;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_C;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_C1;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_C2;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_C3;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_C4;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_C5;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_C6;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_CO5;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_CO6;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_C_CY;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_C_XOR;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_D;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_D1;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_D2;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_D3;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_D4;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_D5;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_D6;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_DO5;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_DO6;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_D_CY;
  wire [0:0] CLBLM_R_X67Y115_SLICE_X101Y115_D_XOR;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_A;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_A1;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_A2;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_A3;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_A4;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_A5;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_A6;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_AO5;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_AO6;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_AQ;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_A_CY;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_A_XOR;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_B;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_B1;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_B2;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_B3;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_B4;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_B5;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_B5Q;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_B6;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_BMUX;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_BO5;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_BO6;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_BQ;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_B_CY;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_B_XOR;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_C;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_C1;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_C2;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_C3;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_C4;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_C5;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_C5Q;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_C6;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_CLK;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_CMUX;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_CO5;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_CO6;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_CQ;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_C_CY;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_C_XOR;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_D;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_D1;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_D2;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_D3;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_D4;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_D5;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_D6;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_DO5;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_DO6;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_D_CY;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_D_XOR;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X100Y116_SR;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_A;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_A1;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_A2;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_A3;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_A4;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_A5;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_A5Q;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_A6;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_AMUX;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_AO5;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_AO6;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_AQ;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_A_CY;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_A_XOR;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_B;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_B1;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_B2;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_B3;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_B4;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_B5;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_B6;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_BO5;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_BO6;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_BQ;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_BX;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_B_CY;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_B_XOR;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_C;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_C1;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_C2;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_C3;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_C4;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_C5;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_C6;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_CLK;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_CO5;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_CO6;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_C_CY;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_C_XOR;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_D;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_D1;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_D2;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_D3;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_D4;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_D5;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_D6;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_DO5;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_DO6;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_D_CY;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_D_XOR;
  wire [0:0] CLBLM_R_X67Y116_SLICE_X101Y116_SR;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_A;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_A1;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_A2;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_A3;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_A4;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_A5;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_A5Q;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_A6;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_AMUX;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_AO5;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_AO6;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_AQ;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_A_CY;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_A_XOR;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_B;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_B1;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_B2;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_B3;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_B4;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_B5;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_B6;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_BO5;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_BO6;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_B_CY;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_B_XOR;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_C;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_C1;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_C2;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_C3;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_C4;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_C5;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_C6;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_CLK;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_CO5;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_CO6;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_C_CY;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_C_XOR;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_D;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_D1;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_D2;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_D3;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_D4;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_D5;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_D6;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_DO5;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_DO6;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_D_CY;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_D_XOR;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X100Y118_SR;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_A;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_A1;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_A2;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_A3;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_A4;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_A5;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_A5Q;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_A6;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_AMUX;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_AO5;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_AO6;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_AQ;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_A_CY;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_A_XOR;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_B;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_B1;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_B2;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_B3;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_B4;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_B5;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_B6;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_BO5;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_BO6;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_BQ;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_BX;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_B_CY;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_B_XOR;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_C;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_C1;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_C2;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_C3;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_C4;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_C5;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_C6;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_CLK;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_CO5;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_CO6;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_C_CY;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_C_XOR;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_D;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_D1;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_D2;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_D3;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_D4;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_D5;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_D6;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_DO5;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_DO6;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_D_CY;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_D_XOR;
  wire [0:0] CLBLM_R_X67Y118_SLICE_X101Y118_SR;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_A;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_A1;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_A2;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_A3;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_A4;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_A5;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_A6;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_AO5;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_AO6;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_A_CY;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_A_XOR;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_B;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_B1;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_B2;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_B3;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_B4;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_B5;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_B6;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_BO5;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_BO6;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_B_CY;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_B_XOR;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_C;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_C1;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_C2;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_C3;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_C4;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_C5;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_C6;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_CO5;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_CO6;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_C_CY;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_C_XOR;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_D;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_D1;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_D2;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_D3;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_D4;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_D5;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_D6;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_DO5;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_DO6;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_D_CY;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X100Y96_D_XOR;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_A;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_A1;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_A2;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_A3;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_A4;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_A5;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_A6;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_AO5;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_AO6;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_AQ;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_A_CY;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_A_XOR;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_B;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_B1;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_B2;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_B3;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_B4;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_B5;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_B6;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_BO5;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_BO6;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_BQ;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_B_CY;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_B_XOR;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_C;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_C1;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_C2;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_C3;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_C4;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_C5;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_C6;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_CLK;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_CO5;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_CO6;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_CQ;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_C_CY;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_C_XOR;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_D;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_D1;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_D2;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_D3;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_D4;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_D5;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_D6;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_DO5;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_DO6;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_DQ;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_D_CY;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_D_XOR;
  wire [0:0] CLBLM_R_X67Y96_SLICE_X101Y96_SR;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_A;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_A1;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_A2;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_A3;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_A4;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_A5;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_A6;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_AO5;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_AO6;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_AQ;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_A_CY;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_A_XOR;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_B;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_B1;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_B2;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_B3;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_B4;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_B5;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_B6;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_BO5;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_BO6;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_B_CY;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_B_XOR;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_C;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_C1;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_C2;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_C3;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_C4;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_C5;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_C6;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_CLK;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_CO5;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_CO6;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_C_CY;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_C_XOR;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_D;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_D1;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_D2;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_D3;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_D4;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_D5;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_D6;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_DO5;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_DO6;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_D_CY;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_D_XOR;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X100Y97_SR;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_A;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_A1;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_A2;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_A3;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_A4;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_A5;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_A6;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_AO5;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_AO6;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_AQ;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_A_CY;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_A_XOR;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_B;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_B1;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_B2;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_B3;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_B4;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_B5;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_B6;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_BO5;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_BO6;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_BQ;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_B_CY;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_B_XOR;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_C;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_C1;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_C2;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_C3;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_C4;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_C5;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_C6;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_CLK;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_CO5;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_CO6;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_CQ;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_C_CY;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_C_XOR;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_D;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_D1;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_D2;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_D3;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_D4;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_D5;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_D6;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_DO5;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_DO6;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_DQ;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_D_CY;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_D_XOR;
  wire [0:0] CLBLM_R_X67Y97_SLICE_X101Y97_SR;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_A;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_A1;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_A2;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_A3;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_A4;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_A5;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_A5Q;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_A6;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_AMUX;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_AO5;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_AO6;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_AQ;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_A_CY;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_A_XOR;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_B;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_B1;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_B2;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_B3;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_B4;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_B5;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_B5Q;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_B6;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_BMUX;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_BO5;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_BO6;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_BQ;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_B_CY;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_B_XOR;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_C;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_C1;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_C2;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_C3;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_C4;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_C5;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_C6;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_CLK;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_CMUX;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_CO5;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_CO6;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_C_CY;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_C_XOR;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_D;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_D1;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_D2;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_D3;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_D4;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_D5;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_D6;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_DO5;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_DO6;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_D_CY;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_D_XOR;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X100Y98_SR;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_A;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_A1;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_A2;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_A3;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_A4;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_A5;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_A6;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_AMUX;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_AO5;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_AO6;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_A_CY;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_A_XOR;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_B;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_B1;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_B2;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_B3;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_B4;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_B5;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_B6;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_BMUX;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_BO5;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_BO6;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_B_CY;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_B_XOR;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_C;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_C1;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_C2;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_C3;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_C4;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_C5;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_C6;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_CLK;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_CMUX;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_CO5;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_CO6;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_C_CY;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_C_XOR;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_D;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_D1;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_D2;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_D3;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_D4;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_D5;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_D6;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_DO5;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_DO6;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_DQ;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_D_CY;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_D_XOR;
  wire [0:0] CLBLM_R_X67Y98_SLICE_X101Y98_SR;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_A;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_A1;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_A2;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_A3;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_A4;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_A5;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_A6;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_AO5;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_AO6;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_AQ;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_A_CY;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_A_XOR;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_B;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_B1;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_B2;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_B3;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_B4;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_B5;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_B6;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_BO5;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_BO6;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_BQ;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_B_CY;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_B_XOR;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_C;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_C1;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_C2;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_C3;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_C4;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_C5;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_C6;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_CLK;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_CO5;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_CO6;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_C_CY;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_C_XOR;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_D;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_D1;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_D2;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_D3;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_D4;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_D5;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_D6;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_DO5;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_DO6;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_D_CY;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_D_XOR;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X100Y99_SR;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_A;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_A1;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_A2;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_A3;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_A4;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_A5;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_A6;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_AO5;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_AO6;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_A_CY;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_A_XOR;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_B;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_B1;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_B2;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_B3;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_B4;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_B5;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_B6;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_BO5;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_BO6;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_B_CY;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_B_XOR;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_C;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_C1;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_C2;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_C3;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_C4;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_C5;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_C6;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_CO5;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_CO6;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_C_CY;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_C_XOR;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_D;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_D1;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_D2;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_D3;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_D4;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_D5;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_D6;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_DO5;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_DO6;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_D_CY;
  wire [0:0] CLBLM_R_X67Y99_SLICE_X101Y99_D_XOR;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_CE;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_I;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  wire [0:0] CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_CE;
  wire [0:0] CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_I;
  wire [0:0] CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_O;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_O;
  wire [0:0] LIOB33_SING_X0Y150_IOB_X0Y150_O;
  wire [0:0] LIOB33_SING_X0Y199_IOB_X0Y199_O;
  wire [0:0] LIOB33_SING_X0Y50_IOB_X0Y50_O;
  wire [0:0] LIOB33_SING_X0Y99_IOB_X0Y99_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_O;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y151_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y152_O;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y153_O;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y154_O;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y155_O;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y156_O;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y157_O;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y158_O;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y159_O;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y160_O;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y161_O;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y162_O;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y163_O;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y164_O;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y165_O;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y166_O;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y167_O;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y168_O;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y169_O;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y170_O;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y171_O;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y172_O;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y173_O;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y174_O;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y175_O;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y176_O;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y177_O;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y178_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y179_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y180_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y181_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y182_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y183_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y184_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y185_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y186_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y187_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y188_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y189_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y190_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y191_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y192_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y193_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y194_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y195_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y196_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y197_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y198_O;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y51_O;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y52_O;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y53_O;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y54_O;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y55_O;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y56_O;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y57_O;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y58_O;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y59_O;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y60_O;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y61_O;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y62_O;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y63_O;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y64_O;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y65_O;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y66_O;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y67_O;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y68_O;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y69_O;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y70_O;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y71_O;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y72_O;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y73_O;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y74_O;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y75_O;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y76_O;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y77_O;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y78_O;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y79_O;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y80_O;
  wire [0:0] LIOB33_X0Y81_IOB_X0Y81_O;
  wire [0:0] LIOB33_X0Y81_IOB_X0Y82_O;
  wire [0:0] LIOB33_X0Y83_IOB_X0Y83_O;
  wire [0:0] LIOB33_X0Y83_IOB_X0Y84_O;
  wire [0:0] LIOB33_X0Y85_IOB_X0Y85_O;
  wire [0:0] LIOB33_X0Y85_IOB_X0Y86_O;
  wire [0:0] LIOB33_X0Y87_IOB_X0Y87_O;
  wire [0:0] LIOB33_X0Y87_IOB_X0Y88_O;
  wire [0:0] LIOB33_X0Y89_IOB_X0Y89_O;
  wire [0:0] LIOB33_X0Y89_IOB_X0Y90_O;
  wire [0:0] LIOB33_X0Y91_IOB_X0Y91_O;
  wire [0:0] LIOB33_X0Y91_IOB_X0Y92_O;
  wire [0:0] LIOB33_X0Y93_IOB_X0Y93_O;
  wire [0:0] LIOB33_X0Y93_IOB_X0Y94_O;
  wire [0:0] LIOB33_X0Y95_IOB_X0Y95_O;
  wire [0:0] LIOB33_X0Y95_IOB_X0Y96_O;
  wire [0:0] LIOB33_X0Y97_IOB_X0Y97_O;
  wire [0:0] LIOB33_X0Y97_IOB_X0Y98_O;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ;
  wire [0:0] LIOI3_SING_X0Y50_OLOGIC_X0Y50_D1;
  wire [0:0] LIOI3_SING_X0Y50_OLOGIC_X0Y50_OQ;
  wire [0:0] LIOI3_SING_X0Y50_OLOGIC_X0Y50_T1;
  wire [0:0] LIOI3_SING_X0Y50_OLOGIC_X0Y50_TQ;
  wire [0:0] LIOI3_SING_X0Y99_OLOGIC_X0Y99_D1;
  wire [0:0] LIOI3_SING_X0Y99_OLOGIC_X0Y99_OQ;
  wire [0:0] LIOI3_SING_X0Y99_OLOGIC_X0Y99_T1;
  wire [0:0] LIOI3_SING_X0Y99_OLOGIC_X0Y99_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y57_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y57_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y57_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y57_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y58_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y58_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y58_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y58_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_OLOGIC_X0Y69_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_OLOGIC_X0Y69_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_OLOGIC_X0Y69_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_OLOGIC_X0Y69_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_OLOGIC_X0Y70_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_OLOGIC_X0Y70_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_OLOGIC_X0Y70_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_OLOGIC_X0Y70_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y81_OLOGIC_X0Y81_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y81_OLOGIC_X0Y81_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y81_OLOGIC_X0Y81_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y81_OLOGIC_X0Y81_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y81_OLOGIC_X0Y82_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y81_OLOGIC_X0Y82_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y81_OLOGIC_X0Y82_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y81_OLOGIC_X0Y82_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y93_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y93_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y93_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y93_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y94_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y94_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y94_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y94_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y63_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y63_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y63_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y63_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y87_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y87_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y87_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y87_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y88_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y88_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y88_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y88_TQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_TQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_TQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_D1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_OQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_T1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_TQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_D1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_OQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_T1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_TQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_D1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_OQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_T1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_TQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_D1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_OQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_T1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_TQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_D1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_OQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_T1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_TQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_D1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_OQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_T1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_TQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_D1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_OQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_T1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_TQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_D1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_OQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_T1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_TQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_D1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_OQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_T1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_TQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_D1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_OQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_T1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_TQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_D1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_OQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_T1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_TQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_D1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_OQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_T1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_TQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_D1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_OQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_T1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_TQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_D1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_OQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_T1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_TQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_D1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_OQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_T1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_TQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_D1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_OQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_T1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_TQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_D1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_OQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_T1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_TQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_D1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_OQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_T1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_TQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_TQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_TQ;
  wire [0:0] LIOI3_X0Y51_OLOGIC_X0Y51_D1;
  wire [0:0] LIOI3_X0Y51_OLOGIC_X0Y51_OQ;
  wire [0:0] LIOI3_X0Y51_OLOGIC_X0Y51_T1;
  wire [0:0] LIOI3_X0Y51_OLOGIC_X0Y51_TQ;
  wire [0:0] LIOI3_X0Y51_OLOGIC_X0Y52_D1;
  wire [0:0] LIOI3_X0Y51_OLOGIC_X0Y52_OQ;
  wire [0:0] LIOI3_X0Y51_OLOGIC_X0Y52_T1;
  wire [0:0] LIOI3_X0Y51_OLOGIC_X0Y52_TQ;
  wire [0:0] LIOI3_X0Y53_OLOGIC_X0Y53_D1;
  wire [0:0] LIOI3_X0Y53_OLOGIC_X0Y53_OQ;
  wire [0:0] LIOI3_X0Y53_OLOGIC_X0Y53_T1;
  wire [0:0] LIOI3_X0Y53_OLOGIC_X0Y53_TQ;
  wire [0:0] LIOI3_X0Y53_OLOGIC_X0Y54_D1;
  wire [0:0] LIOI3_X0Y53_OLOGIC_X0Y54_OQ;
  wire [0:0] LIOI3_X0Y53_OLOGIC_X0Y54_T1;
  wire [0:0] LIOI3_X0Y53_OLOGIC_X0Y54_TQ;
  wire [0:0] LIOI3_X0Y55_OLOGIC_X0Y55_D1;
  wire [0:0] LIOI3_X0Y55_OLOGIC_X0Y55_OQ;
  wire [0:0] LIOI3_X0Y55_OLOGIC_X0Y55_T1;
  wire [0:0] LIOI3_X0Y55_OLOGIC_X0Y55_TQ;
  wire [0:0] LIOI3_X0Y55_OLOGIC_X0Y56_D1;
  wire [0:0] LIOI3_X0Y55_OLOGIC_X0Y56_OQ;
  wire [0:0] LIOI3_X0Y55_OLOGIC_X0Y56_T1;
  wire [0:0] LIOI3_X0Y55_OLOGIC_X0Y56_TQ;
  wire [0:0] LIOI3_X0Y59_OLOGIC_X0Y59_D1;
  wire [0:0] LIOI3_X0Y59_OLOGIC_X0Y59_OQ;
  wire [0:0] LIOI3_X0Y59_OLOGIC_X0Y59_T1;
  wire [0:0] LIOI3_X0Y59_OLOGIC_X0Y59_TQ;
  wire [0:0] LIOI3_X0Y59_OLOGIC_X0Y60_D1;
  wire [0:0] LIOI3_X0Y59_OLOGIC_X0Y60_OQ;
  wire [0:0] LIOI3_X0Y59_OLOGIC_X0Y60_T1;
  wire [0:0] LIOI3_X0Y59_OLOGIC_X0Y60_TQ;
  wire [0:0] LIOI3_X0Y61_OLOGIC_X0Y61_D1;
  wire [0:0] LIOI3_X0Y61_OLOGIC_X0Y61_OQ;
  wire [0:0] LIOI3_X0Y61_OLOGIC_X0Y61_T1;
  wire [0:0] LIOI3_X0Y61_OLOGIC_X0Y61_TQ;
  wire [0:0] LIOI3_X0Y61_OLOGIC_X0Y62_D1;
  wire [0:0] LIOI3_X0Y61_OLOGIC_X0Y62_OQ;
  wire [0:0] LIOI3_X0Y61_OLOGIC_X0Y62_T1;
  wire [0:0] LIOI3_X0Y61_OLOGIC_X0Y62_TQ;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y65_D1;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y65_OQ;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y65_T1;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y65_TQ;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y66_D1;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y66_OQ;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y66_T1;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y66_TQ;
  wire [0:0] LIOI3_X0Y67_OLOGIC_X0Y67_D1;
  wire [0:0] LIOI3_X0Y67_OLOGIC_X0Y67_OQ;
  wire [0:0] LIOI3_X0Y67_OLOGIC_X0Y67_T1;
  wire [0:0] LIOI3_X0Y67_OLOGIC_X0Y67_TQ;
  wire [0:0] LIOI3_X0Y67_OLOGIC_X0Y68_D1;
  wire [0:0] LIOI3_X0Y67_OLOGIC_X0Y68_OQ;
  wire [0:0] LIOI3_X0Y67_OLOGIC_X0Y68_T1;
  wire [0:0] LIOI3_X0Y67_OLOGIC_X0Y68_TQ;
  wire [0:0] LIOI3_X0Y71_OLOGIC_X0Y71_D1;
  wire [0:0] LIOI3_X0Y71_OLOGIC_X0Y71_OQ;
  wire [0:0] LIOI3_X0Y71_OLOGIC_X0Y71_T1;
  wire [0:0] LIOI3_X0Y71_OLOGIC_X0Y71_TQ;
  wire [0:0] LIOI3_X0Y71_OLOGIC_X0Y72_D1;
  wire [0:0] LIOI3_X0Y71_OLOGIC_X0Y72_OQ;
  wire [0:0] LIOI3_X0Y71_OLOGIC_X0Y72_T1;
  wire [0:0] LIOI3_X0Y71_OLOGIC_X0Y72_TQ;
  wire [0:0] LIOI3_X0Y73_OLOGIC_X0Y73_D1;
  wire [0:0] LIOI3_X0Y73_OLOGIC_X0Y73_OQ;
  wire [0:0] LIOI3_X0Y73_OLOGIC_X0Y73_T1;
  wire [0:0] LIOI3_X0Y73_OLOGIC_X0Y73_TQ;
  wire [0:0] LIOI3_X0Y73_OLOGIC_X0Y74_D1;
  wire [0:0] LIOI3_X0Y73_OLOGIC_X0Y74_OQ;
  wire [0:0] LIOI3_X0Y73_OLOGIC_X0Y74_T1;
  wire [0:0] LIOI3_X0Y73_OLOGIC_X0Y74_TQ;
  wire [0:0] LIOI3_X0Y75_OLOGIC_X0Y75_D1;
  wire [0:0] LIOI3_X0Y75_OLOGIC_X0Y75_OQ;
  wire [0:0] LIOI3_X0Y75_OLOGIC_X0Y75_T1;
  wire [0:0] LIOI3_X0Y75_OLOGIC_X0Y75_TQ;
  wire [0:0] LIOI3_X0Y75_OLOGIC_X0Y76_D1;
  wire [0:0] LIOI3_X0Y75_OLOGIC_X0Y76_OQ;
  wire [0:0] LIOI3_X0Y75_OLOGIC_X0Y76_T1;
  wire [0:0] LIOI3_X0Y75_OLOGIC_X0Y76_TQ;
  wire [0:0] LIOI3_X0Y77_OLOGIC_X0Y77_D1;
  wire [0:0] LIOI3_X0Y77_OLOGIC_X0Y77_OQ;
  wire [0:0] LIOI3_X0Y77_OLOGIC_X0Y77_T1;
  wire [0:0] LIOI3_X0Y77_OLOGIC_X0Y77_TQ;
  wire [0:0] LIOI3_X0Y77_OLOGIC_X0Y78_D1;
  wire [0:0] LIOI3_X0Y77_OLOGIC_X0Y78_OQ;
  wire [0:0] LIOI3_X0Y77_OLOGIC_X0Y78_T1;
  wire [0:0] LIOI3_X0Y77_OLOGIC_X0Y78_TQ;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y79_D1;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y79_OQ;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y79_T1;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y79_TQ;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_D1;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_OQ;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_T1;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_TQ;
  wire [0:0] LIOI3_X0Y83_OLOGIC_X0Y83_D1;
  wire [0:0] LIOI3_X0Y83_OLOGIC_X0Y83_OQ;
  wire [0:0] LIOI3_X0Y83_OLOGIC_X0Y83_T1;
  wire [0:0] LIOI3_X0Y83_OLOGIC_X0Y83_TQ;
  wire [0:0] LIOI3_X0Y83_OLOGIC_X0Y84_D1;
  wire [0:0] LIOI3_X0Y83_OLOGIC_X0Y84_OQ;
  wire [0:0] LIOI3_X0Y83_OLOGIC_X0Y84_T1;
  wire [0:0] LIOI3_X0Y83_OLOGIC_X0Y84_TQ;
  wire [0:0] LIOI3_X0Y85_OLOGIC_X0Y85_D1;
  wire [0:0] LIOI3_X0Y85_OLOGIC_X0Y85_OQ;
  wire [0:0] LIOI3_X0Y85_OLOGIC_X0Y85_T1;
  wire [0:0] LIOI3_X0Y85_OLOGIC_X0Y85_TQ;
  wire [0:0] LIOI3_X0Y85_OLOGIC_X0Y86_D1;
  wire [0:0] LIOI3_X0Y85_OLOGIC_X0Y86_OQ;
  wire [0:0] LIOI3_X0Y85_OLOGIC_X0Y86_T1;
  wire [0:0] LIOI3_X0Y85_OLOGIC_X0Y86_TQ;
  wire [0:0] LIOI3_X0Y89_OLOGIC_X0Y89_D1;
  wire [0:0] LIOI3_X0Y89_OLOGIC_X0Y89_OQ;
  wire [0:0] LIOI3_X0Y89_OLOGIC_X0Y89_T1;
  wire [0:0] LIOI3_X0Y89_OLOGIC_X0Y89_TQ;
  wire [0:0] LIOI3_X0Y89_OLOGIC_X0Y90_D1;
  wire [0:0] LIOI3_X0Y89_OLOGIC_X0Y90_OQ;
  wire [0:0] LIOI3_X0Y89_OLOGIC_X0Y90_T1;
  wire [0:0] LIOI3_X0Y89_OLOGIC_X0Y90_TQ;
  wire [0:0] LIOI3_X0Y91_OLOGIC_X0Y91_D1;
  wire [0:0] LIOI3_X0Y91_OLOGIC_X0Y91_OQ;
  wire [0:0] LIOI3_X0Y91_OLOGIC_X0Y91_T1;
  wire [0:0] LIOI3_X0Y91_OLOGIC_X0Y91_TQ;
  wire [0:0] LIOI3_X0Y91_OLOGIC_X0Y92_D1;
  wire [0:0] LIOI3_X0Y91_OLOGIC_X0Y92_OQ;
  wire [0:0] LIOI3_X0Y91_OLOGIC_X0Y92_T1;
  wire [0:0] LIOI3_X0Y91_OLOGIC_X0Y92_TQ;
  wire [0:0] LIOI3_X0Y95_OLOGIC_X0Y95_D1;
  wire [0:0] LIOI3_X0Y95_OLOGIC_X0Y95_OQ;
  wire [0:0] LIOI3_X0Y95_OLOGIC_X0Y95_T1;
  wire [0:0] LIOI3_X0Y95_OLOGIC_X0Y95_TQ;
  wire [0:0] LIOI3_X0Y95_OLOGIC_X0Y96_D1;
  wire [0:0] LIOI3_X0Y95_OLOGIC_X0Y96_OQ;
  wire [0:0] LIOI3_X0Y95_OLOGIC_X0Y96_T1;
  wire [0:0] LIOI3_X0Y95_OLOGIC_X0Y96_TQ;
  wire [0:0] LIOI3_X0Y97_OLOGIC_X0Y97_D1;
  wire [0:0] LIOI3_X0Y97_OLOGIC_X0Y97_OQ;
  wire [0:0] LIOI3_X0Y97_OLOGIC_X0Y97_T1;
  wire [0:0] LIOI3_X0Y97_OLOGIC_X0Y97_TQ;
  wire [0:0] LIOI3_X0Y97_OLOGIC_X0Y98_D1;
  wire [0:0] LIOI3_X0Y97_OLOGIC_X0Y98_OQ;
  wire [0:0] LIOI3_X0Y97_OLOGIC_X0Y98_T1;
  wire [0:0] LIOI3_X0Y97_OLOGIC_X0Y98_TQ;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_O;
  wire [0:0] RIOB33_SING_X105Y149_IOB_X1Y149_O;
  wire [0:0] RIOB33_SING_X105Y150_IOB_X1Y150_O;
  wire [0:0] RIOB33_SING_X105Y199_IOB_X1Y199_O;
  wire [0:0] RIOB33_SING_X105Y50_IOB_X1Y50_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_O;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_O;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_O;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_O;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_O;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_O;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_O;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_O;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_O;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_O;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_O;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_O;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_O;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y114_O;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y115_O;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y116_O;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y117_O;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y118_O;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y119_O;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y120_O;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y121_O;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y122_O;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y123_O;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y124_O;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y125_O;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y126_O;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y127_O;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y128_O;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y129_O;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y130_O;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y131_O;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y132_O;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y133_O;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y134_O;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y135_O;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y136_O;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y137_O;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y138_O;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y139_O;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y140_O;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y141_O;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y142_O;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y143_O;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y144_O;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y145_O;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y146_O;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y147_O;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y148_O;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y151_O;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y152_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y153_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y154_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y155_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y156_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y157_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y158_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y159_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y160_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y161_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y162_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y163_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y164_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y165_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y166_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y167_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y168_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y169_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y170_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y171_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y172_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y173_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y174_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y175_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y176_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y177_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y178_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y179_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y180_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y181_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y182_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y183_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y184_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y185_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y186_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y187_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y188_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y189_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y190_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y191_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y192_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y193_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y194_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y195_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y196_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y197_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y198_O;
  wire [0:0] RIOB33_X105Y51_IOB_X1Y51_I;
  wire [0:0] RIOB33_X105Y51_IOB_X1Y52_I;
  wire [0:0] RIOB33_X105Y53_IOB_X1Y53_I;
  wire [0:0] RIOB33_X105Y53_IOB_X1Y54_I;
  wire [0:0] RIOB33_X105Y55_IOB_X1Y55_I;
  wire [0:0] RIOB33_X105Y55_IOB_X1Y56_I;
  wire [0:0] RIOB33_X105Y57_IOB_X1Y57_I;
  wire [0:0] RIOB33_X105Y57_IOB_X1Y58_I;
  wire [0:0] RIOB33_X105Y59_IOB_X1Y59_I;
  wire [0:0] RIOB33_X105Y59_IOB_X1Y60_I;
  wire [0:0] RIOB33_X105Y61_IOB_X1Y61_I;
  wire [0:0] RIOB33_X105Y61_IOB_X1Y62_I;
  wire [0:0] RIOB33_X105Y63_IOB_X1Y63_O;
  wire [0:0] RIOB33_X105Y63_IOB_X1Y64_O;
  wire [0:0] RIOB33_X105Y65_IOB_X1Y65_O;
  wire [0:0] RIOB33_X105Y65_IOB_X1Y66_O;
  wire [0:0] RIOB33_X105Y67_IOB_X1Y67_O;
  wire [0:0] RIOB33_X105Y67_IOB_X1Y68_O;
  wire [0:0] RIOB33_X105Y69_IOB_X1Y69_O;
  wire [0:0] RIOB33_X105Y69_IOB_X1Y70_O;
  wire [0:0] RIOB33_X105Y71_IOB_X1Y71_O;
  wire [0:0] RIOB33_X105Y71_IOB_X1Y72_O;
  wire [0:0] RIOB33_X105Y73_IOB_X1Y73_O;
  wire [0:0] RIOB33_X105Y73_IOB_X1Y74_O;
  wire [0:0] RIOB33_X105Y75_IOB_X1Y75_O;
  wire [0:0] RIOB33_X105Y75_IOB_X1Y76_O;
  wire [0:0] RIOB33_X105Y77_IOB_X1Y77_O;
  wire [0:0] RIOB33_X105Y77_IOB_X1Y78_I;
  wire [0:0] RIOB33_X105Y79_IOB_X1Y79_O;
  wire [0:0] RIOB33_X105Y79_IOB_X1Y80_O;
  wire [0:0] RIOB33_X105Y81_IOB_X1Y81_O;
  wire [0:0] RIOB33_X105Y81_IOB_X1Y82_O;
  wire [0:0] RIOB33_X105Y83_IOB_X1Y83_O;
  wire [0:0] RIOB33_X105Y83_IOB_X1Y84_O;
  wire [0:0] RIOB33_X105Y85_IOB_X1Y85_O;
  wire [0:0] RIOB33_X105Y85_IOB_X1Y86_O;
  wire [0:0] RIOB33_X105Y87_IOB_X1Y87_O;
  wire [0:0] RIOB33_X105Y87_IOB_X1Y88_O;
  wire [0:0] RIOB33_X105Y89_IOB_X1Y89_O;
  wire [0:0] RIOB33_X105Y89_IOB_X1Y90_O;
  wire [0:0] RIOB33_X105Y91_IOB_X1Y91_O;
  wire [0:0] RIOI3_SING_X105Y100_OLOGIC_X1Y100_D1;
  wire [0:0] RIOI3_SING_X105Y100_OLOGIC_X1Y100_OQ;
  wire [0:0] RIOI3_SING_X105Y100_OLOGIC_X1Y100_T1;
  wire [0:0] RIOI3_SING_X105Y100_OLOGIC_X1Y100_TQ;
  wire [0:0] RIOI3_SING_X105Y149_OLOGIC_X1Y149_D1;
  wire [0:0] RIOI3_SING_X105Y149_OLOGIC_X1Y149_OQ;
  wire [0:0] RIOI3_SING_X105Y149_OLOGIC_X1Y149_T1;
  wire [0:0] RIOI3_SING_X105Y149_OLOGIC_X1Y149_TQ;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ;
  wire [0:0] RIOI3_SING_X105Y50_ILOGIC_X1Y50_D;
  wire [0:0] RIOI3_SING_X105Y50_ILOGIC_X1Y50_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_ILOGIC_X1Y57_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_ILOGIC_X1Y57_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_ILOGIC_X1Y58_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_ILOGIC_X1Y58_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_TQ;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y101_D1;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y101_OQ;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y101_T1;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y101_TQ;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y102_D1;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y102_OQ;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y102_T1;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y102_TQ;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y103_D1;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y103_OQ;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y103_T1;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y103_TQ;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y104_D1;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y104_OQ;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y104_T1;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y104_TQ;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y105_D1;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y105_OQ;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y105_T1;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y105_TQ;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y106_D1;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y106_OQ;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y106_T1;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y106_TQ;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y109_D1;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y109_OQ;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y109_T1;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y109_TQ;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y110_D1;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y110_OQ;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y110_T1;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y110_TQ;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y111_D1;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y111_OQ;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y111_T1;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y111_TQ;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y112_D1;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y112_OQ;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y112_T1;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y112_TQ;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y115_D1;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y115_OQ;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y115_T1;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y115_TQ;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y116_D1;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y116_OQ;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y116_T1;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y116_TQ;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y117_D1;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y117_OQ;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y117_T1;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y117_TQ;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y118_D1;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y118_OQ;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y118_T1;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y118_TQ;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y121_D1;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y121_OQ;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y121_T1;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y121_TQ;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y122_D1;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y122_OQ;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y122_T1;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y122_TQ;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y123_D1;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y123_OQ;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y123_T1;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y123_TQ;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y124_D1;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y124_OQ;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y124_T1;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y124_TQ;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y125_D1;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y125_OQ;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y125_T1;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y125_TQ;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y126_D1;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y126_OQ;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y126_T1;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y126_TQ;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_D1;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_OQ;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_T1;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_TQ;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y128_D1;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y128_OQ;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y128_T1;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y128_TQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_D1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_OQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_T1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_TQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_D1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_OQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_T1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_TQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_D1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_OQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_T1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_TQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_D1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_OQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_T1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_TQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_D1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_OQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_T1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_TQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_D1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_OQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_T1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_TQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_D1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_OQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_T1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_TQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_D1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_OQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_T1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_TQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_D1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_OQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_T1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_TQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_D1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_OQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_T1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_TQ;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_D1;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_OQ;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_T1;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_TQ;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y146_D1;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y146_OQ;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y146_T1;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y146_TQ;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y147_D1;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y147_OQ;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y147_T1;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y147_TQ;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y148_D1;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y148_OQ;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y148_T1;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y148_TQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_TQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_TQ;
  wire [0:0] RIOI3_X105Y51_ILOGIC_X1Y51_D;
  wire [0:0] RIOI3_X105Y51_ILOGIC_X1Y51_O;
  wire [0:0] RIOI3_X105Y51_ILOGIC_X1Y52_D;
  wire [0:0] RIOI3_X105Y51_ILOGIC_X1Y52_O;
  wire [0:0] RIOI3_X105Y53_ILOGIC_X1Y53_D;
  wire [0:0] RIOI3_X105Y53_ILOGIC_X1Y53_O;
  wire [0:0] RIOI3_X105Y53_ILOGIC_X1Y54_D;
  wire [0:0] RIOI3_X105Y53_ILOGIC_X1Y54_O;
  wire [0:0] RIOI3_X105Y55_ILOGIC_X1Y55_D;
  wire [0:0] RIOI3_X105Y55_ILOGIC_X1Y55_O;
  wire [0:0] RIOI3_X105Y55_ILOGIC_X1Y56_D;
  wire [0:0] RIOI3_X105Y55_ILOGIC_X1Y56_O;
  wire [0:0] RIOI3_X105Y59_ILOGIC_X1Y59_D;
  wire [0:0] RIOI3_X105Y59_ILOGIC_X1Y59_O;
  wire [0:0] RIOI3_X105Y59_ILOGIC_X1Y60_D;
  wire [0:0] RIOI3_X105Y59_ILOGIC_X1Y60_O;
  wire [0:0] RIOI3_X105Y61_ILOGIC_X1Y62_D;
  wire [0:0] RIOI3_X105Y61_ILOGIC_X1Y62_O;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y65_D1;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y65_OQ;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y65_T1;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y65_TQ;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y66_D1;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y66_OQ;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y66_T1;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y66_TQ;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y67_D1;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y67_OQ;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y67_T1;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y67_TQ;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y68_D1;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y68_OQ;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y68_T1;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y68_TQ;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y71_D1;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y71_OQ;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y71_T1;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y71_TQ;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y72_D1;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y72_OQ;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y72_T1;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y72_TQ;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y73_D1;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y73_OQ;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y73_T1;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y73_TQ;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y74_D1;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y74_OQ;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y74_T1;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y74_TQ;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y75_D1;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y75_OQ;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y75_T1;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y75_TQ;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y76_D1;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y76_OQ;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y76_T1;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y76_TQ;
  wire [0:0] RIOI3_X105Y77_ILOGIC_X1Y78_D;
  wire [0:0] RIOI3_X105Y77_ILOGIC_X1Y78_O;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y77_D1;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y77_OQ;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y77_T1;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y77_TQ;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y79_D1;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y79_OQ;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y79_T1;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y79_TQ;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y80_D1;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y80_OQ;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y80_T1;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y80_TQ;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y83_D1;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y83_OQ;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y83_T1;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y83_TQ;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y84_D1;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y84_OQ;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y84_T1;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y84_TQ;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y85_D1;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y85_OQ;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y85_T1;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y85_TQ;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y86_D1;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y86_OQ;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y86_T1;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y86_TQ;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y89_D1;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y89_OQ;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y89_T1;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y89_TQ;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y90_D1;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y90_OQ;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y90_T1;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y90_TQ;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y91_D1;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y91_OQ;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y91_T1;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y91_TQ;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X0Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X0Y131_DO5),
.O6(CLBLL_L_X2Y131_SLICE_X0Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X0Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X0Y131_CO5),
.O6(CLBLL_L_X2Y131_SLICE_X0Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X0Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X0Y131_BO5),
.O6(CLBLL_L_X2Y131_SLICE_X0Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffff0000ffff)
  ) CLBLL_L_X2Y131_SLICE_X0Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_R_X73Y123_SLICE_X110Y123_AQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X0Y131_AO5),
.O6(CLBLL_L_X2Y131_SLICE_X0Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X1Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X1Y131_DO5),
.O6(CLBLL_L_X2Y131_SLICE_X1Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X1Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X1Y131_CO5),
.O6(CLBLL_L_X2Y131_SLICE_X1Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X1Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X1Y131_BO5),
.O6(CLBLL_L_X2Y131_SLICE_X1Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X1Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X1Y131_AO5),
.O6(CLBLL_L_X2Y131_SLICE_X1Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y123_SLICE_X50Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y123_SLICE_X50Y123_DO5),
.O6(CLBLL_L_X34Y123_SLICE_X50Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y123_SLICE_X50Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y123_SLICE_X50Y123_CO5),
.O6(CLBLL_L_X34Y123_SLICE_X50Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y123_SLICE_X50Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y123_SLICE_X50Y123_BO5),
.O6(CLBLL_L_X34Y123_SLICE_X50Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffffffff)
  ) CLBLL_L_X34Y123_SLICE_X50Y123_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X53Y122_SLICE_X80Y122_AQ),
.O5(CLBLL_L_X34Y123_SLICE_X50Y123_AO5),
.O6(CLBLL_L_X34Y123_SLICE_X50Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y123_SLICE_X51Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y123_SLICE_X51Y123_DO5),
.O6(CLBLL_L_X34Y123_SLICE_X51Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y123_SLICE_X51Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y123_SLICE_X51Y123_CO5),
.O6(CLBLL_L_X34Y123_SLICE_X51Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y123_SLICE_X51Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y123_SLICE_X51Y123_BO5),
.O6(CLBLL_L_X34Y123_SLICE_X51Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y123_SLICE_X51Y123_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y123_SLICE_X51Y123_AO5),
.O6(CLBLL_L_X34Y123_SLICE_X51Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y126_SLICE_X50Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y126_SLICE_X50Y126_DO5),
.O6(CLBLL_L_X34Y126_SLICE_X50Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y126_SLICE_X50Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y126_SLICE_X50Y126_CO5),
.O6(CLBLL_L_X34Y126_SLICE_X50Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y126_SLICE_X50Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y126_SLICE_X50Y126_BO5),
.O6(CLBLL_L_X34Y126_SLICE_X50Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0f0f0f)
  ) CLBLL_L_X34Y126_SLICE_X50Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_R_X71Y124_SLICE_X106Y124_A5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y126_SLICE_X50Y126_AO5),
.O6(CLBLL_L_X34Y126_SLICE_X50Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y126_SLICE_X51Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y126_SLICE_X51Y126_DO5),
.O6(CLBLL_L_X34Y126_SLICE_X51Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y126_SLICE_X51Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y126_SLICE_X51Y126_CO5),
.O6(CLBLL_L_X34Y126_SLICE_X51Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y126_SLICE_X51Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y126_SLICE_X51Y126_BO5),
.O6(CLBLL_L_X34Y126_SLICE_X51Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y126_SLICE_X51Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y126_SLICE_X51Y126_AO5),
.O6(CLBLL_L_X34Y126_SLICE_X51Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y128_SLICE_X50Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y128_SLICE_X50Y128_DO5),
.O6(CLBLL_L_X34Y128_SLICE_X50Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y128_SLICE_X50Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y128_SLICE_X50Y128_CO5),
.O6(CLBLL_L_X34Y128_SLICE_X50Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y128_SLICE_X50Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y128_SLICE_X50Y128_BO5),
.O6(CLBLL_L_X34Y128_SLICE_X50Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00ff00ff)
  ) CLBLL_L_X34Y128_SLICE_X50Y128_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_R_X73Y125_SLICE_X111Y125_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y128_SLICE_X50Y128_AO5),
.O6(CLBLL_L_X34Y128_SLICE_X50Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y128_SLICE_X51Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y128_SLICE_X51Y128_DO5),
.O6(CLBLL_L_X34Y128_SLICE_X51Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y128_SLICE_X51Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y128_SLICE_X51Y128_CO5),
.O6(CLBLL_L_X34Y128_SLICE_X51Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y128_SLICE_X51Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y128_SLICE_X51Y128_BO5),
.O6(CLBLL_L_X34Y128_SLICE_X51Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y128_SLICE_X51Y128_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y128_SLICE_X51Y128_AO5),
.O6(CLBLL_L_X34Y128_SLICE_X51Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y98_SLICE_X106Y98_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y98_SLICE_X106Y98_AO5),
.Q(CLBLL_R_X71Y98_SLICE_X106Y98_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y98_SLICE_X106Y98_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y98_SLICE_X106Y98_AO6),
.Q(CLBLL_R_X71Y98_SLICE_X106Y98_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y98_SLICE_X106Y98_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y98_SLICE_X106Y98_DO5),
.O6(CLBLL_R_X71Y98_SLICE_X106Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y98_SLICE_X106Y98_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y98_SLICE_X106Y98_CO5),
.O6(CLBLL_R_X71Y98_SLICE_X106Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y98_SLICE_X106Y98_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y98_SLICE_X106Y98_BO5),
.O6(CLBLL_R_X71Y98_SLICE_X106Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee44445f0af5a0)
  ) CLBLL_R_X71Y98_SLICE_X106Y98_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X72Y98_SLICE_X108Y98_AQ),
.I2(CLBLL_R_X71Y100_SLICE_X106Y100_AO5),
.I3(CLBLM_L_X70Y98_SLICE_X104Y98_AQ),
.I4(CLBLL_R_X71Y98_SLICE_X106Y98_A5Q),
.I5(1'b1),
.O5(CLBLL_R_X71Y98_SLICE_X106Y98_AO5),
.O6(CLBLL_R_X71Y98_SLICE_X106Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y98_SLICE_X107Y98_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y98_SLICE_X107Y98_DO5),
.O6(CLBLL_R_X71Y98_SLICE_X107Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y98_SLICE_X107Y98_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y98_SLICE_X107Y98_CO5),
.O6(CLBLL_R_X71Y98_SLICE_X107Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y98_SLICE_X107Y98_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y98_SLICE_X107Y98_BO5),
.O6(CLBLL_R_X71Y98_SLICE_X107Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y98_SLICE_X107Y98_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y98_SLICE_X107Y98_AO5),
.O6(CLBLL_R_X71Y98_SLICE_X107Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y100_SLICE_X106Y100_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y100_SLICE_X106Y100_BO6),
.Q(CLBLL_R_X71Y100_SLICE_X106Y100_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000550030001100)
  ) CLBLL_R_X71Y100_SLICE_X106Y100_DLUT (
.I0(CLBLM_L_X70Y100_SLICE_X105Y100_CQ),
.I1(CLBLM_L_X70Y100_SLICE_X104Y100_A5Q),
.I2(CLBLL_R_X71Y100_SLICE_X106Y100_BQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLL_R_X77Y108_SLICE_X118Y108_AQ),
.I5(CLBLM_L_X60Y97_SLICE_X90Y97_BQ),
.O5(CLBLL_R_X71Y100_SLICE_X106Y100_DO5),
.O6(CLBLL_R_X71Y100_SLICE_X106Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h808080800f000000)
  ) CLBLL_R_X71Y100_SLICE_X106Y100_CLUT (
.I0(CLBLM_L_X70Y100_SLICE_X105Y100_CQ),
.I1(CLBLL_R_X71Y101_SLICE_X106Y101_BQ),
.I2(CLBLM_L_X70Y100_SLICE_X105Y100_A5Q),
.I3(CLBLM_L_X60Y99_SLICE_X90Y99_AQ),
.I4(CLBLL_R_X71Y101_SLICE_X106Y101_CQ),
.I5(CLBLM_L_X70Y100_SLICE_X105Y100_AQ),
.O5(CLBLL_R_X71Y100_SLICE_X106Y100_CO5),
.O6(CLBLL_R_X71Y100_SLICE_X106Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7070000000f000f0)
  ) CLBLL_R_X71Y100_SLICE_X106Y100_BLUT (
.I0(CLBLL_R_X77Y108_SLICE_X118Y108_AQ),
.I1(CLBLL_R_X71Y100_SLICE_X106Y100_BQ),
.I2(CLBLL_R_X71Y100_SLICE_X106Y100_DO6),
.I3(CLBLM_L_X60Y97_SLICE_X90Y97_BQ),
.I4(CLBLM_L_X70Y100_SLICE_X105Y100_CQ),
.I5(CLBLM_L_X60Y99_SLICE_X90Y99_AQ),
.O5(CLBLL_R_X71Y100_SLICE_X106Y100_BO5),
.O6(CLBLL_R_X71Y100_SLICE_X106Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333cccc80008000)
  ) CLBLL_R_X71Y100_SLICE_X106Y100_ALUT (
.I0(CLBLL_R_X77Y108_SLICE_X118Y108_AQ),
.I1(CLBLL_R_X71Y100_SLICE_X106Y100_BQ),
.I2(CLBLM_L_X60Y99_SLICE_X90Y99_AQ),
.I3(CLBLM_L_X70Y100_SLICE_X105Y100_CQ),
.I4(CLBLL_R_X71Y98_SLICE_X106Y98_A5Q),
.I5(1'b1),
.O5(CLBLL_R_X71Y100_SLICE_X106Y100_AO5),
.O6(CLBLL_R_X71Y100_SLICE_X106Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y100_SLICE_X107Y100_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y100_SLICE_X107Y100_DO5),
.O6(CLBLL_R_X71Y100_SLICE_X107Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y100_SLICE_X107Y100_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y100_SLICE_X107Y100_CO5),
.O6(CLBLL_R_X71Y100_SLICE_X107Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y100_SLICE_X107Y100_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y100_SLICE_X107Y100_BO5),
.O6(CLBLL_R_X71Y100_SLICE_X107Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y100_SLICE_X107Y100_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y100_SLICE_X107Y100_AO5),
.O6(CLBLL_R_X71Y100_SLICE_X107Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y101_SLICE_X106Y101_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y101_SLICE_X106Y101_AO6),
.Q(CLBLL_R_X71Y101_SLICE_X106Y101_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y101_SLICE_X106Y101_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y101_SLICE_X106Y101_BO6),
.Q(CLBLL_R_X71Y101_SLICE_X106Y101_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y101_SLICE_X106Y101_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y101_SLICE_X106Y101_CO6),
.Q(CLBLL_R_X71Y101_SLICE_X106Y101_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4450005044000000)
  ) CLBLL_R_X71Y101_SLICE_X106Y101_DLUT (
.I0(CLBLM_L_X70Y100_SLICE_X105Y100_AQ),
.I1(CLBLL_R_X71Y102_SLICE_X106Y102_AQ),
.I2(CLBLL_R_X71Y103_SLICE_X106Y103_AQ),
.I3(CLBLM_L_X70Y100_SLICE_X105Y100_A5Q),
.I4(CLBLM_L_X70Y101_SLICE_X104Y101_AQ),
.I5(CLBLM_L_X70Y100_SLICE_X104Y100_A5Q),
.O5(CLBLL_R_X71Y101_SLICE_X106Y101_DO5),
.O6(CLBLL_R_X71Y101_SLICE_X106Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8d8d8d8fad850)
  ) CLBLL_R_X71Y101_SLICE_X106Y101_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X71Y101_SLICE_X106Y101_CQ),
.I2(CLBLL_R_X71Y101_SLICE_X106Y101_BQ),
.I3(CLBLM_L_X70Y103_SLICE_X105Y103_DO5),
.I4(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I5(CLBLL_R_X71Y103_SLICE_X106Y103_BO6),
.O5(CLBLL_R_X71Y101_SLICE_X106Y101_CO5),
.O6(CLBLL_R_X71Y101_SLICE_X106Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00d8ffd800)
  ) CLBLL_R_X71Y101_SLICE_X106Y101_BLUT (
.I0(CLBLM_L_X70Y103_SLICE_X105Y103_DO6),
.I1(CLBLL_R_X71Y101_SLICE_X106Y101_BQ),
.I2(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLL_R_X71Y102_SLICE_X106Y102_BQ),
.I5(CLBLL_R_X71Y103_SLICE_X106Y103_BO6),
.O5(CLBLL_R_X71Y101_SLICE_X106Y101_BO5),
.O6(CLBLL_R_X71Y101_SLICE_X106Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ccccf0aacccc)
  ) CLBLL_R_X71Y101_SLICE_X106Y101_ALUT (
.I0(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I1(CLBLM_L_X70Y101_SLICE_X104Y101_CQ),
.I2(CLBLL_R_X71Y101_SLICE_X106Y101_AQ),
.I3(CLBLM_L_X70Y103_SLICE_X104Y103_DO5),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X70Y103_SLICE_X105Y103_CO5),
.O5(CLBLL_R_X71Y101_SLICE_X106Y101_AO5),
.O6(CLBLL_R_X71Y101_SLICE_X106Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y101_SLICE_X107Y101_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y101_SLICE_X107Y101_AO6),
.Q(CLBLL_R_X71Y101_SLICE_X107Y101_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y101_SLICE_X107Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y101_SLICE_X107Y101_DO5),
.O6(CLBLL_R_X71Y101_SLICE_X107Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y101_SLICE_X107Y101_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y101_SLICE_X107Y101_CO5),
.O6(CLBLL_R_X71Y101_SLICE_X107Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y101_SLICE_X107Y101_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y101_SLICE_X107Y101_BO5),
.O6(CLBLL_R_X71Y101_SLICE_X107Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1e0f1e0ffff0000)
  ) CLBLL_R_X71Y101_SLICE_X107Y101_ALUT (
.I0(CLBLM_L_X70Y103_SLICE_X105Y103_DO6),
.I1(CLBLM_L_X70Y103_SLICE_X105Y103_CO5),
.I2(CLBLL_R_X71Y101_SLICE_X107Y101_AQ),
.I3(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I4(CLBLL_R_X71Y101_SLICE_X106Y101_AQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLL_R_X71Y101_SLICE_X107Y101_AO5),
.O6(CLBLL_R_X71Y101_SLICE_X107Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y102_SLICE_X106Y102_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y102_SLICE_X106Y102_AO6),
.Q(CLBLL_R_X71Y102_SLICE_X106Y102_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y102_SLICE_X106Y102_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y102_SLICE_X106Y102_BO6),
.Q(CLBLL_R_X71Y102_SLICE_X106Y102_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y102_SLICE_X106Y102_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y102_SLICE_X106Y102_CO6),
.Q(CLBLL_R_X71Y102_SLICE_X106Y102_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h13ff5fff335fff5f)
  ) CLBLL_R_X71Y102_SLICE_X106Y102_DLUT (
.I0(CLBLL_R_X71Y102_SLICE_X106Y102_BQ),
.I1(CLBLL_R_X71Y102_SLICE_X106Y102_CQ),
.I2(CLBLL_R_X77Y108_SLICE_X118Y108_AQ),
.I3(CLBLL_R_X71Y98_SLICE_X106Y98_A5Q),
.I4(CLBLM_L_X70Y101_SLICE_X105Y101_AQ),
.I5(CLBLL_R_X71Y100_SLICE_X106Y100_BQ),
.O5(CLBLL_R_X71Y102_SLICE_X106Y102_DO5),
.O6(CLBLL_R_X71Y102_SLICE_X106Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccf0ccf0aaf0)
  ) CLBLL_R_X71Y102_SLICE_X106Y102_CLUT (
.I0(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I1(CLBLL_R_X71Y102_SLICE_X106Y102_CQ),
.I2(CLBLL_R_X71Y102_SLICE_X106Y102_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X70Y103_SLICE_X105Y103_DO6),
.I5(CLBLL_R_X71Y103_SLICE_X106Y103_BO5),
.O5(CLBLL_R_X71Y102_SLICE_X106Y102_CO5),
.O6(CLBLL_R_X71Y102_SLICE_X106Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddfddd5888a8880)
  ) CLBLL_R_X71Y102_SLICE_X106Y102_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X71Y102_SLICE_X106Y102_BQ),
.I2(CLBLL_R_X71Y103_SLICE_X106Y103_BO6),
.I3(CLBLM_L_X70Y103_SLICE_X104Y103_DO5),
.I4(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I5(CLBLM_L_X70Y102_SLICE_X105Y102_AQ),
.O5(CLBLL_R_X71Y102_SLICE_X106Y102_BO5),
.O6(CLBLL_R_X71Y102_SLICE_X106Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1ffe0fff100e000)
  ) CLBLL_R_X71Y102_SLICE_X106Y102_ALUT (
.I0(CLBLL_R_X71Y103_SLICE_X106Y103_BO5),
.I1(CLBLM_L_X70Y103_SLICE_X104Y103_DO5),
.I2(CLBLL_R_X71Y102_SLICE_X106Y102_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I5(CLBLL_R_X71Y103_SLICE_X106Y103_AQ),
.O5(CLBLL_R_X71Y102_SLICE_X106Y102_AO5),
.O6(CLBLL_R_X71Y102_SLICE_X106Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y102_SLICE_X107Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y102_SLICE_X107Y102_DO5),
.O6(CLBLL_R_X71Y102_SLICE_X107Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y102_SLICE_X107Y102_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y102_SLICE_X107Y102_CO5),
.O6(CLBLL_R_X71Y102_SLICE_X107Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y102_SLICE_X107Y102_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y102_SLICE_X107Y102_BO5),
.O6(CLBLL_R_X71Y102_SLICE_X107Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y102_SLICE_X107Y102_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y102_SLICE_X107Y102_AO5),
.O6(CLBLL_R_X71Y102_SLICE_X107Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y103_SLICE_X106Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y103_SLICE_X106Y103_AO6),
.Q(CLBLL_R_X71Y103_SLICE_X106Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y103_SLICE_X106Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y103_SLICE_X106Y103_DO5),
.O6(CLBLL_R_X71Y103_SLICE_X106Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y103_SLICE_X106Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y103_SLICE_X106Y103_CO5),
.O6(CLBLL_R_X71Y103_SLICE_X106Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafafaffafafafa)
  ) CLBLL_R_X71Y103_SLICE_X106Y103_BLUT (
.I0(CLBLM_L_X70Y104_SLICE_X104Y104_A5Q),
.I1(1'b1),
.I2(CLBLM_L_X70Y103_SLICE_X104Y103_B5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y103_SLICE_X106Y103_BO5),
.O6(CLBLL_R_X71Y103_SLICE_X106Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f1e0aaaaaaaa)
  ) CLBLL_R_X71Y103_SLICE_X106Y103_ALUT (
.I0(CLBLM_L_X70Y104_SLICE_X104Y104_A5Q),
.I1(CLBLM_L_X70Y103_SLICE_X104Y103_DO6),
.I2(CLBLL_R_X71Y103_SLICE_X106Y103_AQ),
.I3(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I4(CLBLM_L_X70Y103_SLICE_X104Y103_B5Q),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLL_R_X71Y103_SLICE_X106Y103_AO5),
.O6(CLBLL_R_X71Y103_SLICE_X106Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y103_SLICE_X107Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y103_SLICE_X107Y103_DO5),
.O6(CLBLL_R_X71Y103_SLICE_X107Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y103_SLICE_X107Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y103_SLICE_X107Y103_CO5),
.O6(CLBLL_R_X71Y103_SLICE_X107Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y103_SLICE_X107Y103_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y103_SLICE_X107Y103_BO5),
.O6(CLBLL_R_X71Y103_SLICE_X107Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y103_SLICE_X107Y103_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y103_SLICE_X107Y103_AO5),
.O6(CLBLL_R_X71Y103_SLICE_X107Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y107_SLICE_X106Y107_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y107_SLICE_X106Y107_CO5),
.Q(CLBLL_R_X71Y107_SLICE_X106Y107_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y107_SLICE_X106Y107_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y107_SLICE_X106Y107_AO6),
.Q(CLBLL_R_X71Y107_SLICE_X106Y107_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y107_SLICE_X106Y107_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y107_SLICE_X106Y107_CO6),
.Q(CLBLL_R_X71Y107_SLICE_X106Y107_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdeccedfcccccccc)
  ) CLBLL_R_X71Y107_SLICE_X106Y107_DLUT (
.I0(CLBLL_R_X71Y107_SLICE_X106Y107_C5Q),
.I1(CLBLM_L_X70Y107_SLICE_X105Y107_BQ),
.I2(CLBLL_R_X71Y107_SLICE_X107Y107_C5Q),
.I3(CLBLL_R_X71Y107_SLICE_X107Y107_CQ),
.I4(CLBLL_R_X71Y107_SLICE_X106Y107_CQ),
.I5(CLBLM_L_X70Y106_SLICE_X105Y106_CO6),
.O5(CLBLL_R_X71Y107_SLICE_X106Y107_DO5),
.O6(CLBLL_R_X71Y107_SLICE_X106Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5afaaa0a5cac5cac)
  ) CLBLL_R_X71Y107_SLICE_X106Y107_CLUT (
.I0(CLBLL_R_X71Y107_SLICE_X106Y107_C5Q),
.I1(CLBLL_R_X71Y107_SLICE_X107Y107_C5Q),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X70Y106_SLICE_X105Y106_CO6),
.I4(CLBLL_R_X71Y107_SLICE_X106Y107_CQ),
.I5(1'b1),
.O5(CLBLL_R_X71Y107_SLICE_X106Y107_CO5),
.O6(CLBLL_R_X71Y107_SLICE_X106Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h800000007f7fffff)
  ) CLBLL_R_X71Y107_SLICE_X106Y107_BLUT (
.I0(CLBLL_R_X73Y108_SLICE_X110Y108_A5Q),
.I1(CLBLM_L_X62Y92_SLICE_X92Y92_AQ),
.I2(CLBLL_R_X71Y107_SLICE_X106Y107_CQ),
.I3(CLBLM_L_X70Y106_SLICE_X105Y106_CO6),
.I4(CLBLL_R_X71Y107_SLICE_X106Y107_C5Q),
.I5(1'b1),
.O5(CLBLL_R_X71Y107_SLICE_X106Y107_BO5),
.O6(CLBLL_R_X71Y107_SLICE_X106Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc3cffffcc3c0000)
  ) CLBLL_R_X71Y107_SLICE_X106Y107_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X72Y106_SLICE_X108Y106_CO6),
.I2(CLBLL_R_X71Y107_SLICE_X106Y107_AQ),
.I3(CLBLL_R_X71Y107_SLICE_X106Y107_BO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X71Y108_SLICE_X106Y108_AQ),
.O5(CLBLL_R_X71Y107_SLICE_X106Y107_AO5),
.O6(CLBLL_R_X71Y107_SLICE_X106Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y107_SLICE_X107Y107_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y107_SLICE_X107Y107_CO5),
.Q(CLBLL_R_X71Y107_SLICE_X107Y107_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y107_SLICE_X107Y107_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y107_SLICE_X107Y107_AO6),
.Q(CLBLL_R_X71Y107_SLICE_X107Y107_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y107_SLICE_X107Y107_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y107_SLICE_X107Y107_BO6),
.Q(CLBLL_R_X71Y107_SLICE_X107Y107_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y107_SLICE_X107Y107_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y107_SLICE_X107Y107_CO6),
.Q(CLBLL_R_X71Y107_SLICE_X107Y107_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0cc0000a0000000)
  ) CLBLL_R_X71Y107_SLICE_X107Y107_DLUT (
.I0(CLBLM_L_X72Y107_SLICE_X108Y107_BQ),
.I1(CLBLM_L_X72Y107_SLICE_X109Y107_BQ),
.I2(CLBLM_L_X72Y108_SLICE_X108Y108_CQ),
.I3(CLBLL_R_X71Y107_SLICE_X106Y107_CQ),
.I4(CLBLL_R_X71Y107_SLICE_X106Y107_C5Q),
.I5(CLBLL_R_X71Y107_SLICE_X107Y107_AQ),
.O5(CLBLL_R_X71Y107_SLICE_X107Y107_DO5),
.O6(CLBLL_R_X71Y107_SLICE_X107Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0555f0f00ccccccc)
  ) CLBLL_R_X71Y107_SLICE_X107Y107_CLUT (
.I0(CLBLL_R_X71Y107_SLICE_X107Y107_C5Q),
.I1(CLBLL_R_X71Y107_SLICE_X107Y107_CQ),
.I2(CLBLL_R_X73Y108_SLICE_X110Y108_A5Q),
.I3(CLBLM_L_X72Y107_SLICE_X109Y107_DO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLL_R_X71Y107_SLICE_X107Y107_CO5),
.O6(CLBLL_R_X71Y107_SLICE_X107Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cfc0dfd08f80)
  ) CLBLL_R_X71Y107_SLICE_X107Y107_BLUT (
.I0(CLBLL_R_X71Y109_SLICE_X106Y109_CO6),
.I1(CLBLL_R_X71Y107_SLICE_X107Y107_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLL_R_X71Y107_SLICE_X107Y107_AQ),
.I4(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I5(CLBLM_L_X72Y108_SLICE_X109Y108_BO5),
.O5(CLBLL_R_X71Y107_SLICE_X107Y107_BO5),
.O6(CLBLL_R_X71Y107_SLICE_X107Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0f7a2d580)
  ) CLBLL_R_X71Y107_SLICE_X107Y107_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X72Y108_SLICE_X109Y108_BO6),
.I2(CLBLL_R_X71Y107_SLICE_X107Y107_AQ),
.I3(CLBLM_L_X72Y108_SLICE_X108Y108_AQ),
.I4(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I5(CLBLL_R_X71Y109_SLICE_X106Y109_CO6),
.O5(CLBLL_R_X71Y107_SLICE_X107Y107_AO5),
.O6(CLBLL_R_X71Y107_SLICE_X107Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y108_SLICE_X106Y108_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y108_SLICE_X106Y108_DO5),
.Q(CLBLL_R_X71Y108_SLICE_X106Y108_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y108_SLICE_X106Y108_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y108_SLICE_X106Y108_AO6),
.Q(CLBLL_R_X71Y108_SLICE_X106Y108_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y108_SLICE_X106Y108_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y108_SLICE_X106Y108_BO6),
.Q(CLBLL_R_X71Y108_SLICE_X106Y108_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y108_SLICE_X106Y108_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y108_SLICE_X106Y108_CO6),
.Q(CLBLL_R_X71Y108_SLICE_X106Y108_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y108_SLICE_X106Y108_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y108_SLICE_X106Y108_DO6),
.Q(CLBLL_R_X71Y108_SLICE_X106Y108_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcce4cce4d2fad250)
  ) CLBLL_R_X71Y108_SLICE_X106Y108_DLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X71Y108_SLICE_X106Y108_CQ),
.I2(CLBLL_R_X71Y108_SLICE_X106Y108_DQ),
.I3(CLBLL_R_X71Y107_SLICE_X106Y107_BO6),
.I4(CLBLL_R_X71Y108_SLICE_X106Y108_D5Q),
.I5(1'b1),
.O5(CLBLL_R_X71Y108_SLICE_X106Y108_DO5),
.O6(CLBLL_R_X71Y108_SLICE_X106Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7d28dd88dd88dd88)
  ) CLBLL_R_X71Y108_SLICE_X106Y108_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X71Y108_SLICE_X106Y108_CQ),
.I2(CLBLM_L_X72Y108_SLICE_X109Y108_A5Q),
.I3(CLBLL_R_X71Y108_SLICE_X106Y108_BQ),
.I4(CLBLL_R_X71Y109_SLICE_X106Y109_B5Q),
.I5(CLBLL_R_X71Y109_SLICE_X106Y109_BQ),
.O5(CLBLL_R_X71Y108_SLICE_X106Y108_CO5),
.O6(CLBLL_R_X71Y108_SLICE_X106Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fccfffff0cc0000)
  ) CLBLL_R_X71Y108_SLICE_X106Y108_BLUT (
.I0(1'b1),
.I1(CLBLL_R_X71Y108_SLICE_X106Y108_BQ),
.I2(CLBLL_R_X71Y108_SLICE_X106Y108_AQ),
.I3(CLBLL_R_X71Y107_SLICE_X106Y107_BO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X71Y107_SLICE_X106Y107_AQ),
.O5(CLBLL_R_X71Y108_SLICE_X106Y108_BO5),
.O6(CLBLL_R_X71Y108_SLICE_X106Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8f070f0ffff0000)
  ) CLBLL_R_X71Y108_SLICE_X106Y108_ALUT (
.I0(CLBLL_R_X71Y109_SLICE_X106Y109_B5Q),
.I1(CLBLL_R_X71Y109_SLICE_X106Y109_BQ),
.I2(CLBLL_R_X71Y108_SLICE_X106Y108_AQ),
.I3(CLBLM_L_X72Y108_SLICE_X109Y108_A5Q),
.I4(CLBLL_R_X71Y108_SLICE_X107Y108_AQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLL_R_X71Y108_SLICE_X106Y108_AO5),
.O6(CLBLL_R_X71Y108_SLICE_X106Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y108_SLICE_X107Y108_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y109_SLICE_X109Y109_DQ),
.Q(CLBLL_R_X71Y108_SLICE_X107Y108_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y108_SLICE_X107Y108_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y108_SLICE_X107Y108_AO6),
.Q(CLBLL_R_X71Y108_SLICE_X107Y108_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y108_SLICE_X107Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y108_SLICE_X107Y108_DO5),
.O6(CLBLL_R_X71Y108_SLICE_X107Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y108_SLICE_X107Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y108_SLICE_X107Y108_CO5),
.O6(CLBLL_R_X71Y108_SLICE_X107Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y108_SLICE_X107Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y108_SLICE_X107Y108_BO5),
.O6(CLBLL_R_X71Y108_SLICE_X107Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h70f000008f0f0000)
  ) CLBLL_R_X71Y108_SLICE_X107Y108_ALUT (
.I0(CLBLL_R_X71Y109_SLICE_X106Y109_B5Q),
.I1(CLBLM_L_X72Y108_SLICE_X109Y108_A5Q),
.I2(CLBLL_R_X71Y108_SLICE_X107Y108_AQ),
.I3(CLBLL_R_X71Y109_SLICE_X106Y109_BQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X79Y99_SLICE_X122Y99_AO6),
.O5(CLBLL_R_X71Y108_SLICE_X107Y108_AO5),
.O6(CLBLL_R_X71Y108_SLICE_X107Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y109_SLICE_X106Y109_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y109_SLICE_X106Y109_BO5),
.Q(CLBLL_R_X71Y109_SLICE_X106Y109_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y109_SLICE_X106Y109_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y109_SLICE_X106Y109_AO6),
.Q(CLBLL_R_X71Y109_SLICE_X106Y109_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y109_SLICE_X106Y109_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y109_SLICE_X106Y109_BO6),
.Q(CLBLL_R_X71Y109_SLICE_X106Y109_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y109_SLICE_X106Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y109_SLICE_X106Y109_DO5),
.O6(CLBLL_R_X71Y109_SLICE_X106Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaaaaaa000000)
  ) CLBLL_R_X71Y109_SLICE_X106Y109_CLUT (
.I0(CLBLL_R_X71Y109_SLICE_X106Y109_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X72Y108_SLICE_X109Y108_A5Q),
.I4(CLBLL_R_X71Y109_SLICE_X106Y109_B5Q),
.I5(1'b1),
.O5(CLBLL_R_X71Y109_SLICE_X106Y109_CO5),
.O6(CLBLL_R_X71Y109_SLICE_X106Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff0ff005fafa0a0)
  ) CLBLL_R_X71Y109_SLICE_X106Y109_BLUT (
.I0(CLBLL_R_X71Y109_SLICE_X106Y109_B5Q),
.I1(1'b1),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X72Y108_SLICE_X109Y108_A5Q),
.I4(CLBLL_R_X71Y109_SLICE_X106Y109_BQ),
.I5(1'b1),
.O5(CLBLL_R_X71Y109_SLICE_X106Y109_BO5),
.O6(CLBLL_R_X71Y109_SLICE_X106Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0cc33ccf0cc)
  ) CLBLL_R_X71Y109_SLICE_X106Y109_ALUT (
.I0(1'b1),
.I1(CLBLL_R_X71Y110_SLICE_X106Y110_BQ),
.I2(CLBLL_R_X71Y109_SLICE_X106Y109_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLL_R_X71Y109_SLICE_X106Y109_CO5),
.I5(CLBLL_R_X71Y110_SLICE_X106Y110_AQ),
.O5(CLBLL_R_X71Y109_SLICE_X106Y109_AO5),
.O6(CLBLL_R_X71Y109_SLICE_X106Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y109_SLICE_X107Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y109_SLICE_X107Y109_DO5),
.O6(CLBLL_R_X71Y109_SLICE_X107Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y109_SLICE_X107Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y109_SLICE_X107Y109_CO5),
.O6(CLBLL_R_X71Y109_SLICE_X107Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y109_SLICE_X107Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y109_SLICE_X107Y109_BO5),
.O6(CLBLL_R_X71Y109_SLICE_X107Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y109_SLICE_X107Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y109_SLICE_X107Y109_AO5),
.O6(CLBLL_R_X71Y109_SLICE_X107Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y110_SLICE_X106Y110_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y110_SLICE_X106Y110_AO5),
.Q(CLBLL_R_X71Y110_SLICE_X106Y110_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y110_SLICE_X106Y110_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y110_SLICE_X106Y110_AO6),
.Q(CLBLL_R_X71Y110_SLICE_X106Y110_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y110_SLICE_X106Y110_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y110_SLICE_X106Y110_BO6),
.Q(CLBLL_R_X71Y110_SLICE_X106Y110_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y110_SLICE_X106Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y110_SLICE_X106Y110_DO5),
.O6(CLBLL_R_X71Y110_SLICE_X106Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y110_SLICE_X106Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y110_SLICE_X106Y110_CO5),
.O6(CLBLL_R_X71Y110_SLICE_X106Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he4ccf0f0ccccf0f0)
  ) CLBLL_R_X71Y110_SLICE_X106Y110_BLUT (
.I0(CLBLL_R_X71Y109_SLICE_X106Y109_B5Q),
.I1(CLBLL_R_X71Y110_SLICE_X106Y110_BQ),
.I2(CLBLL_R_X71Y110_SLICE_X106Y110_AQ),
.I3(CLBLM_L_X72Y108_SLICE_X109Y108_A5Q),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X71Y109_SLICE_X106Y109_BQ),
.O5(CLBLL_R_X71Y110_SLICE_X106Y110_BO5),
.O6(CLBLL_R_X71Y110_SLICE_X106Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff0aaaa33330000)
  ) CLBLL_R_X71Y110_SLICE_X106Y110_ALUT (
.I0(CLBLL_R_X71Y108_SLICE_X106Y108_D5Q),
.I1(CLBLL_R_X71Y114_SLICE_X106Y114_AQ),
.I2(CLBLL_R_X71Y110_SLICE_X106Y110_AQ),
.I3(CLBLL_R_X71Y107_SLICE_X106Y107_BO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLL_R_X71Y110_SLICE_X106Y110_AO5),
.O6(CLBLL_R_X71Y110_SLICE_X106Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y110_SLICE_X107Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y110_SLICE_X107Y110_DO5),
.O6(CLBLL_R_X71Y110_SLICE_X107Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y110_SLICE_X107Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y110_SLICE_X107Y110_CO5),
.O6(CLBLL_R_X71Y110_SLICE_X107Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y110_SLICE_X107Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y110_SLICE_X107Y110_BO5),
.O6(CLBLL_R_X71Y110_SLICE_X107Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y110_SLICE_X107Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y110_SLICE_X107Y110_AO5),
.O6(CLBLL_R_X71Y110_SLICE_X107Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y111_SLICE_X106Y111_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y111_SLICE_X106Y111_AO5),
.Q(CLBLL_R_X71Y111_SLICE_X106Y111_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y111_SLICE_X106Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y111_SLICE_X106Y111_AO6),
.Q(CLBLL_R_X71Y111_SLICE_X106Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y111_SLICE_X106Y111_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y111_SLICE_X106Y111_BO6),
.Q(CLBLL_R_X71Y111_SLICE_X106Y111_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y111_SLICE_X106Y111_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y111_SLICE_X106Y111_CO6),
.Q(CLBLL_R_X71Y111_SLICE_X106Y111_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb1b1001fb1b1001f)
  ) CLBLL_R_X71Y111_SLICE_X106Y111_DLUT (
.I0(CLBLL_R_X71Y111_SLICE_X107Y111_AQ),
.I1(CLBLL_R_X71Y111_SLICE_X107Y111_CO6),
.I2(CLBLM_L_X70Y112_SLICE_X104Y112_AQ),
.I3(CLBLM_L_X70Y111_SLICE_X104Y111_DO6),
.I4(CLBLM_L_X70Y112_SLICE_X104Y112_A5Q),
.I5(1'b1),
.O5(CLBLL_R_X71Y111_SLICE_X106Y111_DO5),
.O6(CLBLL_R_X71Y111_SLICE_X106Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h57085708dd88dd88)
  ) CLBLL_R_X71Y111_SLICE_X106Y111_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X71Y111_SLICE_X106Y111_CQ),
.I2(CLBLM_L_X70Y111_SLICE_X105Y111_BQ),
.I3(CLBLL_R_X71Y111_SLICE_X106Y111_BQ),
.I4(1'b1),
.I5(CLBLM_L_X70Y111_SLICE_X104Y111_BO5),
.O5(CLBLL_R_X71Y111_SLICE_X106Y111_CO5),
.O6(CLBLL_R_X71Y111_SLICE_X106Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ccaaaa33ccaaaa)
  ) CLBLL_R_X71Y111_SLICE_X106Y111_BLUT (
.I0(CLBLM_L_X70Y111_SLICE_X104Y111_AQ),
.I1(CLBLL_R_X71Y111_SLICE_X106Y111_BQ),
.I2(1'b1),
.I3(CLBLM_L_X70Y111_SLICE_X104Y111_BO5),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X70Y111_SLICE_X105Y111_BQ),
.O5(CLBLL_R_X71Y111_SLICE_X106Y111_BO5),
.O6(CLBLL_R_X71Y111_SLICE_X106Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h03030000aaaaff00)
  ) CLBLL_R_X71Y111_SLICE_X106Y111_ALUT (
.I0(CLBLL_R_X71Y111_SLICE_X106Y111_DO6),
.I1(CLBLM_L_X72Y108_SLICE_X109Y108_A5Q),
.I2(CLBLL_R_X71Y111_SLICE_X106Y111_AQ),
.I3(CLBLL_R_X71Y112_SLICE_X106Y112_AQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLL_R_X71Y111_SLICE_X106Y111_AO5),
.O6(CLBLL_R_X71Y111_SLICE_X106Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y111_SLICE_X107Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y111_SLICE_X107Y111_AO6),
.Q(CLBLL_R_X71Y111_SLICE_X107Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffcfffffffc)
  ) CLBLL_R_X71Y111_SLICE_X107Y111_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X70Y111_SLICE_X105Y111_BQ),
.I2(CLBLM_L_X70Y112_SLICE_X104Y112_A5Q),
.I3(CLBLL_R_X71Y111_SLICE_X106Y111_CQ),
.I4(CLBLM_L_X70Y112_SLICE_X104Y112_AQ),
.I5(1'b1),
.O5(CLBLL_R_X71Y111_SLICE_X107Y111_DO5),
.O6(CLBLL_R_X71Y111_SLICE_X107Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hef6def6df3b2f3b2)
  ) CLBLL_R_X71Y111_SLICE_X107Y111_CLUT (
.I0(CLBLL_R_X71Y111_SLICE_X106Y111_CQ),
.I1(CLBLM_L_X70Y111_SLICE_X105Y111_AQ),
.I2(CLBLM_L_X70Y111_SLICE_X104Y111_AQ),
.I3(CLBLM_L_X70Y111_SLICE_X105Y111_BQ),
.I4(1'b1),
.I5(CLBLL_R_X71Y111_SLICE_X106Y111_BQ),
.O5(CLBLL_R_X71Y111_SLICE_X107Y111_CO5),
.O6(CLBLL_R_X71Y111_SLICE_X107Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffef)
  ) CLBLL_R_X71Y111_SLICE_X107Y111_BLUT (
.I0(CLBLL_R_X71Y111_SLICE_X107Y111_DO6),
.I1(CLBLM_L_X70Y111_SLICE_X105Y111_AQ),
.I2(CLBLL_R_X71Y111_SLICE_X107Y111_AQ),
.I3(CLBLL_R_X71Y111_SLICE_X106Y111_BQ),
.I4(CLBLM_L_X72Y111_SLICE_X108Y111_AO6),
.I5(CLBLM_L_X70Y111_SLICE_X104Y111_AQ),
.O5(CLBLL_R_X71Y111_SLICE_X107Y111_BO5),
.O6(CLBLL_R_X71Y111_SLICE_X107Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa3faa00aac0aa)
  ) CLBLL_R_X71Y111_SLICE_X107Y111_ALUT (
.I0(CLBLM_L_X72Y111_SLICE_X109Y111_CQ),
.I1(CLBLM_L_X72Y111_SLICE_X109Y111_A5Q),
.I2(CLBLM_L_X72Y111_SLICE_X109Y111_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X70Y111_SLICE_X104Y111_BQ),
.I5(CLBLL_R_X71Y111_SLICE_X107Y111_AQ),
.O5(CLBLL_R_X71Y111_SLICE_X107Y111_AO5),
.O6(CLBLL_R_X71Y111_SLICE_X107Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y112_SLICE_X106Y112_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y112_SLICE_X106Y112_BO5),
.Q(CLBLL_R_X71Y112_SLICE_X106Y112_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y112_SLICE_X106Y112_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y112_SLICE_X106Y112_AO6),
.Q(CLBLL_R_X71Y112_SLICE_X106Y112_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y112_SLICE_X106Y112_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y112_SLICE_X106Y112_BO6),
.Q(CLBLL_R_X71Y112_SLICE_X106Y112_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y112_SLICE_X106Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y112_SLICE_X106Y112_DO5),
.O6(CLBLL_R_X71Y112_SLICE_X106Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y112_SLICE_X106Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y112_SLICE_X106Y112_CO5),
.O6(CLBLL_R_X71Y112_SLICE_X106Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha2aaaaaaececffff)
  ) CLBLL_R_X71Y112_SLICE_X106Y112_BLUT (
.I0(CLBLM_L_X70Y112_SLICE_X105Y112_A5Q),
.I1(CLBLL_R_X71Y112_SLICE_X106Y112_BQ),
.I2(CLBLL_R_X71Y112_SLICE_X106Y112_B5Q),
.I3(CLBLM_L_X72Y111_SLICE_X109Y111_CQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLL_R_X71Y112_SLICE_X106Y112_BO5),
.O6(CLBLL_R_X71Y112_SLICE_X106Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0b0f0f0f0f0f0)
  ) CLBLL_R_X71Y112_SLICE_X106Y112_ALUT (
.I0(CLBLL_R_X71Y111_SLICE_X107Y111_CO6),
.I1(CLBLM_L_X70Y112_SLICE_X104Y112_A5Q),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X70Y112_SLICE_X104Y112_AQ),
.I4(CLBLM_L_X72Y111_SLICE_X108Y111_AO6),
.I5(CLBLL_R_X71Y111_SLICE_X107Y111_AQ),
.O5(CLBLL_R_X71Y112_SLICE_X106Y112_AO5),
.O6(CLBLL_R_X71Y112_SLICE_X106Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y112_SLICE_X107Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y112_SLICE_X107Y112_DO5),
.O6(CLBLL_R_X71Y112_SLICE_X107Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y112_SLICE_X107Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y112_SLICE_X107Y112_CO5),
.O6(CLBLL_R_X71Y112_SLICE_X107Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y112_SLICE_X107Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y112_SLICE_X107Y112_BO5),
.O6(CLBLL_R_X71Y112_SLICE_X107Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y112_SLICE_X107Y112_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y112_SLICE_X107Y112_AO5),
.O6(CLBLL_R_X71Y112_SLICE_X107Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y114_SLICE_X106Y114_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y110_SLICE_X106Y110_A5Q),
.Q(CLBLL_R_X71Y114_SLICE_X106Y114_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y114_SLICE_X106Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y114_SLICE_X106Y114_DO5),
.O6(CLBLL_R_X71Y114_SLICE_X106Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y114_SLICE_X106Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y114_SLICE_X106Y114_CO5),
.O6(CLBLL_R_X71Y114_SLICE_X106Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y114_SLICE_X106Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y114_SLICE_X106Y114_BO5),
.O6(CLBLL_R_X71Y114_SLICE_X106Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y114_SLICE_X106Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y114_SLICE_X106Y114_AO5),
.O6(CLBLL_R_X71Y114_SLICE_X106Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y114_SLICE_X107Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y114_SLICE_X107Y114_DO5),
.O6(CLBLL_R_X71Y114_SLICE_X107Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y114_SLICE_X107Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y114_SLICE_X107Y114_CO5),
.O6(CLBLL_R_X71Y114_SLICE_X107Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y114_SLICE_X107Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y114_SLICE_X107Y114_BO5),
.O6(CLBLL_R_X71Y114_SLICE_X107Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y114_SLICE_X107Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y114_SLICE_X107Y114_AO5),
.O6(CLBLL_R_X71Y114_SLICE_X107Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y117_SLICE_X106Y117_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y117_SLICE_X106Y117_AO5),
.Q(CLBLL_R_X71Y117_SLICE_X106Y117_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y117_SLICE_X106Y117_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y117_SLICE_X106Y117_BO5),
.Q(CLBLL_R_X71Y117_SLICE_X106Y117_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y117_SLICE_X106Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y117_SLICE_X106Y117_AO6),
.Q(CLBLL_R_X71Y117_SLICE_X106Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y117_SLICE_X106Y117_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y117_SLICE_X106Y117_BO6),
.Q(CLBLL_R_X71Y117_SLICE_X106Y117_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y117_SLICE_X106Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y117_SLICE_X106Y117_DO5),
.O6(CLBLL_R_X71Y117_SLICE_X106Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y117_SLICE_X106Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y117_SLICE_X106Y117_CO5),
.O6(CLBLL_R_X71Y117_SLICE_X106Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafad8d8aa00aa00)
  ) CLBLL_R_X71Y117_SLICE_X106Y117_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X71Y117_SLICE_X106Y117_BQ),
.I2(CLBLL_R_X71Y117_SLICE_X106Y117_AQ),
.I3(CLBLM_R_X67Y111_SLICE_X100Y111_A5Q),
.I4(CLBLM_L_X68Y105_SLICE_X102Y105_DO6),
.I5(1'b1),
.O5(CLBLL_R_X71Y117_SLICE_X106Y117_BO5),
.O6(CLBLL_R_X71Y117_SLICE_X106Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccf3c088888888)
  ) CLBLL_R_X71Y117_SLICE_X106Y117_ALUT (
.I0(CLBLL_R_X71Y109_SLICE_X106Y109_B5Q),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLL_R_X71Y117_SLICE_X106Y117_AQ),
.I3(CLBLM_L_X72Y123_SLICE_X108Y123_A5Q),
.I4(CLBLM_L_X68Y107_SLICE_X103Y107_AO6),
.I5(1'b1),
.O5(CLBLL_R_X71Y117_SLICE_X106Y117_AO5),
.O6(CLBLL_R_X71Y117_SLICE_X106Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y117_SLICE_X107Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y117_SLICE_X107Y117_DO5),
.O6(CLBLL_R_X71Y117_SLICE_X107Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y117_SLICE_X107Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y117_SLICE_X107Y117_CO5),
.O6(CLBLL_R_X71Y117_SLICE_X107Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y117_SLICE_X107Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y117_SLICE_X107Y117_BO5),
.O6(CLBLL_R_X71Y117_SLICE_X107Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y117_SLICE_X107Y117_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y117_SLICE_X107Y117_AO5),
.O6(CLBLL_R_X71Y117_SLICE_X107Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y119_SLICE_X106Y119_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y119_SLICE_X106Y119_AO5),
.Q(CLBLL_R_X71Y119_SLICE_X106Y119_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y119_SLICE_X106Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y119_SLICE_X106Y119_AO6),
.Q(CLBLL_R_X71Y119_SLICE_X106Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y119_SLICE_X106Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y119_SLICE_X106Y119_DO5),
.O6(CLBLL_R_X71Y119_SLICE_X106Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y119_SLICE_X106Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y119_SLICE_X106Y119_CO5),
.O6(CLBLL_R_X71Y119_SLICE_X106Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y119_SLICE_X106Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y119_SLICE_X106Y119_BO5),
.O6(CLBLL_R_X71Y119_SLICE_X106Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4e455ffaa00)
  ) CLBLL_R_X71Y119_SLICE_X106Y119_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X71Y124_SLICE_X106Y124_A5Q),
.I2(CLBLL_R_X71Y125_SLICE_X106Y125_DO6),
.I3(CLBLL_R_X71Y110_SLICE_X106Y110_A5Q),
.I4(CLBLL_R_X71Y114_SLICE_X106Y114_AQ),
.I5(1'b1),
.O5(CLBLL_R_X71Y119_SLICE_X106Y119_AO5),
.O6(CLBLL_R_X71Y119_SLICE_X106Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y119_SLICE_X107Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y119_SLICE_X107Y119_DO5),
.O6(CLBLL_R_X71Y119_SLICE_X107Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y119_SLICE_X107Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y119_SLICE_X107Y119_CO5),
.O6(CLBLL_R_X71Y119_SLICE_X107Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y119_SLICE_X107Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y119_SLICE_X107Y119_BO5),
.O6(CLBLL_R_X71Y119_SLICE_X107Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y119_SLICE_X107Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y119_SLICE_X107Y119_AO5),
.O6(CLBLL_R_X71Y119_SLICE_X107Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y121_SLICE_X106Y121_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y121_SLICE_X106Y121_BO5),
.Q(CLBLL_R_X71Y121_SLICE_X106Y121_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y121_SLICE_X106Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y121_SLICE_X106Y121_AO6),
.Q(CLBLL_R_X71Y121_SLICE_X106Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y121_SLICE_X106Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y121_SLICE_X106Y121_DO5),
.O6(CLBLL_R_X71Y121_SLICE_X106Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y121_SLICE_X106Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y121_SLICE_X106Y121_CO5),
.O6(CLBLL_R_X71Y121_SLICE_X106Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaffaafcfcb8b8)
  ) CLBLL_R_X71Y121_SLICE_X106Y121_BLUT (
.I0(CLBLL_R_X71Y126_SLICE_X107Y126_CO6),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_R_X63Y122_SLICE_X95Y122_CQ),
.I3(CLBLL_R_X83Y94_SLICE_X130Y94_AQ),
.I4(CLBLL_R_X71Y121_SLICE_X106Y121_A5Q),
.I5(1'b1),
.O5(CLBLL_R_X71Y121_SLICE_X106Y121_BO5),
.O6(CLBLL_R_X71Y121_SLICE_X106Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffccccfffbccc8)
  ) CLBLL_R_X71Y121_SLICE_X106Y121_ALUT (
.I0(CLBLM_L_X72Y123_SLICE_X108Y123_CO6),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_L_X68Y107_SLICE_X103Y107_AO6),
.I3(CLBLL_R_X71Y121_SLICE_X106Y121_BO6),
.I4(CLBLM_L_X72Y118_SLICE_X108Y118_AQ),
.I5(CLBLM_L_X68Y105_SLICE_X102Y105_DO6),
.O5(CLBLL_R_X71Y121_SLICE_X106Y121_AO5),
.O6(CLBLL_R_X71Y121_SLICE_X106Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y121_SLICE_X107Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y121_SLICE_X107Y121_DO5),
.O6(CLBLL_R_X71Y121_SLICE_X107Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y121_SLICE_X107Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y121_SLICE_X107Y121_CO5),
.O6(CLBLL_R_X71Y121_SLICE_X107Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y121_SLICE_X107Y121_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y121_SLICE_X107Y121_BO5),
.O6(CLBLL_R_X71Y121_SLICE_X107Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y121_SLICE_X107Y121_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y121_SLICE_X107Y121_AO5),
.O6(CLBLL_R_X71Y121_SLICE_X107Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y124_SLICE_X106Y124_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y124_SLICE_X106Y124_AO5),
.Q(CLBLL_R_X71Y124_SLICE_X106Y124_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y124_SLICE_X106Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y124_SLICE_X106Y124_AO6),
.Q(CLBLL_R_X71Y124_SLICE_X106Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y124_SLICE_X106Y124_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y124_SLICE_X106Y124_BO5),
.Q(CLBLL_R_X71Y124_SLICE_X106Y124_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y124_SLICE_X106Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y124_SLICE_X106Y124_DO5),
.O6(CLBLL_R_X71Y124_SLICE_X106Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0054005500000000)
  ) CLBLL_R_X71Y124_SLICE_X106Y124_CLUT (
.I0(CLBLL_R_X71Y126_SLICE_X107Y126_AQ),
.I1(CLBLL_R_X71Y126_SLICE_X107Y126_BQ),
.I2(CLBLM_L_X70Y123_SLICE_X104Y123_AQ),
.I3(CLBLM_L_X70Y124_SLICE_X105Y124_BO6),
.I4(CLBLM_L_X70Y126_SLICE_X104Y126_CQ),
.I5(CLBLM_L_X70Y125_SLICE_X105Y125_AQ),
.O5(CLBLL_R_X71Y124_SLICE_X106Y124_CO5),
.O6(CLBLL_R_X71Y124_SLICE_X106Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffafffafdfffd0f0)
  ) CLBLL_R_X71Y124_SLICE_X106Y124_BLUT (
.I0(CLBLL_R_X73Y125_SLICE_X110Y125_DO6),
.I1(CLBLL_R_X71Y124_SLICE_X106Y124_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLL_R_X71Y129_SLICE_X107Y129_BO6),
.I4(CLBLL_R_X71Y117_SLICE_X106Y117_BQ),
.I5(1'b1),
.O5(CLBLL_R_X71Y124_SLICE_X106Y124_BO5),
.O6(CLBLL_R_X71Y124_SLICE_X106Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88bb88fcfc3030)
  ) CLBLL_R_X71Y124_SLICE_X106Y124_ALUT (
.I0(CLBLM_L_X70Y125_SLICE_X105Y125_CO6),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_L_X70Y124_SLICE_X104Y124_BQ),
.I3(CLBLL_R_X73Y125_SLICE_X111Y125_A5Q),
.I4(CLBLL_R_X71Y125_SLICE_X106Y125_DO6),
.I5(1'b1),
.O5(CLBLL_R_X71Y124_SLICE_X106Y124_AO5),
.O6(CLBLL_R_X71Y124_SLICE_X106Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y124_SLICE_X107Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y124_SLICE_X107Y124_DO5),
.O6(CLBLL_R_X71Y124_SLICE_X107Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y124_SLICE_X107Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y124_SLICE_X107Y124_CO5),
.O6(CLBLL_R_X71Y124_SLICE_X107Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y124_SLICE_X107Y124_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y124_SLICE_X107Y124_BO5),
.O6(CLBLL_R_X71Y124_SLICE_X107Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y124_SLICE_X107Y124_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y124_SLICE_X107Y124_AO5),
.O6(CLBLL_R_X71Y124_SLICE_X107Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y125_SLICE_X106Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y125_SLICE_X106Y125_AO6),
.Q(CLBLL_R_X71Y125_SLICE_X106Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y125_SLICE_X106Y125_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y125_SLICE_X106Y125_BO6),
.Q(CLBLL_R_X71Y125_SLICE_X106Y125_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y125_SLICE_X106Y125_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y125_SLICE_X106Y125_CO6),
.Q(CLBLL_R_X71Y125_SLICE_X106Y125_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fcfff0f0fdfd)
  ) CLBLL_R_X71Y125_SLICE_X106Y125_DLUT (
.I0(CLBLM_L_X70Y124_SLICE_X104Y124_BQ),
.I1(CLBLL_R_X71Y126_SLICE_X107Y126_AQ),
.I2(CLBLL_R_X71Y125_SLICE_X107Y125_DO6),
.I3(CLBLM_L_X70Y126_SLICE_X104Y126_CQ),
.I4(CLBLL_R_X71Y126_SLICE_X106Y126_DO6),
.I5(CLBLM_L_X70Y125_SLICE_X105Y125_AQ),
.O5(CLBLL_R_X71Y125_SLICE_X106Y125_DO5),
.O6(CLBLL_R_X71Y125_SLICE_X106Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccdd0000fcfdf0f0)
  ) CLBLL_R_X71Y125_SLICE_X106Y125_CLUT (
.I0(CLBLL_R_X71Y132_SLICE_X107Y132_BQ),
.I1(CLBLL_R_X71Y125_SLICE_X106Y125_CQ),
.I2(CLBLL_R_X71Y125_SLICE_X106Y125_BQ),
.I3(CLBLM_L_X70Y125_SLICE_X105Y125_BO6),
.I4(CLBLM_L_X70Y125_SLICE_X105Y125_AO5),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLL_R_X71Y125_SLICE_X106Y125_CO5),
.O6(CLBLL_R_X71Y125_SLICE_X106Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888ff888a8aff8a)
  ) CLBLL_R_X71Y125_SLICE_X106Y125_BLUT (
.I0(CLBLM_L_X70Y125_SLICE_X105Y125_AO5),
.I1(CLBLL_R_X71Y125_SLICE_X106Y125_BQ),
.I2(CLBLM_L_X70Y125_SLICE_X105Y125_BO6),
.I3(CLBLM_L_X70Y126_SLICE_X104Y126_BQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X71Y130_SLICE_X106Y130_CQ),
.O5(CLBLL_R_X71Y125_SLICE_X106Y125_BO5),
.O6(CLBLL_R_X71Y125_SLICE_X106Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a077772222)
  ) CLBLL_R_X71Y125_SLICE_X106Y125_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X71Y125_SLICE_X106Y125_BQ),
.I2(CLBLL_R_X71Y125_SLICE_X106Y125_AQ),
.I3(1'b1),
.I4(CLBLL_R_X71Y125_SLICE_X107Y125_AQ),
.I5(CLBLM_L_X70Y124_SLICE_X105Y124_CO6),
.O5(CLBLL_R_X71Y125_SLICE_X106Y125_AO5),
.O6(CLBLL_R_X71Y125_SLICE_X106Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y125_SLICE_X107Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y125_SLICE_X107Y125_AO6),
.Q(CLBLL_R_X71Y125_SLICE_X107Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000f0a00000f0c)
  ) CLBLL_R_X71Y125_SLICE_X107Y125_DLUT (
.I0(CLBLM_L_X72Y123_SLICE_X108Y123_AQ),
.I1(CLBLM_L_X72Y125_SLICE_X108Y125_AQ),
.I2(CLBLL_R_X71Y126_SLICE_X107Y126_BO5),
.I3(CLBLL_R_X71Y126_SLICE_X107Y126_AQ),
.I4(CLBLM_L_X70Y124_SLICE_X105Y124_DO6),
.I5(CLBLM_L_X70Y125_SLICE_X105Y125_AQ),
.O5(CLBLL_R_X71Y125_SLICE_X107Y125_DO5),
.O6(CLBLL_R_X71Y125_SLICE_X107Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5000500040005000)
  ) CLBLL_R_X71Y125_SLICE_X107Y125_CLUT (
.I0(CLBLM_L_X70Y124_SLICE_X105Y124_BO6),
.I1(CLBLM_L_X70Y123_SLICE_X104Y123_AQ),
.I2(CLBLM_L_X70Y125_SLICE_X105Y125_AQ),
.I3(CLBLL_R_X71Y126_SLICE_X107Y126_AQ),
.I4(CLBLL_R_X71Y125_SLICE_X107Y125_AQ),
.I5(CLBLL_R_X71Y126_SLICE_X107Y126_BQ),
.O5(CLBLL_R_X71Y125_SLICE_X107Y125_CO5),
.O6(CLBLL_R_X71Y125_SLICE_X107Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0050005000400050)
  ) CLBLL_R_X71Y125_SLICE_X107Y125_BLUT (
.I0(CLBLM_L_X70Y125_SLICE_X105Y125_AQ),
.I1(CLBLM_L_X70Y123_SLICE_X104Y123_AQ),
.I2(CLBLL_R_X71Y126_SLICE_X107Y126_AQ),
.I3(CLBLM_L_X70Y124_SLICE_X105Y124_BO6),
.I4(CLBLL_R_X71Y125_SLICE_X106Y125_AQ),
.I5(CLBLL_R_X71Y126_SLICE_X107Y126_BQ),
.O5(CLBLL_R_X71Y125_SLICE_X107Y125_BO5),
.O6(CLBLL_R_X71Y125_SLICE_X107Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafaf2fafa0a0e0a0)
  ) CLBLL_R_X71Y125_SLICE_X107Y125_ALUT (
.I0(CLBLL_R_X71Y125_SLICE_X107Y125_AQ),
.I1(CLBLM_L_X70Y123_SLICE_X104Y123_AQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLL_R_X71Y126_SLICE_X107Y126_BQ),
.I4(CLBLM_L_X70Y125_SLICE_X105Y125_BO5),
.I5(CLBLL_R_X71Y125_SLICE_X106Y125_CQ),
.O5(CLBLL_R_X71Y125_SLICE_X107Y125_AO5),
.O6(CLBLL_R_X71Y125_SLICE_X107Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y126_SLICE_X106Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y126_SLICE_X106Y126_AO6),
.Q(CLBLL_R_X71Y126_SLICE_X106Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y126_SLICE_X106Y126_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y126_SLICE_X106Y126_BO6),
.Q(CLBLL_R_X71Y126_SLICE_X106Y126_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha2ffa2ff80ff80ff)
  ) CLBLL_R_X71Y126_SLICE_X106Y126_DLUT (
.I0(CLBLL_R_X71Y126_SLICE_X107Y126_AQ),
.I1(CLBLM_L_X70Y125_SLICE_X105Y125_AQ),
.I2(CLBLL_R_X71Y126_SLICE_X106Y126_AQ),
.I3(CLBLM_L_X70Y124_SLICE_X105Y124_DO6),
.I4(1'b1),
.I5(CLBLM_L_X70Y126_SLICE_X105Y126_AQ),
.O5(CLBLL_R_X71Y126_SLICE_X106Y126_DO5),
.O6(CLBLL_R_X71Y126_SLICE_X106Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0500040005000500)
  ) CLBLL_R_X71Y126_SLICE_X106Y126_CLUT (
.I0(CLBLM_L_X70Y124_SLICE_X105Y124_BO6),
.I1(CLBLM_L_X70Y123_SLICE_X104Y123_AQ),
.I2(CLBLM_L_X70Y125_SLICE_X105Y125_AQ),
.I3(CLBLL_R_X71Y126_SLICE_X107Y126_AQ),
.I4(CLBLL_R_X71Y126_SLICE_X107Y126_BQ),
.I5(CLBLM_L_X70Y126_SLICE_X105Y126_AQ),
.O5(CLBLL_R_X71Y126_SLICE_X106Y126_CO5),
.O6(CLBLL_R_X71Y126_SLICE_X106Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcd00cd00ffffcd00)
  ) CLBLL_R_X71Y126_SLICE_X106Y126_BLUT (
.I0(CLBLM_L_X72Y128_SLICE_X108Y128_AQ),
.I1(CLBLL_R_X71Y126_SLICE_X106Y126_BQ),
.I2(CLBLM_L_X70Y125_SLICE_X105Y125_BO6),
.I3(CLBLM_L_X70Y125_SLICE_X105Y125_AO5),
.I4(CLBLM_L_X70Y126_SLICE_X105Y126_BQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLL_R_X71Y126_SLICE_X106Y126_BO5),
.O6(CLBLL_R_X71Y126_SLICE_X106Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e466e4e4e4e4e4)
  ) CLBLL_R_X71Y126_SLICE_X106Y126_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X71Y126_SLICE_X106Y126_BQ),
.I2(CLBLL_R_X71Y126_SLICE_X106Y126_AQ),
.I3(CLBLL_R_X71Y126_SLICE_X107Y126_BQ),
.I4(CLBLM_L_X70Y125_SLICE_X105Y125_BO5),
.I5(CLBLM_L_X70Y123_SLICE_X104Y123_AQ),
.O5(CLBLL_R_X71Y126_SLICE_X106Y126_AO5),
.O6(CLBLL_R_X71Y126_SLICE_X106Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y126_SLICE_X107Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y126_SLICE_X107Y126_AO6),
.Q(CLBLL_R_X71Y126_SLICE_X107Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y126_SLICE_X107Y126_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y126_SLICE_X107Y126_BO6),
.Q(CLBLL_R_X71Y126_SLICE_X107Y126_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccc8ccccccc8)
  ) CLBLL_R_X71Y126_SLICE_X107Y126_DLUT (
.I0(CLBLL_R_X73Y124_SLICE_X111Y124_BQ),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_L_X72Y128_SLICE_X108Y128_DQ),
.I3(CLBLM_L_X72Y125_SLICE_X109Y125_AQ),
.I4(CLBLL_R_X71Y127_SLICE_X107Y127_DQ),
.I5(1'b1),
.O5(CLBLL_R_X71Y126_SLICE_X107Y126_DO5),
.O6(CLBLL_R_X71Y126_SLICE_X107Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccc8cccccccc)
  ) CLBLL_R_X71Y126_SLICE_X107Y126_CLUT (
.I0(CLBLL_R_X73Y124_SLICE_X111Y124_BQ),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLL_R_X71Y127_SLICE_X107Y127_DQ),
.I3(CLBLM_L_X72Y125_SLICE_X109Y125_AQ),
.I4(CLBLM_L_X72Y128_SLICE_X108Y128_DQ),
.I5(CLBLL_R_X71Y130_SLICE_X106Y130_DO5),
.O5(CLBLL_R_X71Y126_SLICE_X107Y126_CO5),
.O6(CLBLL_R_X71Y126_SLICE_X107Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000f0f050305030)
  ) CLBLL_R_X71Y126_SLICE_X107Y126_BLUT (
.I0(CLBLM_L_X72Y127_SLICE_X108Y127_CQ),
.I1(CLBLL_R_X71Y127_SLICE_X107Y127_BQ),
.I2(CLBLL_R_X71Y126_SLICE_X107Y126_AQ),
.I3(CLBLM_L_X70Y125_SLICE_X105Y125_AQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLL_R_X71Y126_SLICE_X107Y126_BO5),
.O6(CLBLL_R_X71Y126_SLICE_X107Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaaaa1b001b00)
  ) CLBLL_R_X71Y126_SLICE_X107Y126_ALUT (
.I0(CLBLM_L_X70Y125_SLICE_X105Y125_AQ),
.I1(CLBLM_L_X72Y129_SLICE_X108Y129_BQ),
.I2(CLBLL_R_X71Y132_SLICE_X107Y132_CQ),
.I3(CLBLL_R_X71Y126_SLICE_X107Y126_AQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLL_R_X71Y126_SLICE_X107Y126_AO5),
.O6(CLBLL_R_X71Y126_SLICE_X107Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y127_SLICE_X106Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y127_SLICE_X106Y127_DO5),
.O6(CLBLL_R_X71Y127_SLICE_X106Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y127_SLICE_X106Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y127_SLICE_X106Y127_CO5),
.O6(CLBLL_R_X71Y127_SLICE_X106Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y127_SLICE_X106Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y127_SLICE_X106Y127_BO5),
.O6(CLBLL_R_X71Y127_SLICE_X106Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y127_SLICE_X106Y127_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y127_SLICE_X106Y127_AO5),
.O6(CLBLL_R_X71Y127_SLICE_X106Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y127_SLICE_X107Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y127_SLICE_X107Y127_AO6),
.Q(CLBLL_R_X71Y127_SLICE_X107Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y127_SLICE_X107Y127_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y127_SLICE_X107Y127_BO6),
.Q(CLBLL_R_X71Y127_SLICE_X107Y127_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y127_SLICE_X107Y127_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y127_SLICE_X107Y127_CO6),
.Q(CLBLL_R_X71Y127_SLICE_X107Y127_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y127_SLICE_X107Y127_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y127_SLICE_X107Y127_DO6),
.Q(CLBLL_R_X71Y127_SLICE_X107Y127_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff3ccccc003ccccc)
  ) CLBLL_R_X71Y127_SLICE_X107Y127_DLUT (
.I0(1'b1),
.I1(CLBLL_R_X71Y127_SLICE_X107Y127_CQ),
.I2(CLBLL_R_X75Y127_SLICE_X114Y127_DQ),
.I3(CLBLL_R_X71Y127_SLICE_X107Y127_AO5),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X71Y127_SLICE_X107Y127_DQ),
.O5(CLBLL_R_X71Y127_SLICE_X107Y127_DO5),
.O6(CLBLL_R_X71Y127_SLICE_X107Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6aaa6a6acacacaca)
  ) CLBLL_R_X71Y127_SLICE_X107Y127_CLUT (
.I0(CLBLL_R_X71Y127_SLICE_X107Y127_BQ),
.I1(CLBLL_R_X71Y127_SLICE_X107Y127_CQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X72Y126_SLICE_X109Y126_AQ),
.I4(CLBLL_R_X71Y127_SLICE_X107Y127_AQ),
.I5(CLBLL_R_X71Y126_SLICE_X106Y126_CO6),
.O5(CLBLL_R_X71Y127_SLICE_X107Y127_CO5),
.O6(CLBLL_R_X71Y127_SLICE_X107Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ccccaaaaaaaa)
  ) CLBLL_R_X71Y127_SLICE_X107Y127_BLUT (
.I0(CLBLL_R_X73Y126_SLICE_X110Y126_A5Q),
.I1(CLBLL_R_X71Y127_SLICE_X107Y127_BQ),
.I2(1'b1),
.I3(CLBLM_L_X72Y127_SLICE_X109Y127_AO6),
.I4(CLBLL_R_X71Y126_SLICE_X106Y126_CO6),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLL_R_X71Y127_SLICE_X107Y127_BO5),
.O6(CLBLL_R_X71Y127_SLICE_X107Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff500a0ffff0fff)
  ) CLBLL_R_X71Y127_SLICE_X107Y127_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(1'b1),
.I2(CLBLL_R_X71Y127_SLICE_X107Y127_AQ),
.I3(CLBLL_R_X71Y126_SLICE_X106Y126_CO6),
.I4(CLBLM_L_X72Y126_SLICE_X109Y126_AQ),
.I5(1'b1),
.O5(CLBLL_R_X71Y127_SLICE_X107Y127_AO5),
.O6(CLBLL_R_X71Y127_SLICE_X107Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y128_SLICE_X106Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y128_SLICE_X106Y128_AO6),
.Q(CLBLL_R_X71Y128_SLICE_X106Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y128_SLICE_X106Y128_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y128_SLICE_X106Y128_BO6),
.Q(CLBLL_R_X71Y128_SLICE_X106Y128_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y128_SLICE_X106Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y128_SLICE_X106Y128_DO5),
.O6(CLBLL_R_X71Y128_SLICE_X106Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha000a000a000a000)
  ) CLBLL_R_X71Y128_SLICE_X106Y128_CLUT (
.I0(CLBLM_L_X70Y128_SLICE_X104Y128_BQ),
.I1(1'b1),
.I2(CLBLM_L_X70Y129_SLICE_X104Y129_AQ),
.I3(CLBLM_L_X70Y126_SLICE_X105Y126_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y128_SLICE_X106Y128_CO5),
.O6(CLBLL_R_X71Y128_SLICE_X106Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a5f0f0ccccf0f0)
  ) CLBLL_R_X71Y128_SLICE_X106Y128_BLUT (
.I0(CLBLM_L_X70Y129_SLICE_X105Y129_DQ),
.I1(CLBLL_R_X71Y128_SLICE_X106Y128_BQ),
.I2(CLBLL_R_X71Y128_SLICE_X106Y128_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X71Y128_SLICE_X106Y128_CO6),
.O5(CLBLL_R_X71Y128_SLICE_X106Y128_BO5),
.O6(CLBLL_R_X71Y128_SLICE_X106Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haae2e2e2e2e2e2e2)
  ) CLBLL_R_X71Y128_SLICE_X106Y128_ALUT (
.I0(CLBLM_L_X70Y129_SLICE_X105Y129_DQ),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLL_R_X71Y128_SLICE_X106Y128_AQ),
.I3(CLBLM_L_X70Y126_SLICE_X105Y126_CO6),
.I4(CLBLM_L_X70Y128_SLICE_X104Y128_BQ),
.I5(CLBLM_L_X70Y129_SLICE_X104Y129_AQ),
.O5(CLBLL_R_X71Y128_SLICE_X106Y128_AO5),
.O6(CLBLL_R_X71Y128_SLICE_X106Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y128_SLICE_X107Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y128_SLICE_X107Y128_DO5),
.O6(CLBLL_R_X71Y128_SLICE_X107Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y128_SLICE_X107Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y128_SLICE_X107Y128_CO5),
.O6(CLBLL_R_X71Y128_SLICE_X107Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y128_SLICE_X107Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y128_SLICE_X107Y128_BO5),
.O6(CLBLL_R_X71Y128_SLICE_X107Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y128_SLICE_X107Y128_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y128_SLICE_X107Y128_AO5),
.O6(CLBLL_R_X71Y128_SLICE_X107Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y129_SLICE_X106Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y129_SLICE_X106Y129_AO5),
.Q(CLBLL_R_X71Y129_SLICE_X106Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y129_SLICE_X106Y129_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y129_SLICE_X106Y129_BO6),
.Q(CLBLL_R_X71Y129_SLICE_X106Y129_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y129_SLICE_X106Y129_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y129_SLICE_X106Y129_CO6),
.Q(CLBLL_R_X71Y129_SLICE_X106Y129_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800880088008800)
  ) CLBLL_R_X71Y129_SLICE_X106Y129_DLUT (
.I0(CLBLL_R_X71Y125_SLICE_X107Y125_BO6),
.I1(CLBLL_R_X71Y129_SLICE_X106Y129_AQ),
.I2(1'b1),
.I3(CLBLL_R_X71Y130_SLICE_X106Y130_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y129_SLICE_X106Y129_DO5),
.O6(CLBLL_R_X71Y129_SLICE_X106Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf05ad8d8f05ad8d8)
  ) CLBLL_R_X71Y129_SLICE_X106Y129_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X71Y129_SLICE_X106Y129_CQ),
.I2(CLBLL_R_X71Y129_SLICE_X106Y129_BQ),
.I3(CLBLM_L_X72Y130_SLICE_X109Y130_CQ),
.I4(CLBLL_R_X71Y129_SLICE_X106Y129_DO6),
.I5(1'b1),
.O5(CLBLL_R_X71Y129_SLICE_X106Y129_CO5),
.O6(CLBLL_R_X71Y129_SLICE_X106Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfaaffaa80aa00aa)
  ) CLBLL_R_X71Y129_SLICE_X106Y129_BLUT (
.I0(CLBLM_L_X72Y130_SLICE_X109Y130_CQ),
.I1(CLBLL_R_X71Y130_SLICE_X106Y130_BQ),
.I2(CLBLL_R_X71Y129_SLICE_X106Y129_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLL_R_X71Y125_SLICE_X107Y125_BO6),
.I5(CLBLL_R_X71Y129_SLICE_X106Y129_BQ),
.O5(CLBLL_R_X71Y129_SLICE_X106Y129_BO5),
.O6(CLBLL_R_X71Y129_SLICE_X106Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f5f5b8b8ff00)
  ) CLBLL_R_X71Y129_SLICE_X106Y129_ALUT (
.I0(CLBLM_L_X72Y129_SLICE_X108Y129_AQ),
.I1(CLBLL_R_X71Y125_SLICE_X107Y125_BO6),
.I2(CLBLL_R_X71Y129_SLICE_X106Y129_AQ),
.I3(CLBLL_R_X71Y129_SLICE_X107Y129_BQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLL_R_X71Y129_SLICE_X106Y129_AO5),
.O6(CLBLL_R_X71Y129_SLICE_X106Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y129_SLICE_X107Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y130_SLICE_X105Y130_AQ),
.Q(CLBLL_R_X71Y129_SLICE_X107Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y129_SLICE_X107Y129_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y129_SLICE_X108Y129_AQ),
.Q(CLBLL_R_X71Y129_SLICE_X107Y129_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y129_SLICE_X107Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y129_SLICE_X107Y129_DO5),
.O6(CLBLL_R_X71Y129_SLICE_X107Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffafa)
  ) CLBLL_R_X71Y129_SLICE_X107Y129_CLUT (
.I0(CLBLL_R_X71Y130_SLICE_X107Y130_BQ),
.I1(1'b1),
.I2(CLBLL_R_X71Y129_SLICE_X107Y129_BQ),
.I3(1'b1),
.I4(CLBLM_L_X70Y128_SLICE_X105Y128_AQ),
.I5(CLBLM_L_X70Y132_SLICE_X105Y132_AQ),
.O5(CLBLL_R_X71Y129_SLICE_X107Y129_CO5),
.O6(CLBLL_R_X71Y129_SLICE_X107Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000101)
  ) CLBLL_R_X71Y129_SLICE_X107Y129_BLUT (
.I0(CLBLM_L_X72Y132_SLICE_X109Y132_AQ),
.I1(CLBLM_L_X70Y132_SLICE_X105Y132_BQ),
.I2(CLBLL_R_X71Y129_SLICE_X107Y129_AQ),
.I3(1'b1),
.I4(CLBLL_R_X71Y130_SLICE_X107Y130_AQ),
.I5(CLBLL_R_X71Y129_SLICE_X107Y129_CO6),
.O5(CLBLL_R_X71Y129_SLICE_X107Y129_BO5),
.O6(CLBLL_R_X71Y129_SLICE_X107Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0f0f0f0e0)
  ) CLBLL_R_X71Y129_SLICE_X107Y129_ALUT (
.I0(CLBLL_R_X71Y130_SLICE_X107Y130_DO6),
.I1(CLBLM_L_X72Y130_SLICE_X109Y130_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLL_R_X71Y128_SLICE_X106Y128_BQ),
.I4(CLBLL_R_X71Y133_SLICE_X106Y133_DQ),
.I5(CLBLL_R_X71Y129_SLICE_X106Y129_CQ),
.O5(CLBLL_R_X71Y129_SLICE_X107Y129_AO5),
.O6(CLBLL_R_X71Y129_SLICE_X107Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y130_SLICE_X106Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y130_SLICE_X106Y130_AO5),
.Q(CLBLL_R_X71Y130_SLICE_X106Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y130_SLICE_X106Y130_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y130_SLICE_X106Y130_BO6),
.Q(CLBLL_R_X71Y130_SLICE_X106Y130_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y130_SLICE_X106Y130_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y130_SLICE_X106Y130_CO6),
.Q(CLBLL_R_X71Y130_SLICE_X106Y130_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333700000005)
  ) CLBLL_R_X71Y130_SLICE_X106Y130_DLUT (
.I0(CLBLM_L_X70Y129_SLICE_X104Y129_CQ),
.I1(CLBLL_R_X71Y126_SLICE_X107Y126_DO6),
.I2(CLBLM_L_X72Y130_SLICE_X108Y130_CQ),
.I3(CLBLL_R_X71Y132_SLICE_X106Y132_BQ),
.I4(CLBLM_L_X70Y133_SLICE_X105Y133_DQ),
.I5(1'b1),
.O5(CLBLL_R_X71Y130_SLICE_X106Y130_DO5),
.O6(CLBLL_R_X71Y130_SLICE_X106Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa3a0a3afafa0a0a)
  ) CLBLL_R_X71Y130_SLICE_X106Y130_CLUT (
.I0(CLBLL_R_X71Y131_SLICE_X107Y131_AQ),
.I1(CLBLM_L_X72Y130_SLICE_X108Y130_AO6),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLL_R_X71Y129_SLICE_X106Y129_AO6),
.I4(CLBLL_R_X71Y130_SLICE_X106Y130_CQ),
.I5(CLBLL_R_X71Y125_SLICE_X107Y125_BO6),
.O5(CLBLL_R_X71Y130_SLICE_X106Y130_CO5),
.O6(CLBLL_R_X71Y130_SLICE_X106Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ccaaaacfccaaaa)
  ) CLBLL_R_X71Y130_SLICE_X106Y130_BLUT (
.I0(CLBLL_R_X71Y130_SLICE_X106Y130_CQ),
.I1(CLBLL_R_X71Y130_SLICE_X106Y130_BQ),
.I2(CLBLM_L_X72Y129_SLICE_X108Y129_AQ),
.I3(CLBLL_R_X71Y125_SLICE_X107Y125_BO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X71Y129_SLICE_X106Y129_AQ),
.O5(CLBLL_R_X71Y130_SLICE_X106Y130_BO5),
.O6(CLBLL_R_X71Y130_SLICE_X106Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f000f0f5a0cccc)
  ) CLBLL_R_X71Y130_SLICE_X106Y130_ALUT (
.I0(CLBLM_L_X72Y132_SLICE_X109Y132_AO6),
.I1(CLBLL_R_X71Y129_SLICE_X107Y129_AQ),
.I2(CLBLL_R_X71Y130_SLICE_X106Y130_AQ),
.I3(CLBLM_L_X70Y130_SLICE_X105Y130_AQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLL_R_X71Y130_SLICE_X106Y130_AO5),
.O6(CLBLL_R_X71Y130_SLICE_X106Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y130_SLICE_X107Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y131_SLICE_X108Y131_AQ),
.Q(CLBLL_R_X71Y130_SLICE_X107Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y130_SLICE_X107Y130_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y132_SLICE_X106Y132_AQ),
.Q(CLBLL_R_X71Y130_SLICE_X107Y130_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffefefefe)
  ) CLBLL_R_X71Y130_SLICE_X107Y130_DLUT (
.I0(CLBLL_R_X71Y133_SLICE_X107Y133_BQ),
.I1(CLBLM_L_X70Y130_SLICE_X104Y130_DQ),
.I2(CLBLL_R_X71Y131_SLICE_X106Y131_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_R_X71Y134_SLICE_X107Y134_BQ),
.O5(CLBLL_R_X71Y130_SLICE_X107Y130_DO5),
.O6(CLBLL_R_X71Y130_SLICE_X107Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaabbffbbffbbff)
  ) CLBLL_R_X71Y130_SLICE_X107Y130_CLUT (
.I0(CLBLM_L_X72Y129_SLICE_X108Y129_AQ),
.I1(CLBLL_R_X71Y129_SLICE_X106Y129_AQ),
.I2(1'b1),
.I3(CLBLM_L_X72Y131_SLICE_X108Y131_CQ),
.I4(CLBLL_R_X71Y131_SLICE_X107Y131_BQ),
.I5(CLBLL_R_X71Y130_SLICE_X106Y130_BQ),
.O5(CLBLL_R_X71Y130_SLICE_X107Y130_CO5),
.O6(CLBLL_R_X71Y130_SLICE_X107Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h50d050d000c000c0)
  ) CLBLL_R_X71Y130_SLICE_X107Y130_BLUT (
.I0(CLBLL_R_X71Y129_SLICE_X106Y129_AQ),
.I1(CLBLM_L_X72Y131_SLICE_X108Y131_BQ),
.I2(CLBLM_L_X72Y129_SLICE_X108Y129_AQ),
.I3(CLBLL_R_X71Y130_SLICE_X106Y130_BQ),
.I4(1'b1),
.I5(CLBLL_R_X71Y131_SLICE_X107Y131_CQ),
.O5(CLBLL_R_X71Y130_SLICE_X107Y130_BO5),
.O6(CLBLL_R_X71Y130_SLICE_X107Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff85ff80ffffffff)
  ) CLBLL_R_X71Y130_SLICE_X107Y130_ALUT (
.I0(CLBLL_R_X71Y129_SLICE_X106Y129_AQ),
.I1(CLBLM_L_X72Y131_SLICE_X109Y131_BQ),
.I2(CLBLL_R_X71Y130_SLICE_X106Y130_BQ),
.I3(CLBLL_R_X71Y130_SLICE_X107Y130_BO6),
.I4(CLBLL_R_X71Y131_SLICE_X107Y131_AQ),
.I5(CLBLL_R_X71Y130_SLICE_X107Y130_CO6),
.O5(CLBLL_R_X71Y130_SLICE_X107Y130_AO5),
.O6(CLBLL_R_X71Y130_SLICE_X107Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y131_SLICE_X106Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y131_SLICE_X106Y131_AO6),
.Q(CLBLL_R_X71Y131_SLICE_X106Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y131_SLICE_X106Y131_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y131_SLICE_X106Y131_BO6),
.Q(CLBLL_R_X71Y131_SLICE_X106Y131_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y131_SLICE_X106Y131_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y131_SLICE_X106Y131_CO6),
.Q(CLBLL_R_X71Y131_SLICE_X106Y131_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0000000000000)
  ) CLBLL_R_X71Y131_SLICE_X106Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_R_X71Y131_SLICE_X106Y131_AQ),
.I3(1'b1),
.I4(CLBLL_R_X71Y131_SLICE_X107Y131_A5Q),
.I5(CLBLL_R_X71Y125_SLICE_X107Y125_CO6),
.O5(CLBLL_R_X71Y131_SLICE_X106Y131_DO5),
.O6(CLBLL_R_X71Y131_SLICE_X106Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf50add88f50add88)
  ) CLBLL_R_X71Y131_SLICE_X106Y131_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X71Y131_SLICE_X106Y131_CQ),
.I2(CLBLL_R_X71Y132_SLICE_X106Y132_DQ),
.I3(CLBLL_R_X71Y131_SLICE_X106Y131_BQ),
.I4(CLBLL_R_X71Y131_SLICE_X106Y131_DO6),
.I5(1'b1),
.O5(CLBLL_R_X71Y131_SLICE_X106Y131_CO5),
.O6(CLBLL_R_X71Y131_SLICE_X106Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hecccffff4ccc0000)
  ) CLBLL_R_X71Y131_SLICE_X106Y131_BLUT (
.I0(CLBLL_R_X71Y131_SLICE_X107Y131_A5Q),
.I1(CLBLL_R_X71Y131_SLICE_X106Y131_BQ),
.I2(CLBLL_R_X71Y131_SLICE_X106Y131_AQ),
.I3(CLBLL_R_X71Y125_SLICE_X107Y125_CO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X71Y132_SLICE_X106Y132_DQ),
.O5(CLBLL_R_X71Y131_SLICE_X106Y131_BO5),
.O6(CLBLL_R_X71Y131_SLICE_X106Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h50f0cccc55f0cccc)
  ) CLBLL_R_X71Y131_SLICE_X106Y131_ALUT (
.I0(CLBLL_R_X71Y131_SLICE_X107Y131_A5Q),
.I1(CLBLL_R_X71Y132_SLICE_X107Y132_BQ),
.I2(CLBLL_R_X71Y131_SLICE_X106Y131_AQ),
.I3(CLBLL_R_X71Y125_SLICE_X107Y125_CO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X71Y132_SLICE_X106Y132_AQ),
.O5(CLBLL_R_X71Y131_SLICE_X106Y131_AO5),
.O6(CLBLL_R_X71Y131_SLICE_X106Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y131_SLICE_X107Y131_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y131_SLICE_X107Y131_DO5),
.Q(CLBLL_R_X71Y131_SLICE_X107Y131_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y131_SLICE_X107Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y131_SLICE_X107Y131_AO6),
.Q(CLBLL_R_X71Y131_SLICE_X107Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y131_SLICE_X107Y131_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y131_SLICE_X107Y131_BO6),
.Q(CLBLL_R_X71Y131_SLICE_X107Y131_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y131_SLICE_X107Y131_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y131_SLICE_X107Y131_CO6),
.Q(CLBLL_R_X71Y131_SLICE_X107Y131_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33ff33d8d8fa50)
  ) CLBLL_R_X71Y131_SLICE_X107Y131_DLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X71Y132_SLICE_X106Y132_AQ),
.I2(CLBLL_R_X71Y130_SLICE_X107Y130_BQ),
.I3(CLBLL_R_X71Y131_SLICE_X107Y131_A5Q),
.I4(CLBLL_R_X71Y125_SLICE_X107Y125_CO6),
.I5(1'b1),
.O5(CLBLL_R_X71Y131_SLICE_X107Y131_DO5),
.O6(CLBLL_R_X71Y131_SLICE_X107Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafafad8505050d8)
  ) CLBLL_R_X71Y131_SLICE_X107Y131_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X72Y134_SLICE_X109Y134_AO5),
.I2(CLBLM_L_X72Y131_SLICE_X108Y131_CQ),
.I3(CLBLM_L_X72Y131_SLICE_X108Y131_DO5),
.I4(CLBLM_L_X72Y133_SLICE_X109Y133_DO6),
.I5(CLBLL_R_X71Y131_SLICE_X107Y131_CQ),
.O5(CLBLL_R_X71Y131_SLICE_X107Y131_CO5),
.O6(CLBLL_R_X71Y131_SLICE_X107Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hddccf0f088ccf0f0)
  ) CLBLL_R_X71Y131_SLICE_X107Y131_BLUT (
.I0(CLBLM_L_X72Y133_SLICE_X109Y133_DO6),
.I1(CLBLL_R_X71Y131_SLICE_X107Y131_BQ),
.I2(CLBLL_R_X71Y131_SLICE_X107Y131_CQ),
.I3(CLBLM_L_X72Y130_SLICE_X108Y130_AO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X72Y134_SLICE_X109Y134_AO5),
.O5(CLBLL_R_X71Y131_SLICE_X107Y131_BO5),
.O6(CLBLL_R_X71Y131_SLICE_X107Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0faccccf050cccc)
  ) CLBLL_R_X71Y131_SLICE_X107Y131_ALUT (
.I0(CLBLM_L_X72Y131_SLICE_X108Y131_A5Q),
.I1(CLBLL_R_X71Y131_SLICE_X107Y131_BQ),
.I2(CLBLL_R_X71Y131_SLICE_X107Y131_AQ),
.I3(CLBLM_L_X72Y131_SLICE_X109Y131_AO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X72Y134_SLICE_X109Y134_AO5),
.O5(CLBLL_R_X71Y131_SLICE_X107Y131_AO5),
.O6(CLBLL_R_X71Y131_SLICE_X107Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y132_SLICE_X106Y132_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y132_SLICE_X106Y132_AO6),
.Q(CLBLL_R_X71Y132_SLICE_X106Y132_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y132_SLICE_X106Y132_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y132_SLICE_X106Y132_BO6),
.Q(CLBLL_R_X71Y132_SLICE_X106Y132_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y132_SLICE_X106Y132_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y132_SLICE_X106Y132_CO6),
.Q(CLBLL_R_X71Y132_SLICE_X106Y132_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y132_SLICE_X106Y132_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y132_SLICE_X106Y132_DO6),
.Q(CLBLL_R_X71Y132_SLICE_X106Y132_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a0f5d7a082)
  ) CLBLL_R_X71Y132_SLICE_X106Y132_DLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X72Y133_SLICE_X108Y133_AQ),
.I2(CLBLL_R_X71Y132_SLICE_X106Y132_DQ),
.I3(CLBLL_R_X73Y132_SLICE_X110Y132_BO6),
.I4(CLBLL_R_X71Y133_SLICE_X106Y133_DQ),
.I5(CLBLM_L_X72Y133_SLICE_X108Y133_A5Q),
.O5(CLBLL_R_X71Y132_SLICE_X106Y132_DO5),
.O6(CLBLL_R_X71Y132_SLICE_X106Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h66ccf0f0ccccf0f0)
  ) CLBLL_R_X71Y132_SLICE_X106Y132_CLUT (
.I0(CLBLL_R_X71Y125_SLICE_X107Y125_CO6),
.I1(CLBLL_R_X71Y132_SLICE_X106Y132_CQ),
.I2(CLBLL_R_X71Y132_SLICE_X106Y132_BQ),
.I3(CLBLL_R_X71Y131_SLICE_X107Y131_A5Q),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X71Y131_SLICE_X106Y131_AQ),
.O5(CLBLL_R_X71Y132_SLICE_X106Y132_CO5),
.O6(CLBLL_R_X71Y132_SLICE_X106Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacacaca5aaa5aaa)
  ) CLBLL_R_X71Y132_SLICE_X106Y132_BLUT (
.I0(CLBLL_R_X71Y132_SLICE_X107Y132_DQ),
.I1(CLBLL_R_X71Y132_SLICE_X106Y132_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X72Y133_SLICE_X109Y133_BQ),
.I4(1'b1),
.I5(CLBLL_R_X71Y132_SLICE_X106Y132_AO5),
.O5(CLBLL_R_X71Y132_SLICE_X106Y132_BO5),
.O6(CLBLL_R_X71Y132_SLICE_X106Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f3c0ff0fffff)
  ) CLBLL_R_X71Y132_SLICE_X106Y132_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLL_R_X71Y132_SLICE_X106Y132_AQ),
.I3(CLBLL_R_X71Y131_SLICE_X106Y131_AQ),
.I4(CLBLL_R_X71Y125_SLICE_X107Y125_CO6),
.I5(1'b1),
.O5(CLBLL_R_X71Y132_SLICE_X106Y132_AO5),
.O6(CLBLL_R_X71Y132_SLICE_X106Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y132_SLICE_X107Y132_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y132_SLICE_X107Y132_AO5),
.Q(CLBLL_R_X71Y132_SLICE_X107Y132_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y132_SLICE_X107Y132_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y132_SLICE_X107Y132_BO6),
.Q(CLBLL_R_X71Y132_SLICE_X107Y132_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y132_SLICE_X107Y132_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y132_SLICE_X107Y132_CO6),
.Q(CLBLL_R_X71Y132_SLICE_X107Y132_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y132_SLICE_X107Y132_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y132_SLICE_X107Y132_DO6),
.Q(CLBLL_R_X71Y132_SLICE_X107Y132_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3ccc9cccf0ccf0cc)
  ) CLBLL_R_X71Y132_SLICE_X107Y132_DLUT (
.I0(CLBLL_R_X71Y132_SLICE_X106Y132_AQ),
.I1(CLBLL_R_X71Y132_SLICE_X107Y132_CQ),
.I2(CLBLL_R_X71Y132_SLICE_X107Y132_DQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLL_R_X71Y131_SLICE_X106Y131_AQ),
.I5(CLBLL_R_X71Y125_SLICE_X107Y125_CO6),
.O5(CLBLL_R_X71Y132_SLICE_X107Y132_DO5),
.O6(CLBLL_R_X71Y132_SLICE_X107Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafa0a0cfcfc0c0)
  ) CLBLL_R_X71Y132_SLICE_X107Y132_CLUT (
.I0(CLBLM_L_X72Y132_SLICE_X109Y132_BO6),
.I1(CLBLL_R_X71Y132_SLICE_X107Y132_CQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(1'b1),
.I4(CLBLL_R_X71Y131_SLICE_X107Y131_A5Q),
.I5(CLBLL_R_X71Y125_SLICE_X107Y125_CO6),
.O5(CLBLL_R_X71Y132_SLICE_X107Y132_CO5),
.O6(CLBLL_R_X71Y132_SLICE_X107Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8cffdcff8c00dc00)
  ) CLBLL_R_X71Y132_SLICE_X107Y132_BLUT (
.I0(CLBLL_R_X71Y131_SLICE_X107Y131_DO6),
.I1(CLBLL_R_X71Y132_SLICE_X107Y132_BQ),
.I2(CLBLL_R_X71Y125_SLICE_X107Y125_CO6),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLL_R_X71Y132_SLICE_X107Y132_AO6),
.I5(CLBLM_L_X72Y132_SLICE_X108Y132_BQ),
.O5(CLBLL_R_X71Y132_SLICE_X107Y132_BO5),
.O6(CLBLL_R_X71Y132_SLICE_X107Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000f0f0f3aac0aa)
  ) CLBLL_R_X71Y132_SLICE_X107Y132_ALUT (
.I0(CLBLM_L_X72Y132_SLICE_X109Y132_AQ),
.I1(CLBLL_R_X73Y132_SLICE_X110Y132_BO6),
.I2(CLBLL_R_X71Y132_SLICE_X107Y132_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X72Y133_SLICE_X108Y133_AQ),
.I5(1'b1),
.O5(CLBLL_R_X71Y132_SLICE_X107Y132_AO5),
.O6(CLBLL_R_X71Y132_SLICE_X107Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y133_SLICE_X106Y133_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y133_SLICE_X106Y133_AO5),
.Q(CLBLL_R_X71Y133_SLICE_X106Y133_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y133_SLICE_X106Y133_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y133_SLICE_X106Y133_BO6),
.Q(CLBLL_R_X71Y133_SLICE_X106Y133_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y133_SLICE_X106Y133_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y133_SLICE_X106Y133_CO6),
.Q(CLBLL_R_X71Y133_SLICE_X106Y133_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y133_SLICE_X106Y133_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y133_SLICE_X106Y133_DO6),
.Q(CLBLL_R_X71Y133_SLICE_X106Y133_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc66e4e4cc66e4e4)
  ) CLBLL_R_X71Y133_SLICE_X106Y133_DLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X71Y133_SLICE_X106Y133_CQ),
.I2(CLBLL_R_X71Y133_SLICE_X106Y133_DQ),
.I3(CLBLL_R_X71Y132_SLICE_X106Y132_CQ),
.I4(CLBLM_L_X72Y133_SLICE_X108Y133_BO5),
.I5(1'b1),
.O5(CLBLL_R_X71Y133_SLICE_X106Y133_DO5),
.O6(CLBLL_R_X71Y133_SLICE_X106Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88dd88df80)
  ) CLBLL_R_X71Y133_SLICE_X106Y133_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X71Y133_SLICE_X106Y133_CQ),
.I2(CLBLM_L_X72Y133_SLICE_X108Y133_A5Q),
.I3(CLBLL_R_X71Y132_SLICE_X106Y132_CQ),
.I4(CLBLM_L_X72Y133_SLICE_X108Y133_AQ),
.I5(CLBLL_R_X73Y132_SLICE_X110Y132_BO6),
.O5(CLBLL_R_X71Y133_SLICE_X106Y133_CO5),
.O6(CLBLL_R_X71Y133_SLICE_X106Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c6cff00ccccff00)
  ) CLBLL_R_X71Y133_SLICE_X106Y133_BLUT (
.I0(CLBLM_L_X70Y124_SLICE_X105Y124_AO6),
.I1(CLBLL_R_X71Y133_SLICE_X106Y133_BQ),
.I2(CLBLM_L_X70Y133_SLICE_X105Y133_AQ),
.I3(CLBLM_L_X70Y133_SLICE_X105Y133_DQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X70Y133_SLICE_X104Y133_AQ),
.O5(CLBLL_R_X71Y133_SLICE_X106Y133_BO5),
.O6(CLBLL_R_X71Y133_SLICE_X106Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h30303030f5dda088)
  ) CLBLL_R_X71Y133_SLICE_X106Y133_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X70Y135_SLICE_X105Y135_AQ),
.I2(CLBLL_R_X71Y133_SLICE_X106Y133_AQ),
.I3(CLBLM_L_X72Y133_SLICE_X109Y133_CO6),
.I4(CLBLM_L_X70Y132_SLICE_X105Y132_AQ),
.I5(1'b1),
.O5(CLBLL_R_X71Y133_SLICE_X106Y133_AO5),
.O6(CLBLL_R_X71Y133_SLICE_X106Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y133_SLICE_X107Y133_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y133_SLICE_X107Y133_AO6),
.Q(CLBLL_R_X71Y133_SLICE_X107Y133_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y133_SLICE_X107Y133_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y133_SLICE_X107Y133_BO6),
.Q(CLBLL_R_X71Y133_SLICE_X107Y133_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y133_SLICE_X107Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y133_SLICE_X107Y133_DO5),
.O6(CLBLL_R_X71Y133_SLICE_X107Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8080808080808080)
  ) CLBLL_R_X71Y133_SLICE_X107Y133_CLUT (
.I0(CLBLM_L_X70Y133_SLICE_X105Y133_AQ),
.I1(CLBLM_L_X70Y133_SLICE_X104Y133_AQ),
.I2(CLBLM_L_X70Y124_SLICE_X105Y124_AO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y133_SLICE_X107Y133_CO5),
.O6(CLBLL_R_X71Y133_SLICE_X107Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ccf00ff0ccf0)
  ) CLBLL_R_X71Y133_SLICE_X107Y133_BLUT (
.I0(1'b1),
.I1(CLBLL_R_X71Y133_SLICE_X107Y133_BQ),
.I2(CLBLL_R_X71Y133_SLICE_X107Y133_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLL_R_X71Y133_SLICE_X107Y133_CO6),
.I5(CLBLL_R_X71Y134_SLICE_X107Y134_CQ),
.O5(CLBLL_R_X71Y133_SLICE_X107Y133_BO5),
.O6(CLBLL_R_X71Y133_SLICE_X107Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8fff0ff7000f000)
  ) CLBLL_R_X71Y133_SLICE_X107Y133_ALUT (
.I0(CLBLM_L_X70Y124_SLICE_X105Y124_AO6),
.I1(CLBLM_L_X70Y133_SLICE_X104Y133_AQ),
.I2(CLBLL_R_X71Y133_SLICE_X107Y133_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X70Y133_SLICE_X105Y133_AQ),
.I5(CLBLL_R_X71Y134_SLICE_X107Y134_CQ),
.O5(CLBLL_R_X71Y133_SLICE_X107Y133_AO5),
.O6(CLBLL_R_X71Y133_SLICE_X107Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y134_SLICE_X106Y134_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y134_SLICE_X106Y134_AO6),
.Q(CLBLL_R_X71Y134_SLICE_X106Y134_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y134_SLICE_X106Y134_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y134_SLICE_X106Y134_BO6),
.Q(CLBLL_R_X71Y134_SLICE_X106Y134_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y134_SLICE_X106Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y134_SLICE_X106Y134_DO5),
.O6(CLBLL_R_X71Y134_SLICE_X106Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y134_SLICE_X106Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y134_SLICE_X106Y134_CO5),
.O6(CLBLL_R_X71Y134_SLICE_X106Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc3ccaaaac7c8aaaa)
  ) CLBLL_R_X71Y134_SLICE_X106Y134_BLUT (
.I0(CLBLM_L_X70Y135_SLICE_X105Y135_A5Q),
.I1(CLBLL_R_X71Y134_SLICE_X106Y134_BQ),
.I2(CLBLM_L_X72Y133_SLICE_X109Y133_CO6),
.I3(CLBLM_L_X72Y134_SLICE_X109Y134_BO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X70Y135_SLICE_X105Y135_AQ),
.O5(CLBLL_R_X71Y134_SLICE_X106Y134_BO5),
.O6(CLBLL_R_X71Y134_SLICE_X106Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000d00)
  ) CLBLL_R_X71Y134_SLICE_X106Y134_ALUT (
.I0(CLBLM_L_X70Y136_SLICE_X105Y136_BO5),
.I1(CLBLL_R_X75Y134_SLICE_X114Y134_CO6),
.I2(CLBLL_R_X71Y134_SLICE_X106Y134_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X60Y92_SLICE_X90Y92_AQ),
.I5(CLBLM_L_X60Y94_SLICE_X90Y94_AQ),
.O5(CLBLL_R_X71Y134_SLICE_X106Y134_AO5),
.O6(CLBLL_R_X71Y134_SLICE_X106Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y134_SLICE_X107Y134_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y134_SLICE_X107Y134_AO6),
.Q(CLBLL_R_X71Y134_SLICE_X107Y134_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y134_SLICE_X107Y134_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y134_SLICE_X107Y134_BO6),
.Q(CLBLL_R_X71Y134_SLICE_X107Y134_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y134_SLICE_X107Y134_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y134_SLICE_X107Y134_CO6),
.Q(CLBLL_R_X71Y134_SLICE_X107Y134_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y134_SLICE_X107Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y134_SLICE_X107Y134_DO5),
.O6(CLBLL_R_X71Y134_SLICE_X107Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccff00c9c9ff00)
  ) CLBLL_R_X71Y134_SLICE_X107Y134_CLUT (
.I0(CLBLM_L_X72Y133_SLICE_X109Y133_CO6),
.I1(CLBLL_R_X71Y134_SLICE_X107Y134_CQ),
.I2(CLBLM_L_X70Y135_SLICE_X105Y135_A5Q),
.I3(CLBLL_R_X71Y134_SLICE_X107Y134_BQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X70Y135_SLICE_X105Y135_AQ),
.O5(CLBLL_R_X71Y134_SLICE_X107Y134_CO5),
.O6(CLBLL_R_X71Y134_SLICE_X107Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf00ff0f0ccccf0f0)
  ) CLBLL_R_X71Y134_SLICE_X107Y134_BLUT (
.I0(1'b1),
.I1(CLBLL_R_X71Y134_SLICE_X107Y134_BQ),
.I2(CLBLL_R_X71Y134_SLICE_X107Y134_AQ),
.I3(CLBLL_R_X71Y133_SLICE_X106Y133_BQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X70Y134_SLICE_X105Y134_DO6),
.O5(CLBLL_R_X71Y134_SLICE_X107Y134_BO5),
.O6(CLBLL_R_X71Y134_SLICE_X107Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0f5a0f780)
  ) CLBLL_R_X71Y134_SLICE_X107Y134_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X70Y135_SLICE_X105Y135_AQ),
.I2(CLBLL_R_X71Y134_SLICE_X107Y134_AQ),
.I3(CLBLL_R_X71Y133_SLICE_X106Y133_BQ),
.I4(CLBLM_L_X72Y133_SLICE_X109Y133_CO6),
.I5(CLBLM_L_X70Y135_SLICE_X105Y135_A5Q),
.O5(CLBLL_R_X71Y134_SLICE_X107Y134_AO5),
.O6(CLBLL_R_X71Y134_SLICE_X107Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y101_SLICE_X110Y101_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y101_SLICE_X110Y101_AO6),
.Q(CLBLL_R_X73Y101_SLICE_X110Y101_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y101_SLICE_X110Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y101_SLICE_X110Y101_DO5),
.O6(CLBLL_R_X73Y101_SLICE_X110Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y101_SLICE_X110Y101_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y101_SLICE_X110Y101_CO5),
.O6(CLBLL_R_X73Y101_SLICE_X110Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y101_SLICE_X110Y101_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y101_SLICE_X110Y101_BO5),
.O6(CLBLL_R_X73Y101_SLICE_X110Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0e2e2ff00ff00)
  ) CLBLL_R_X73Y101_SLICE_X110Y101_ALUT (
.I0(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I1(CLBLM_L_X72Y103_SLICE_X108Y103_CO6),
.I2(CLBLL_R_X73Y101_SLICE_X110Y101_AQ),
.I3(CLBLL_R_X73Y103_SLICE_X110Y103_BQ),
.I4(CLBLM_L_X72Y103_SLICE_X108Y103_DO6),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLL_R_X73Y101_SLICE_X110Y101_AO5),
.O6(CLBLL_R_X73Y101_SLICE_X110Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y101_SLICE_X111Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y101_SLICE_X111Y101_DO5),
.O6(CLBLL_R_X73Y101_SLICE_X111Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y101_SLICE_X111Y101_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y101_SLICE_X111Y101_CO5),
.O6(CLBLL_R_X73Y101_SLICE_X111Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y101_SLICE_X111Y101_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y101_SLICE_X111Y101_BO5),
.O6(CLBLL_R_X73Y101_SLICE_X111Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y101_SLICE_X111Y101_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y101_SLICE_X111Y101_AO5),
.O6(CLBLL_R_X73Y101_SLICE_X111Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y102_SLICE_X110Y102_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y102_SLICE_X111Y102_A5Q),
.Q(CLBLL_R_X73Y102_SLICE_X110Y102_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y102_SLICE_X110Y102_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y102_SLICE_X110Y102_AO6),
.Q(CLBLL_R_X73Y102_SLICE_X110Y102_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y102_SLICE_X110Y102_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y102_SLICE_X110Y102_BO6),
.Q(CLBLL_R_X73Y102_SLICE_X110Y102_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y102_SLICE_X110Y102_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y102_SLICE_X110Y102_CO6),
.Q(CLBLL_R_X73Y102_SLICE_X110Y102_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0ff00ff00ff00ff)
  ) CLBLL_R_X73Y102_SLICE_X110Y102_DLUT (
.I0(1'b1),
.I1(CLBLL_R_X73Y102_SLICE_X111Y102_A5Q),
.I2(CLBLM_L_X72Y104_SLICE_X109Y104_BQ),
.I3(CLBLL_R_X73Y104_SLICE_X110Y104_A5Q),
.I4(CLBLL_R_X73Y102_SLICE_X110Y102_CQ),
.I5(CLBLM_L_X72Y104_SLICE_X109Y104_B5Q),
.O5(CLBLL_R_X73Y102_SLICE_X110Y102_DO5),
.O6(CLBLL_R_X73Y102_SLICE_X110Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88df8add88d580)
  ) CLBLL_R_X73Y102_SLICE_X110Y102_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X73Y102_SLICE_X110Y102_CQ),
.I2(CLBLM_L_X72Y103_SLICE_X108Y103_CO5),
.I3(CLBLL_R_X73Y102_SLICE_X110Y102_BQ),
.I4(CLBLM_L_X72Y103_SLICE_X108Y103_DO5),
.I5(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.O5(CLBLL_R_X73Y102_SLICE_X110Y102_CO5),
.O6(CLBLL_R_X73Y102_SLICE_X110Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcdcdff00c8c8ff00)
  ) CLBLL_R_X73Y102_SLICE_X110Y102_BLUT (
.I0(CLBLM_L_X72Y103_SLICE_X108Y103_CO5),
.I1(CLBLL_R_X73Y102_SLICE_X110Y102_BQ),
.I2(CLBLM_L_X72Y103_SLICE_X108Y103_DO6),
.I3(CLBLM_L_X72Y103_SLICE_X109Y103_BQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.O5(CLBLL_R_X73Y102_SLICE_X110Y102_BO5),
.O6(CLBLL_R_X73Y102_SLICE_X110Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2eee2e2e222e2)
  ) CLBLL_R_X73Y102_SLICE_X110Y102_ALUT (
.I0(CLBLL_R_X73Y102_SLICE_X110Y102_CQ),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLL_R_X73Y102_SLICE_X110Y102_AQ),
.I3(CLBLM_L_X72Y103_SLICE_X108Y103_A5Q),
.I4(CLBLM_L_X72Y103_SLICE_X108Y103_CO5),
.I5(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.O5(CLBLL_R_X73Y102_SLICE_X110Y102_AO5),
.O6(CLBLL_R_X73Y102_SLICE_X110Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y102_SLICE_X111Y102_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y103_SLICE_X110Y103_B5Q),
.Q(CLBLL_R_X73Y102_SLICE_X111Y102_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y102_SLICE_X111Y102_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y102_SLICE_X111Y102_AO6),
.Q(CLBLL_R_X73Y102_SLICE_X111Y102_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0f0f0faf0)
  ) CLBLL_R_X73Y102_SLICE_X111Y102_DLUT (
.I0(CLBLL_R_X73Y103_SLICE_X110Y103_B5Q),
.I1(1'b1),
.I2(CLBLL_R_X73Y104_SLICE_X110Y104_A5Q),
.I3(CLBLM_L_X74Y103_SLICE_X113Y103_BQ),
.I4(CLBLM_L_X72Y104_SLICE_X109Y104_BQ),
.I5(CLBLM_L_X72Y104_SLICE_X109Y104_B5Q),
.O5(CLBLL_R_X73Y102_SLICE_X111Y102_DO5),
.O6(CLBLL_R_X73Y102_SLICE_X111Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafafac8fafafafa)
  ) CLBLL_R_X73Y102_SLICE_X111Y102_CLUT (
.I0(CLBLM_L_X72Y103_SLICE_X109Y103_DO6),
.I1(CLBLM_L_X74Y103_SLICE_X112Y103_DO6),
.I2(CLBLL_R_X73Y102_SLICE_X110Y102_DO6),
.I3(CLBLM_L_X74Y103_SLICE_X112Y103_CO6),
.I4(CLBLL_R_X73Y102_SLICE_X111Y102_DO6),
.I5(CLBLL_R_X73Y102_SLICE_X111Y102_BO6),
.O5(CLBLL_R_X73Y102_SLICE_X111Y102_CO5),
.O6(CLBLL_R_X73Y102_SLICE_X111Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'habffafffbbffffff)
  ) CLBLL_R_X73Y102_SLICE_X111Y102_BLUT (
.I0(CLBLM_L_X72Y104_SLICE_X109Y104_BQ),
.I1(CLBLL_R_X73Y103_SLICE_X111Y103_AQ),
.I2(CLBLL_R_X73Y102_SLICE_X111Y102_AQ),
.I3(CLBLM_L_X72Y104_SLICE_X109Y104_B5Q),
.I4(CLBLL_R_X73Y102_SLICE_X111Y102_A5Q),
.I5(CLBLM_L_X60Y101_SLICE_X90Y101_AQ),
.O5(CLBLL_R_X73Y102_SLICE_X111Y102_BO5),
.O6(CLBLL_R_X73Y102_SLICE_X111Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0fda8f5a07520)
  ) CLBLL_R_X73Y102_SLICE_X111Y102_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X72Y103_SLICE_X108Y103_A5Q),
.I2(CLBLL_R_X73Y102_SLICE_X111Y102_AQ),
.I3(CLBLM_L_X74Y102_SLICE_X112Y102_AQ),
.I4(CLBLM_L_X72Y103_SLICE_X108Y103_CO6),
.I5(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.O5(CLBLL_R_X73Y102_SLICE_X111Y102_AO5),
.O6(CLBLL_R_X73Y102_SLICE_X111Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y103_SLICE_X110Y103_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X60Y101_SLICE_X90Y101_AQ),
.Q(CLBLL_R_X73Y103_SLICE_X110Y103_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y103_SLICE_X110Y103_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y103_SLICE_X109Y103_AQ),
.Q(CLBLL_R_X73Y103_SLICE_X110Y103_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y103_SLICE_X110Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y103_SLICE_X110Y103_AO6),
.Q(CLBLL_R_X73Y103_SLICE_X110Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y103_SLICE_X110Y103_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y103_SLICE_X110Y103_BO6),
.Q(CLBLL_R_X73Y103_SLICE_X110Y103_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff8fff0fff0fff0)
  ) CLBLL_R_X73Y103_SLICE_X110Y103_DLUT (
.I0(CLBLL_R_X73Y102_SLICE_X110Y102_AQ),
.I1(CLBLL_R_X73Y104_SLICE_X110Y104_A5Q),
.I2(CLBLL_R_X73Y103_SLICE_X111Y103_DO6),
.I3(CLBLL_R_X73Y103_SLICE_X110Y103_CO6),
.I4(CLBLM_L_X72Y103_SLICE_X109Y103_AO5),
.I5(CLBLL_R_X73Y102_SLICE_X110Y102_A5Q),
.O5(CLBLL_R_X73Y103_SLICE_X110Y103_DO5),
.O6(CLBLL_R_X73Y103_SLICE_X110Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h400000000ff00ff0)
  ) CLBLL_R_X73Y103_SLICE_X110Y103_CLUT (
.I0(CLBLM_L_X72Y104_SLICE_X109Y104_BQ),
.I1(CLBLL_R_X73Y103_SLICE_X110Y103_AQ),
.I2(CLBLL_R_X75Y103_SLICE_X115Y103_AQ),
.I3(CLBLL_R_X73Y104_SLICE_X110Y104_A5Q),
.I4(CLBLM_L_X72Y104_SLICE_X109Y104_B5Q),
.I5(1'b1),
.O5(CLBLL_R_X73Y103_SLICE_X110Y103_CO5),
.O6(CLBLL_R_X73Y103_SLICE_X110Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccaaf0f0f0f0)
  ) CLBLL_R_X73Y103_SLICE_X110Y103_BLUT (
.I0(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I1(CLBLL_R_X73Y103_SLICE_X110Y103_BQ),
.I2(CLBLL_R_X73Y103_SLICE_X110Y103_AQ),
.I3(CLBLM_L_X72Y103_SLICE_X108Y103_BO5),
.I4(CLBLM_L_X72Y103_SLICE_X108Y103_CO6),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLL_R_X73Y103_SLICE_X110Y103_BO5),
.O6(CLBLL_R_X73Y103_SLICE_X110Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1e0f1e0ffff0000)
  ) CLBLL_R_X73Y103_SLICE_X110Y103_ALUT (
.I0(CLBLM_L_X72Y103_SLICE_X108Y103_BO6),
.I1(CLBLM_L_X72Y103_SLICE_X108Y103_CO6),
.I2(CLBLL_R_X73Y103_SLICE_X110Y103_AQ),
.I3(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I4(CLBLL_R_X73Y102_SLICE_X110Y102_AQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLL_R_X73Y103_SLICE_X110Y103_AO5),
.O6(CLBLL_R_X73Y103_SLICE_X110Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y103_SLICE_X111Y103_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X79Y104_SLICE_X122Y104_A5Q),
.Q(CLBLL_R_X73Y103_SLICE_X111Y103_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y103_SLICE_X111Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y103_SLICE_X111Y103_AO6),
.Q(CLBLL_R_X73Y103_SLICE_X111Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8080000000000000)
  ) CLBLL_R_X73Y103_SLICE_X111Y103_DLUT (
.I0(CLBLM_L_X60Y101_SLICE_X90Y101_AQ),
.I1(CLBLL_R_X73Y104_SLICE_X110Y104_A5Q),
.I2(CLBLM_L_X72Y104_SLICE_X109Y104_BQ),
.I3(1'b1),
.I4(CLBLM_L_X72Y104_SLICE_X109Y104_B5Q),
.I5(CLBLL_R_X73Y104_SLICE_X111Y104_BQ),
.O5(CLBLL_R_X73Y103_SLICE_X111Y103_DO5),
.O6(CLBLL_R_X73Y103_SLICE_X111Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfdfdddfdfdfdfdf)
  ) CLBLL_R_X73Y103_SLICE_X111Y103_CLUT (
.I0(CLBLM_L_X72Y104_SLICE_X109Y104_BQ),
.I1(CLBLM_L_X72Y104_SLICE_X109Y104_B5Q),
.I2(CLBLL_R_X73Y104_SLICE_X111Y104_CO6),
.I3(CLBLL_R_X79Y104_SLICE_X122Y104_A5Q),
.I4(CLBLL_R_X73Y103_SLICE_X110Y103_CO5),
.I5(CLBLL_R_X73Y103_SLICE_X110Y103_BQ),
.O5(CLBLL_R_X73Y103_SLICE_X111Y103_CO5),
.O6(CLBLL_R_X73Y103_SLICE_X111Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0c0e0f0f0f0f0)
  ) CLBLL_R_X73Y103_SLICE_X111Y103_BLUT (
.I0(CLBLM_L_X74Y103_SLICE_X113Y103_DO6),
.I1(CLBLL_R_X73Y103_SLICE_X110Y103_DO6),
.I2(CLBLM_L_X70Y105_SLICE_X104Y105_BO6),
.I3(CLBLL_R_X75Y103_SLICE_X114Y103_BO6),
.I4(CLBLL_R_X73Y102_SLICE_X111Y102_CO6),
.I5(CLBLL_R_X73Y103_SLICE_X111Y103_CO6),
.O5(CLBLL_R_X73Y103_SLICE_X111Y103_BO5),
.O6(CLBLL_R_X73Y103_SLICE_X111Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f7b3c0c0c480)
  ) CLBLL_R_X73Y103_SLICE_X111Y103_ALUT (
.I0(CLBLL_R_X73Y104_SLICE_X110Y104_DO6),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLL_R_X73Y103_SLICE_X111Y103_AQ),
.I3(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I4(CLBLM_L_X72Y103_SLICE_X108Y103_DO5),
.I5(CLBLM_L_X74Y103_SLICE_X113Y103_BQ),
.O5(CLBLL_R_X73Y103_SLICE_X111Y103_AO5),
.O6(CLBLL_R_X73Y103_SLICE_X111Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y104_SLICE_X110Y104_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y104_SLICE_X110Y104_AO5),
.Q(CLBLL_R_X73Y104_SLICE_X110Y104_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y104_SLICE_X110Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y104_SLICE_X110Y104_AO6),
.Q(CLBLL_R_X73Y104_SLICE_X110Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y104_SLICE_X110Y104_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y104_SLICE_X110Y104_BO6),
.Q(CLBLL_R_X73Y104_SLICE_X110Y104_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y104_SLICE_X110Y104_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y104_SLICE_X110Y104_CO6),
.Q(CLBLL_R_X73Y104_SLICE_X110Y104_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff0ff0fff0fff)
  ) CLBLL_R_X73Y104_SLICE_X110Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X72Y104_SLICE_X109Y104_A5Q),
.I3(CLBLL_R_X73Y104_SLICE_X110Y104_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y104_SLICE_X110Y104_DO5),
.O6(CLBLL_R_X73Y104_SLICE_X110Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccaf0f0f0f0)
  ) CLBLL_R_X73Y104_SLICE_X110Y104_CLUT (
.I0(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I1(CLBLL_R_X73Y104_SLICE_X110Y104_CQ),
.I2(CLBLL_R_X73Y104_SLICE_X110Y104_BQ),
.I3(CLBLM_L_X72Y103_SLICE_X108Y103_BO6),
.I4(CLBLM_L_X72Y104_SLICE_X109Y104_A5Q),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLL_R_X73Y104_SLICE_X110Y104_CO5),
.O6(CLBLL_R_X73Y104_SLICE_X110Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6aca6aca88008800)
  ) CLBLL_R_X73Y104_SLICE_X110Y104_BLUT (
.I0(CLBLM_L_X72Y104_SLICE_X109Y104_A5Q),
.I1(CLBLL_R_X73Y104_SLICE_X110Y104_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X72Y103_SLICE_X108Y103_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y104_SLICE_X110Y104_BO5),
.O6(CLBLL_R_X73Y104_SLICE_X110Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa50507722dd88)
  ) CLBLL_R_X73Y104_SLICE_X110Y104_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X73Y104_SLICE_X111Y104_DO6),
.I2(CLBLL_R_X73Y111_SLICE_X110Y111_AQ),
.I3(CLBLL_R_X73Y102_SLICE_X110Y102_A5Q),
.I4(CLBLL_R_X73Y104_SLICE_X110Y104_A5Q),
.I5(1'b1),
.O5(CLBLL_R_X73Y104_SLICE_X110Y104_AO5),
.O6(CLBLL_R_X73Y104_SLICE_X110Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y104_SLICE_X111Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y104_SLICE_X111Y104_AO6),
.Q(CLBLL_R_X73Y104_SLICE_X111Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y104_SLICE_X111Y104_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y104_SLICE_X111Y104_BO6),
.Q(CLBLL_R_X73Y104_SLICE_X111Y104_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc000c00000000000)
  ) CLBLL_R_X73Y104_SLICE_X111Y104_DLUT (
.I0(1'b1),
.I1(CLBLL_R_X79Y104_SLICE_X122Y104_A5Q),
.I2(CLBLM_L_X62Y95_SLICE_X92Y95_AQ),
.I3(CLBLL_R_X73Y103_SLICE_X111Y103_A5Q),
.I4(1'b1),
.I5(CLBLL_R_X75Y103_SLICE_X115Y103_AQ),
.O5(CLBLL_R_X73Y104_SLICE_X111Y104_DO5),
.O6(CLBLL_R_X73Y104_SLICE_X111Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8883000c888c000)
  ) CLBLL_R_X73Y104_SLICE_X111Y104_CLUT (
.I0(CLBLL_R_X73Y102_SLICE_X110Y102_BQ),
.I1(CLBLL_R_X73Y104_SLICE_X110Y104_A5Q),
.I2(CLBLM_L_X62Y95_SLICE_X92Y95_AQ),
.I3(CLBLL_R_X73Y104_SLICE_X111Y104_AQ),
.I4(CLBLL_R_X73Y103_SLICE_X110Y103_B5Q),
.I5(CLBLL_R_X75Y103_SLICE_X115Y103_AQ),
.O5(CLBLL_R_X73Y104_SLICE_X111Y104_CO5),
.O6(CLBLL_R_X73Y104_SLICE_X111Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccaaaaf0ccaaaa)
  ) CLBLL_R_X73Y104_SLICE_X111Y104_BLUT (
.I0(CLBLL_R_X73Y104_SLICE_X111Y104_AQ),
.I1(CLBLL_R_X73Y104_SLICE_X111Y104_BQ),
.I2(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I3(CLBLL_R_X73Y104_SLICE_X110Y104_BO5),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLL_R_X73Y104_SLICE_X111Y104_BO5),
.O6(CLBLL_R_X73Y104_SLICE_X111Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaafcaa00aa30aa)
  ) CLBLL_R_X73Y104_SLICE_X111Y104_ALUT (
.I0(CLBLM_L_X74Y104_SLICE_X112Y104_CQ),
.I1(CLBLL_R_X73Y104_SLICE_X110Y104_DO5),
.I2(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X72Y103_SLICE_X108Y103_DO5),
.I5(CLBLL_R_X73Y104_SLICE_X111Y104_AQ),
.O5(CLBLL_R_X73Y104_SLICE_X111Y104_AO5),
.O6(CLBLL_R_X73Y104_SLICE_X111Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y106_SLICE_X110Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y106_SLICE_X110Y106_DO5),
.O6(CLBLL_R_X73Y106_SLICE_X110Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y106_SLICE_X110Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y106_SLICE_X110Y106_CO5),
.O6(CLBLL_R_X73Y106_SLICE_X110Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555000051550000)
  ) CLBLL_R_X73Y106_SLICE_X110Y106_BLUT (
.I0(CLBLL_R_X73Y108_SLICE_X110Y108_A5Q),
.I1(CLBLM_L_X72Y107_SLICE_X108Y107_A5Q),
.I2(CLBLL_R_X71Y107_SLICE_X106Y107_C5Q),
.I3(CLBLM_L_X74Y107_SLICE_X112Y107_CQ),
.I4(CLBLL_R_X73Y106_SLICE_X110Y106_AO6),
.I5(CLBLL_R_X71Y107_SLICE_X106Y107_CQ),
.O5(CLBLL_R_X73Y106_SLICE_X110Y106_BO5),
.O6(CLBLL_R_X73Y106_SLICE_X110Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff153fffff)
  ) CLBLL_R_X73Y106_SLICE_X110Y106_ALUT (
.I0(CLBLM_L_X74Y107_SLICE_X113Y107_AQ),
.I1(CLBLL_R_X73Y107_SLICE_X111Y107_BQ),
.I2(CLBLM_L_X62Y92_SLICE_X92Y92_AQ),
.I3(CLBLM_L_X72Y107_SLICE_X108Y107_BQ),
.I4(CLBLL_R_X71Y107_SLICE_X106Y107_C5Q),
.I5(CLBLL_R_X71Y107_SLICE_X106Y107_CQ),
.O5(CLBLL_R_X73Y106_SLICE_X110Y106_AO5),
.O6(CLBLL_R_X73Y106_SLICE_X110Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y106_SLICE_X111Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y106_SLICE_X111Y106_DO5),
.O6(CLBLL_R_X73Y106_SLICE_X111Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y106_SLICE_X111Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y106_SLICE_X111Y106_CO5),
.O6(CLBLL_R_X73Y106_SLICE_X111Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y106_SLICE_X111Y106_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y106_SLICE_X111Y106_BO5),
.O6(CLBLL_R_X73Y106_SLICE_X111Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y106_SLICE_X111Y106_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y106_SLICE_X111Y106_AO5),
.O6(CLBLL_R_X73Y106_SLICE_X111Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y107_SLICE_X110Y107_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y107_SLICE_X110Y107_AO6),
.Q(CLBLL_R_X73Y107_SLICE_X110Y107_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y107_SLICE_X110Y107_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y107_SLICE_X110Y107_BO6),
.Q(CLBLL_R_X73Y107_SLICE_X110Y107_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffecffa0ff00ff00)
  ) CLBLL_R_X73Y107_SLICE_X110Y107_DLUT (
.I0(CLBLM_L_X72Y106_SLICE_X108Y106_AQ),
.I1(CLBLM_L_X72Y107_SLICE_X109Y107_BQ),
.I2(CLBLM_L_X74Y107_SLICE_X112Y107_AQ),
.I3(CLBLL_R_X73Y107_SLICE_X110Y107_CO6),
.I4(CLBLL_R_X73Y107_SLICE_X111Y107_DQ),
.I5(CLBLM_L_X72Y107_SLICE_X109Y107_BO5),
.O5(CLBLL_R_X73Y107_SLICE_X110Y107_DO5),
.O6(CLBLL_R_X73Y107_SLICE_X110Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000cc808080)
  ) CLBLL_R_X73Y107_SLICE_X110Y107_CLUT (
.I0(CLBLL_R_X73Y107_SLICE_X111Y107_AQ),
.I1(CLBLL_R_X71Y107_SLICE_X106Y107_CQ),
.I2(CLBLM_L_X72Y107_SLICE_X109Y107_A5Q),
.I3(CLBLL_R_X73Y107_SLICE_X111Y107_CQ),
.I4(CLBLM_L_X72Y107_SLICE_X108Y107_CQ),
.I5(CLBLL_R_X71Y107_SLICE_X106Y107_C5Q),
.O5(CLBLL_R_X73Y107_SLICE_X110Y107_CO5),
.O6(CLBLL_R_X73Y107_SLICE_X110Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffd8ffcc00d800)
  ) CLBLL_R_X73Y107_SLICE_X110Y107_BLUT (
.I0(CLBLM_L_X72Y109_SLICE_X108Y109_BO6),
.I1(CLBLL_R_X73Y107_SLICE_X110Y107_BQ),
.I2(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X72Y108_SLICE_X109Y108_BO6),
.I5(CLBLM_L_X74Y107_SLICE_X112Y107_AQ),
.O5(CLBLL_R_X73Y107_SLICE_X110Y107_BO5),
.O6(CLBLL_R_X73Y107_SLICE_X110Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0ccaaaaaaaa)
  ) CLBLL_R_X73Y107_SLICE_X110Y107_ALUT (
.I0(CLBLM_L_X72Y107_SLICE_X109Y107_AQ),
.I1(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I2(CLBLL_R_X73Y107_SLICE_X110Y107_AQ),
.I3(CLBLM_L_X72Y108_SLICE_X108Y108_BO6),
.I4(CLBLM_L_X72Y108_SLICE_X109Y108_BO6),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLL_R_X73Y107_SLICE_X110Y107_AO5),
.O6(CLBLL_R_X73Y107_SLICE_X110Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y107_SLICE_X111Y107_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y107_SLICE_X111Y107_AO6),
.Q(CLBLL_R_X73Y107_SLICE_X111Y107_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y107_SLICE_X111Y107_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y107_SLICE_X111Y107_BO6),
.Q(CLBLL_R_X73Y107_SLICE_X111Y107_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y107_SLICE_X111Y107_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y107_SLICE_X111Y107_CO6),
.Q(CLBLL_R_X73Y107_SLICE_X111Y107_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y107_SLICE_X111Y107_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y107_SLICE_X111Y107_DO6),
.Q(CLBLL_R_X73Y107_SLICE_X111Y107_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf5ccf0cca0cc)
  ) CLBLL_R_X73Y107_SLICE_X111Y107_DLUT (
.I0(CLBLM_L_X72Y108_SLICE_X109Y108_BO6),
.I1(CLBLL_R_X73Y107_SLICE_X111Y107_AQ),
.I2(CLBLL_R_X73Y107_SLICE_X111Y107_DQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X72Y108_SLICE_X108Y108_BO5),
.I5(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.O5(CLBLL_R_X73Y107_SLICE_X111Y107_DO5),
.O6(CLBLL_R_X73Y107_SLICE_X111Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaaccf0f0f0f0)
  ) CLBLL_R_X73Y107_SLICE_X111Y107_CLUT (
.I0(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I1(CLBLL_R_X73Y107_SLICE_X111Y107_CQ),
.I2(CLBLM_L_X74Y107_SLICE_X113Y107_AQ),
.I3(CLBLM_L_X72Y108_SLICE_X109Y108_A5Q),
.I4(CLBLM_L_X72Y108_SLICE_X108Y108_BO5),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLL_R_X73Y107_SLICE_X111Y107_CO5),
.O6(CLBLL_R_X73Y107_SLICE_X111Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcafaca0acacacaca)
  ) CLBLL_R_X73Y107_SLICE_X111Y107_BLUT (
.I0(CLBLM_L_X74Y107_SLICE_X112Y107_DQ),
.I1(CLBLL_R_X73Y107_SLICE_X111Y107_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X72Y108_SLICE_X108Y108_BO6),
.I4(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I5(CLBLM_L_X72Y108_SLICE_X109Y108_A5Q),
.O5(CLBLL_R_X73Y107_SLICE_X111Y107_BO5),
.O6(CLBLL_R_X73Y107_SLICE_X111Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff05fa00cccccccc)
  ) CLBLL_R_X73Y107_SLICE_X111Y107_ALUT (
.I0(CLBLM_L_X72Y108_SLICE_X108Y108_BO5),
.I1(CLBLL_R_X73Y107_SLICE_X111Y107_BQ),
.I2(CLBLM_L_X72Y108_SLICE_X109Y108_CO5),
.I3(CLBLL_R_X73Y107_SLICE_X111Y107_AQ),
.I4(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLL_R_X73Y107_SLICE_X111Y107_AO5),
.O6(CLBLL_R_X73Y107_SLICE_X111Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y108_SLICE_X110Y108_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y108_SLICE_X110Y108_AO5),
.Q(CLBLL_R_X73Y108_SLICE_X110Y108_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y108_SLICE_X110Y108_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y108_SLICE_X110Y108_AO6),
.Q(CLBLL_R_X73Y108_SLICE_X110Y108_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y108_SLICE_X110Y108_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y108_SLICE_X110Y108_BO6),
.Q(CLBLL_R_X73Y108_SLICE_X110Y108_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y108_SLICE_X110Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y108_SLICE_X110Y108_DO5),
.O6(CLBLL_R_X73Y108_SLICE_X110Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y108_SLICE_X110Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y108_SLICE_X110Y108_CO5),
.O6(CLBLL_R_X73Y108_SLICE_X110Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcdffcd00c8ffc800)
  ) CLBLL_R_X73Y108_SLICE_X110Y108_BLUT (
.I0(CLBLM_L_X72Y109_SLICE_X108Y109_BO6),
.I1(CLBLL_R_X73Y108_SLICE_X110Y108_BQ),
.I2(CLBLM_L_X72Y108_SLICE_X109Y108_BO5),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLL_R_X73Y107_SLICE_X110Y107_BQ),
.I5(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.O5(CLBLL_R_X73Y108_SLICE_X110Y108_BO5),
.O6(CLBLL_R_X73Y108_SLICE_X110Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccf066ff6600)
  ) CLBLL_R_X73Y108_SLICE_X110Y108_ALUT (
.I0(CLBLM_L_X72Y107_SLICE_X109Y107_DO6),
.I1(CLBLL_R_X73Y108_SLICE_X110Y108_A5Q),
.I2(CLBLL_R_X73Y113_SLICE_X110Y113_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X72Y107_SLICE_X108Y107_CQ),
.I5(1'b1),
.O5(CLBLL_R_X73Y108_SLICE_X110Y108_AO5),
.O6(CLBLL_R_X73Y108_SLICE_X110Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y108_SLICE_X111Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y108_SLICE_X111Y108_DO5),
.O6(CLBLL_R_X73Y108_SLICE_X111Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y108_SLICE_X111Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y108_SLICE_X111Y108_CO5),
.O6(CLBLL_R_X73Y108_SLICE_X111Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y108_SLICE_X111Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y108_SLICE_X111Y108_BO5),
.O6(CLBLL_R_X73Y108_SLICE_X111Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y108_SLICE_X111Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y108_SLICE_X111Y108_AO5),
.O6(CLBLL_R_X73Y108_SLICE_X111Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y109_SLICE_X110Y109_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y109_SLICE_X110Y109_AO6),
.Q(CLBLL_R_X73Y109_SLICE_X110Y109_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y109_SLICE_X110Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y109_SLICE_X110Y109_DO5),
.O6(CLBLL_R_X73Y109_SLICE_X110Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y109_SLICE_X110Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y109_SLICE_X110Y109_CO5),
.O6(CLBLL_R_X73Y109_SLICE_X110Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y109_SLICE_X110Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y109_SLICE_X110Y109_BO5),
.O6(CLBLL_R_X73Y109_SLICE_X110Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8f0ff00f0f0ff00)
  ) CLBLL_R_X73Y109_SLICE_X110Y109_ALUT (
.I0(CLBLM_L_X72Y109_SLICE_X109Y109_A5Q),
.I1(CLBLM_L_X72Y109_SLICE_X108Y109_AQ),
.I2(CLBLM_L_X72Y116_SLICE_X108Y116_AQ),
.I3(CLBLM_L_X72Y109_SLICE_X109Y109_C5Q),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X72Y109_SLICE_X109Y109_B5Q),
.O5(CLBLL_R_X73Y109_SLICE_X110Y109_AO5),
.O6(CLBLL_R_X73Y109_SLICE_X110Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y109_SLICE_X111Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y109_SLICE_X111Y109_DO5),
.O6(CLBLL_R_X73Y109_SLICE_X111Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y109_SLICE_X111Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y109_SLICE_X111Y109_CO5),
.O6(CLBLL_R_X73Y109_SLICE_X111Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y109_SLICE_X111Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y109_SLICE_X111Y109_BO5),
.O6(CLBLL_R_X73Y109_SLICE_X111Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y109_SLICE_X111Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y109_SLICE_X111Y109_AO5),
.O6(CLBLL_R_X73Y109_SLICE_X111Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y111_SLICE_X110Y111_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y118_SLICE_X109Y118_A5Q),
.Q(CLBLL_R_X73Y111_SLICE_X110Y111_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y111_SLICE_X110Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y111_SLICE_X110Y111_AO6),
.Q(CLBLL_R_X73Y111_SLICE_X110Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y111_SLICE_X110Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y111_SLICE_X110Y111_DO5),
.O6(CLBLL_R_X73Y111_SLICE_X110Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y111_SLICE_X110Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y111_SLICE_X110Y111_CO5),
.O6(CLBLL_R_X73Y111_SLICE_X110Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y111_SLICE_X110Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y111_SLICE_X110Y111_BO5),
.O6(CLBLL_R_X73Y111_SLICE_X110Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3030ffff33300000)
  ) CLBLL_R_X73Y111_SLICE_X110Y111_ALUT (
.I0(1'b1),
.I1(CLBLL_R_X73Y104_SLICE_X110Y104_AQ),
.I2(CLBLL_R_X73Y111_SLICE_X110Y111_AQ),
.I3(CLBLM_L_X72Y118_SLICE_X109Y118_A5Q),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X73Y111_SLICE_X110Y111_A5Q),
.O5(CLBLL_R_X73Y111_SLICE_X110Y111_AO5),
.O6(CLBLL_R_X73Y111_SLICE_X110Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y111_SLICE_X111Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y111_SLICE_X111Y111_DO5),
.O6(CLBLL_R_X73Y111_SLICE_X111Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y111_SLICE_X111Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y111_SLICE_X111Y111_CO5),
.O6(CLBLL_R_X73Y111_SLICE_X111Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y111_SLICE_X111Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y111_SLICE_X111Y111_BO5),
.O6(CLBLL_R_X73Y111_SLICE_X111Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y111_SLICE_X111Y111_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y111_SLICE_X111Y111_AO5),
.O6(CLBLL_R_X73Y111_SLICE_X111Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y113_SLICE_X110Y113_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y117_SLICE_X106Y117_A5Q),
.Q(CLBLL_R_X73Y113_SLICE_X110Y113_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y113_SLICE_X110Y113_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y113_SLICE_X110Y113_AO6),
.Q(CLBLL_R_X73Y113_SLICE_X110Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y113_SLICE_X110Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y113_SLICE_X110Y113_DO5),
.O6(CLBLL_R_X73Y113_SLICE_X110Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y113_SLICE_X110Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y113_SLICE_X110Y113_CO5),
.O6(CLBLL_R_X73Y113_SLICE_X110Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y113_SLICE_X110Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y113_SLICE_X110Y113_BO5),
.O6(CLBLL_R_X73Y113_SLICE_X110Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3030ffff33300000)
  ) CLBLL_R_X73Y113_SLICE_X110Y113_ALUT (
.I0(1'b1),
.I1(CLBLL_R_X73Y108_SLICE_X110Y108_AQ),
.I2(CLBLL_R_X73Y113_SLICE_X110Y113_AQ),
.I3(CLBLL_R_X71Y117_SLICE_X106Y117_A5Q),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X73Y113_SLICE_X110Y113_A5Q),
.O5(CLBLL_R_X73Y113_SLICE_X110Y113_AO5),
.O6(CLBLL_R_X73Y113_SLICE_X110Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y113_SLICE_X111Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y113_SLICE_X111Y113_DO5),
.O6(CLBLL_R_X73Y113_SLICE_X111Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y113_SLICE_X111Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y113_SLICE_X111Y113_CO5),
.O6(CLBLL_R_X73Y113_SLICE_X111Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y113_SLICE_X111Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y113_SLICE_X111Y113_BO5),
.O6(CLBLL_R_X73Y113_SLICE_X111Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y113_SLICE_X111Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y113_SLICE_X111Y113_AO5),
.O6(CLBLL_R_X73Y113_SLICE_X111Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y118_SLICE_X110Y118_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y118_SLICE_X110Y118_BO5),
.Q(CLBLL_R_X73Y118_SLICE_X110Y118_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y118_SLICE_X110Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y118_SLICE_X110Y118_AO6),
.Q(CLBLL_R_X73Y118_SLICE_X110Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y118_SLICE_X110Y118_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y118_SLICE_X110Y118_BO6),
.Q(CLBLL_R_X73Y118_SLICE_X110Y118_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y118_SLICE_X110Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y118_SLICE_X110Y118_DO5),
.O6(CLBLL_R_X73Y118_SLICE_X110Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y118_SLICE_X110Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y118_SLICE_X110Y118_CO5),
.O6(CLBLL_R_X73Y118_SLICE_X110Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff4022222222)
  ) CLBLL_R_X73Y118_SLICE_X110Y118_BLUT (
.I0(CLBLL_R_X73Y118_SLICE_X111Y118_A5Q),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLL_R_X73Y118_SLICE_X110Y118_AQ),
.I3(CLBLL_R_X73Y119_SLICE_X111Y119_AQ),
.I4(CLBLL_R_X73Y119_SLICE_X110Y119_CO6),
.I5(1'b1),
.O5(CLBLL_R_X73Y118_SLICE_X110Y118_BO5),
.O6(CLBLL_R_X73Y118_SLICE_X110Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccffcc08cc08cc)
  ) CLBLL_R_X73Y118_SLICE_X110Y118_ALUT (
.I0(CLBLL_R_X73Y118_SLICE_X111Y118_A5Q),
.I1(CLBLL_R_X73Y118_SLICE_X110Y118_BQ),
.I2(CLBLL_R_X73Y119_SLICE_X110Y119_CO6),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(1'b1),
.I5(CLBLL_R_X73Y119_SLICE_X110Y119_A5Q),
.O5(CLBLL_R_X73Y118_SLICE_X110Y118_AO5),
.O6(CLBLL_R_X73Y118_SLICE_X110Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y118_SLICE_X111Y118_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y118_SLICE_X111Y118_AO5),
.Q(CLBLL_R_X73Y118_SLICE_X111Y118_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y118_SLICE_X111Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y118_SLICE_X111Y118_AO6),
.Q(CLBLL_R_X73Y118_SLICE_X111Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y118_SLICE_X111Y118_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y118_SLICE_X110Y118_B5Q),
.Q(CLBLL_R_X73Y118_SLICE_X111Y118_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y118_SLICE_X111Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y118_SLICE_X111Y118_DO5),
.O6(CLBLL_R_X73Y118_SLICE_X111Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y118_SLICE_X111Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y118_SLICE_X111Y118_CO5),
.O6(CLBLL_R_X73Y118_SLICE_X111Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y118_SLICE_X111Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y118_SLICE_X111Y118_BO5),
.O6(CLBLL_R_X73Y118_SLICE_X111Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0cc05ccf0aa05aa)
  ) CLBLL_R_X73Y118_SLICE_X111Y118_ALUT (
.I0(CLBLL_R_X73Y119_SLICE_X110Y119_B5Q),
.I1(CLBLL_R_X73Y118_SLICE_X111Y118_BQ),
.I2(CLBLL_R_X73Y119_SLICE_X110Y119_CO6),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLL_R_X73Y118_SLICE_X111Y118_A5Q),
.I5(1'b1),
.O5(CLBLL_R_X73Y118_SLICE_X111Y118_AO5),
.O6(CLBLL_R_X73Y118_SLICE_X111Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y119_SLICE_X110Y119_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y119_SLICE_X110Y119_BQ),
.Q(CLBLL_R_X73Y119_SLICE_X110Y119_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y119_SLICE_X110Y119_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y119_SLICE_X110Y119_BO5),
.Q(CLBLL_R_X73Y119_SLICE_X110Y119_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y119_SLICE_X110Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y119_SLICE_X110Y119_AO6),
.Q(CLBLL_R_X73Y119_SLICE_X110Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y119_SLICE_X110Y119_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y119_SLICE_X110Y119_BO6),
.Q(CLBLL_R_X73Y119_SLICE_X110Y119_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y119_SLICE_X110Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y119_SLICE_X110Y119_DO5),
.O6(CLBLL_R_X73Y119_SLICE_X110Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffefffe)
  ) CLBLL_R_X73Y119_SLICE_X110Y119_CLUT (
.I0(CLBLL_R_X73Y119_SLICE_X111Y119_AQ),
.I1(CLBLL_R_X73Y119_SLICE_X110Y119_AQ),
.I2(CLBLL_R_X73Y119_SLICE_X110Y119_BQ),
.I3(CLBLL_R_X73Y119_SLICE_X110Y119_A5Q),
.I4(1'b1),
.I5(CLBLM_L_X72Y113_SLICE_X108Y113_AQ),
.O5(CLBLL_R_X73Y119_SLICE_X110Y119_CO5),
.O6(CLBLL_R_X73Y119_SLICE_X110Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa22eae233003300)
  ) CLBLL_R_X73Y119_SLICE_X110Y119_BLUT (
.I0(CLBLM_L_X72Y113_SLICE_X108Y113_AQ),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLL_R_X73Y118_SLICE_X111Y118_A5Q),
.I3(CLBLM_L_X72Y119_SLICE_X109Y119_AQ),
.I4(CLBLL_R_X73Y119_SLICE_X110Y119_CO6),
.I5(1'b1),
.O5(CLBLL_R_X73Y119_SLICE_X110Y119_BO5),
.O6(CLBLL_R_X73Y119_SLICE_X110Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h44ee4eee44444e4e)
  ) CLBLL_R_X73Y119_SLICE_X110Y119_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X73Y119_SLICE_X110Y119_A5Q),
.I2(CLBLL_R_X73Y118_SLICE_X111Y118_A5Q),
.I3(CLBLM_L_X72Y119_SLICE_X109Y119_AQ),
.I4(CLBLL_R_X73Y119_SLICE_X110Y119_CO6),
.I5(CLBLM_L_X72Y113_SLICE_X108Y113_AQ),
.O5(CLBLL_R_X73Y119_SLICE_X110Y119_AO5),
.O6(CLBLL_R_X73Y119_SLICE_X110Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y119_SLICE_X111Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y119_SLICE_X110Y119_AQ),
.Q(CLBLL_R_X73Y119_SLICE_X111Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y119_SLICE_X111Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y119_SLICE_X111Y119_DO5),
.O6(CLBLL_R_X73Y119_SLICE_X111Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y119_SLICE_X111Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y119_SLICE_X111Y119_CO5),
.O6(CLBLL_R_X73Y119_SLICE_X111Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y119_SLICE_X111Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y119_SLICE_X111Y119_BO5),
.O6(CLBLL_R_X73Y119_SLICE_X111Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y119_SLICE_X111Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y119_SLICE_X111Y119_AO5),
.O6(CLBLL_R_X73Y119_SLICE_X111Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y121_SLICE_X110Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y121_SLICE_X110Y121_AO6),
.Q(CLBLL_R_X73Y121_SLICE_X110Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y121_SLICE_X110Y121_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y121_SLICE_X110Y121_BO6),
.Q(CLBLL_R_X73Y121_SLICE_X110Y121_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h08aa080808aa0808)
  ) CLBLL_R_X73Y121_SLICE_X110Y121_DLUT (
.I0(CLBLL_R_X73Y123_SLICE_X111Y123_AQ),
.I1(CLBLL_R_X73Y121_SLICE_X110Y121_AQ),
.I2(CLBLM_L_X72Y122_SLICE_X109Y122_AQ),
.I3(CLBLM_L_X72Y122_SLICE_X109Y122_A5Q),
.I4(CLBLL_R_X73Y121_SLICE_X110Y121_BQ),
.I5(1'b1),
.O5(CLBLL_R_X73Y121_SLICE_X110Y121_DO5),
.O6(CLBLL_R_X73Y121_SLICE_X110Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff33bffff333b)
  ) CLBLL_R_X73Y121_SLICE_X110Y121_CLUT (
.I0(CLBLL_R_X73Y121_SLICE_X111Y121_AQ),
.I1(CLBLL_R_X73Y121_SLICE_X111Y121_CO6),
.I2(CLBLM_L_X72Y122_SLICE_X109Y122_AQ),
.I3(CLBLM_L_X72Y122_SLICE_X109Y122_A5Q),
.I4(CLBLL_R_X73Y121_SLICE_X110Y121_DO6),
.I5(CLBLL_R_X73Y122_SLICE_X110Y122_BQ),
.O5(CLBLL_R_X73Y121_SLICE_X110Y121_CO5),
.O6(CLBLL_R_X73Y121_SLICE_X110Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccaffffccca0000)
  ) CLBLL_R_X73Y121_SLICE_X110Y121_BLUT (
.I0(CLBLL_R_X75Y128_SLICE_X114Y128_AO5),
.I1(CLBLL_R_X73Y121_SLICE_X110Y121_BQ),
.I2(CLBLL_R_X75Y128_SLICE_X115Y128_BO6),
.I3(CLBLL_R_X73Y122_SLICE_X110Y122_DO5),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X73Y122_SLICE_X110Y122_CQ),
.O5(CLBLL_R_X73Y121_SLICE_X110Y121_BO5),
.O6(CLBLL_R_X73Y121_SLICE_X110Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4e4e4e4ee44)
  ) CLBLL_R_X73Y121_SLICE_X110Y121_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X73Y122_SLICE_X110Y122_BQ),
.I2(CLBLL_R_X73Y121_SLICE_X110Y121_AQ),
.I3(CLBLL_R_X75Y128_SLICE_X114Y128_AO5),
.I4(CLBLL_R_X73Y122_SLICE_X111Y122_AQ),
.I5(CLBLL_R_X73Y122_SLICE_X110Y122_AO6),
.O5(CLBLL_R_X73Y121_SLICE_X110Y121_AO5),
.O6(CLBLL_R_X73Y121_SLICE_X110Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y121_SLICE_X111Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y121_SLICE_X111Y121_AO6),
.Q(CLBLL_R_X73Y121_SLICE_X111Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y121_SLICE_X111Y121_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y121_SLICE_X111Y121_BO6),
.Q(CLBLL_R_X73Y121_SLICE_X111Y121_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y121_SLICE_X111Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y121_SLICE_X111Y121_DO5),
.O6(CLBLL_R_X73Y121_SLICE_X111Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'habafbbffabafbbff)
  ) CLBLL_R_X73Y121_SLICE_X111Y121_CLUT (
.I0(CLBLL_R_X73Y123_SLICE_X111Y123_AQ),
.I1(CLBLL_R_X73Y122_SLICE_X110Y122_CQ),
.I2(CLBLL_R_X73Y121_SLICE_X111Y121_BQ),
.I3(CLBLM_L_X72Y122_SLICE_X109Y122_A5Q),
.I4(CLBLM_L_X72Y122_SLICE_X109Y122_AQ),
.I5(1'b1),
.O5(CLBLL_R_X73Y121_SLICE_X111Y121_CO5),
.O6(CLBLL_R_X73Y121_SLICE_X111Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88fda8dd885d08)
  ) CLBLL_R_X73Y121_SLICE_X111Y121_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X73Y121_SLICE_X111Y121_BQ),
.I2(CLBLL_R_X73Y122_SLICE_X111Y122_AO6),
.I3(CLBLL_R_X73Y121_SLICE_X110Y121_BQ),
.I4(CLBLL_R_X75Y128_SLICE_X115Y128_BO6),
.I5(CLBLL_R_X75Y128_SLICE_X114Y128_AO5),
.O5(CLBLL_R_X73Y121_SLICE_X111Y121_BO5),
.O6(CLBLL_R_X73Y121_SLICE_X111Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf2d0fffff2d00000)
  ) CLBLL_R_X73Y121_SLICE_X111Y121_ALUT (
.I0(CLBLM_L_X74Y122_SLICE_X112Y122_A5Q),
.I1(CLBLL_R_X73Y122_SLICE_X110Y122_AO6),
.I2(CLBLL_R_X73Y121_SLICE_X111Y121_AQ),
.I3(CLBLL_R_X75Y128_SLICE_X114Y128_AO5),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X73Y121_SLICE_X111Y121_BQ),
.O5(CLBLL_R_X73Y121_SLICE_X111Y121_AO5),
.O6(CLBLL_R_X73Y121_SLICE_X111Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y122_SLICE_X110Y122_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y122_SLICE_X110Y122_BO6),
.Q(CLBLL_R_X73Y122_SLICE_X110Y122_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y122_SLICE_X110Y122_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y122_SLICE_X110Y122_CO6),
.Q(CLBLL_R_X73Y122_SLICE_X110Y122_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccffccbbbbbbbb)
  ) CLBLL_R_X73Y122_SLICE_X110Y122_DLUT (
.I0(CLBLL_R_X73Y122_SLICE_X111Y122_AQ),
.I1(CLBLM_L_X74Y122_SLICE_X112Y122_A5Q),
.I2(1'b1),
.I3(CLBLL_R_X75Y128_SLICE_X115Y128_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y122_SLICE_X110Y122_DO5),
.O6(CLBLL_R_X73Y122_SLICE_X110Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffe4ffcc00e400)
  ) CLBLL_R_X73Y122_SLICE_X110Y122_CLUT (
.I0(CLBLL_R_X73Y122_SLICE_X111Y122_AQ),
.I1(CLBLL_R_X73Y122_SLICE_X110Y122_CQ),
.I2(CLBLL_R_X75Y128_SLICE_X114Y128_AO5),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLL_R_X73Y122_SLICE_X110Y122_DO6),
.I5(CLBLL_R_X73Y121_SLICE_X110Y121_AQ),
.O5(CLBLL_R_X73Y122_SLICE_X110Y122_CO5),
.O6(CLBLL_R_X73Y122_SLICE_X110Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa0a0acacacaca)
  ) CLBLL_R_X73Y122_SLICE_X110Y122_BLUT (
.I0(CLBLL_R_X73Y123_SLICE_X111Y123_CQ),
.I1(CLBLL_R_X73Y122_SLICE_X110Y122_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(1'b1),
.I4(CLBLL_R_X75Y128_SLICE_X114Y128_AO5),
.I5(CLBLL_R_X73Y122_SLICE_X110Y122_AO5),
.O5(CLBLL_R_X73Y122_SLICE_X110Y122_BO5),
.O6(CLBLL_R_X73Y122_SLICE_X110Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff333300001111)
  ) CLBLL_R_X73Y122_SLICE_X110Y122_ALUT (
.I0(CLBLM_L_X74Y122_SLICE_X112Y122_A5Q),
.I1(CLBLM_L_X74Y122_SLICE_X112Y122_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_R_X75Y128_SLICE_X115Y128_BO6),
.I5(1'b1),
.O5(CLBLL_R_X73Y122_SLICE_X110Y122_AO5),
.O6(CLBLL_R_X73Y122_SLICE_X110Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y122_SLICE_X111Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y122_SLICE_X111Y122_AO5),
.Q(CLBLL_R_X73Y122_SLICE_X111Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y122_SLICE_X111Y122_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y122_SLICE_X111Y122_BO6),
.Q(CLBLL_R_X73Y122_SLICE_X111Y122_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y122_SLICE_X111Y122_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y122_SLICE_X111Y122_CO6),
.Q(CLBLL_R_X73Y122_SLICE_X111Y122_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y122_SLICE_X111Y122_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y122_SLICE_X111Y122_DO6),
.Q(CLBLL_R_X73Y122_SLICE_X111Y122_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc66e4e4cc66e4e4)
  ) CLBLL_R_X73Y122_SLICE_X111Y122_DLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X73Y122_SLICE_X111Y122_CQ),
.I2(CLBLL_R_X73Y122_SLICE_X111Y122_DQ),
.I3(CLBLL_R_X73Y122_SLICE_X111Y122_BQ),
.I4(CLBLL_R_X73Y122_SLICE_X110Y122_AO5),
.I5(1'b1),
.O5(CLBLL_R_X73Y122_SLICE_X111Y122_DO5),
.O6(CLBLL_R_X73Y122_SLICE_X111Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88dd88df80)
  ) CLBLL_R_X73Y122_SLICE_X111Y122_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X73Y122_SLICE_X111Y122_CQ),
.I2(CLBLM_L_X74Y122_SLICE_X112Y122_A5Q),
.I3(CLBLL_R_X73Y122_SLICE_X111Y122_BQ),
.I4(CLBLL_R_X75Y128_SLICE_X115Y128_BO6),
.I5(CLBLM_L_X74Y122_SLICE_X112Y122_AQ),
.O5(CLBLL_R_X73Y122_SLICE_X111Y122_CO5),
.O6(CLBLL_R_X73Y122_SLICE_X111Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4eeeeeeee4444444)
  ) CLBLL_R_X73Y122_SLICE_X111Y122_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X73Y124_SLICE_X111Y124_BQ),
.I2(CLBLL_R_X71Y124_SLICE_X106Y124_CO6),
.I3(CLBLM_L_X72Y122_SLICE_X109Y122_AQ),
.I4(CLBLM_L_X72Y122_SLICE_X109Y122_A5Q),
.I5(CLBLL_R_X73Y122_SLICE_X111Y122_BQ),
.O5(CLBLL_R_X73Y122_SLICE_X111Y122_BO5),
.O6(CLBLL_R_X73Y122_SLICE_X111Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h30303030e4ffe400)
  ) CLBLL_R_X73Y122_SLICE_X111Y122_ALUT (
.I0(CLBLL_R_X75Y128_SLICE_X115Y128_BO6),
.I1(CLBLM_L_X74Y122_SLICE_X112Y122_AQ),
.I2(CLBLL_R_X73Y122_SLICE_X111Y122_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLL_R_X73Y123_SLICE_X110Y123_BQ),
.I5(1'b1),
.O5(CLBLL_R_X73Y122_SLICE_X111Y122_AO5),
.O6(CLBLL_R_X73Y122_SLICE_X111Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y123_SLICE_X110Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y124_SLICE_X114Y124_C5Q),
.Q(CLBLL_R_X73Y123_SLICE_X110Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y123_SLICE_X110Y123_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y122_SLICE_X112Y122_AQ),
.Q(CLBLL_R_X73Y123_SLICE_X110Y123_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y123_SLICE_X110Y123_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y123_SLICE_X111Y123_AQ),
.Q(CLBLL_R_X73Y123_SLICE_X110Y123_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y123_SLICE_X110Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y123_SLICE_X110Y123_DO5),
.O6(CLBLL_R_X73Y123_SLICE_X110Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y123_SLICE_X110Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y123_SLICE_X110Y123_CO5),
.O6(CLBLL_R_X73Y123_SLICE_X110Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y123_SLICE_X110Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y123_SLICE_X110Y123_BO5),
.O6(CLBLL_R_X73Y123_SLICE_X110Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y123_SLICE_X110Y123_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y123_SLICE_X110Y123_AO5),
.O6(CLBLL_R_X73Y123_SLICE_X110Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y123_SLICE_X111Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y123_SLICE_X111Y123_AO6),
.Q(CLBLL_R_X73Y123_SLICE_X111Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y123_SLICE_X111Y123_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y123_SLICE_X111Y123_BO6),
.Q(CLBLL_R_X73Y123_SLICE_X111Y123_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y123_SLICE_X111Y123_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y123_SLICE_X111Y123_CO6),
.Q(CLBLL_R_X73Y123_SLICE_X111Y123_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y123_SLICE_X111Y123_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y123_SLICE_X111Y123_DO6),
.Q(CLBLL_R_X73Y123_SLICE_X111Y123_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000e1ffe100)
  ) CLBLL_R_X73Y123_SLICE_X111Y123_DLUT (
.I0(CLBLM_L_X74Y122_SLICE_X112Y122_AQ),
.I1(CLBLM_L_X74Y122_SLICE_X112Y122_A5Q),
.I2(CLBLL_R_X73Y123_SLICE_X111Y123_DQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLL_R_X73Y122_SLICE_X111Y122_DQ),
.I5(CLBLL_R_X75Y128_SLICE_X115Y128_BO6),
.O5(CLBLL_R_X73Y123_SLICE_X111Y123_DO5),
.O6(CLBLL_R_X73Y123_SLICE_X111Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cfc0cfc0df80)
  ) CLBLL_R_X73Y123_SLICE_X111Y123_CLUT (
.I0(CLBLM_L_X74Y122_SLICE_X112Y122_AQ),
.I1(CLBLL_R_X73Y123_SLICE_X111Y123_CQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLL_R_X73Y123_SLICE_X111Y123_BQ),
.I4(CLBLM_L_X74Y122_SLICE_X112Y122_A5Q),
.I5(CLBLL_R_X75Y128_SLICE_X115Y128_BO6),
.O5(CLBLL_R_X73Y123_SLICE_X111Y123_CO5),
.O6(CLBLL_R_X73Y123_SLICE_X111Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc37aaaaccc8aaaa)
  ) CLBLL_R_X73Y123_SLICE_X111Y123_BLUT (
.I0(CLBLM_L_X74Y122_SLICE_X112Y122_A5Q),
.I1(CLBLL_R_X73Y123_SLICE_X111Y123_BQ),
.I2(CLBLM_L_X74Y122_SLICE_X112Y122_AQ),
.I3(CLBLL_R_X75Y128_SLICE_X115Y128_BO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X74Y128_SLICE_X113Y128_AO5),
.O5(CLBLL_R_X73Y123_SLICE_X111Y123_BO5),
.O6(CLBLL_R_X73Y123_SLICE_X111Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hef20ef20ff77ff77)
  ) CLBLL_R_X73Y123_SLICE_X111Y123_ALUT (
.I0(CLBLL_R_X73Y123_SLICE_X111Y123_AQ),
.I1(CLBLL_R_X71Y124_SLICE_X106Y124_CO6),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X72Y122_SLICE_X109Y122_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y123_SLICE_X111Y123_AO5),
.O6(CLBLL_R_X73Y123_SLICE_X111Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y124_SLICE_X110Y124_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y124_SLICE_X110Y124_CO6),
.Q(CLBLL_R_X73Y124_SLICE_X110Y124_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y124_SLICE_X110Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y124_SLICE_X110Y124_AO6),
.Q(CLBLL_R_X73Y124_SLICE_X110Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y124_SLICE_X110Y124_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y124_SLICE_X110Y124_BO5),
.Q(CLBLL_R_X73Y124_SLICE_X110Y124_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y124_SLICE_X110Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y124_SLICE_X110Y124_DO5),
.O6(CLBLL_R_X73Y124_SLICE_X110Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffdd2200ffff33ff)
  ) CLBLL_R_X73Y124_SLICE_X110Y124_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X72Y124_SLICE_X108Y124_BO6),
.I2(1'b1),
.I3(CLBLL_R_X73Y124_SLICE_X110Y124_A5Q),
.I4(CLBLM_L_X72Y124_SLICE_X109Y124_AQ),
.I5(1'b1),
.O5(CLBLL_R_X73Y124_SLICE_X110Y124_CO5),
.O6(CLBLL_R_X73Y124_SLICE_X110Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccffffefe04f40)
  ) CLBLL_R_X73Y124_SLICE_X110Y124_BLUT (
.I0(CLBLM_L_X72Y124_SLICE_X108Y124_BO6),
.I1(CLBLL_R_X73Y124_SLICE_X110Y124_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLL_R_X73Y125_SLICE_X110Y125_AQ),
.I4(CLBLL_R_X73Y124_SLICE_X110Y124_A5Q),
.I5(1'b1),
.O5(CLBLL_R_X73Y124_SLICE_X110Y124_BO5),
.O6(CLBLL_R_X73Y124_SLICE_X110Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf050ccccf0facccc)
  ) CLBLL_R_X73Y124_SLICE_X110Y124_ALUT (
.I0(CLBLM_L_X72Y124_SLICE_X108Y124_BO6),
.I1(CLBLL_R_X73Y126_SLICE_X110Y126_AQ),
.I2(CLBLL_R_X73Y124_SLICE_X110Y124_AQ),
.I3(CLBLL_R_X73Y124_SLICE_X110Y124_BO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X74Y126_SLICE_X112Y126_CO6),
.O5(CLBLL_R_X73Y124_SLICE_X110Y124_AO5),
.O6(CLBLL_R_X73Y124_SLICE_X110Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y124_SLICE_X111Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y124_SLICE_X111Y124_AO6),
.Q(CLBLL_R_X73Y124_SLICE_X111Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y124_SLICE_X111Y124_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y124_SLICE_X111Y124_BO6),
.Q(CLBLL_R_X73Y124_SLICE_X111Y124_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y124_SLICE_X111Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y124_SLICE_X111Y124_DO5),
.O6(CLBLL_R_X73Y124_SLICE_X111Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y124_SLICE_X111Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y124_SLICE_X111Y124_CO5),
.O6(CLBLL_R_X73Y124_SLICE_X111Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc0fccf0f0f0f0f0)
  ) CLBLL_R_X73Y124_SLICE_X111Y124_BLUT (
.I0(1'b1),
.I1(CLBLL_R_X73Y124_SLICE_X111Y124_BQ),
.I2(CLBLL_R_X73Y124_SLICE_X111Y124_AQ),
.I3(CLBLL_R_X73Y123_SLICE_X111Y123_AO5),
.I4(CLBLL_R_X73Y123_SLICE_X111Y123_CQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLL_R_X73Y124_SLICE_X111Y124_BO5),
.O6(CLBLL_R_X73Y124_SLICE_X111Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5fdfa020f5f5a0a0)
  ) CLBLL_R_X73Y124_SLICE_X111Y124_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X73Y123_SLICE_X111Y123_AQ),
.I2(CLBLL_R_X73Y124_SLICE_X111Y124_AQ),
.I3(CLBLM_L_X72Y122_SLICE_X109Y122_AQ),
.I4(CLBLM_L_X72Y123_SLICE_X108Y123_AQ),
.I5(CLBLL_R_X71Y124_SLICE_X106Y124_CO6),
.O5(CLBLL_R_X73Y124_SLICE_X111Y124_AO5),
.O6(CLBLL_R_X73Y124_SLICE_X111Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y125_SLICE_X110Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y124_SLICE_X110Y124_A5Q),
.Q(CLBLL_R_X73Y125_SLICE_X110Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000010001)
  ) CLBLL_R_X73Y125_SLICE_X110Y125_DLUT (
.I0(CLBLL_R_X73Y123_SLICE_X110Y123_BQ),
.I1(CLBLM_L_X72Y127_SLICE_X109Y127_BQ),
.I2(CLBLL_R_X73Y125_SLICE_X110Y125_AQ),
.I3(CLBLM_L_X74Y125_SLICE_X112Y125_BO6),
.I4(1'b1),
.I5(CLBLM_L_X72Y127_SLICE_X109Y127_AQ),
.O5(CLBLL_R_X73Y125_SLICE_X110Y125_DO5),
.O6(CLBLL_R_X73Y125_SLICE_X110Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00a000a0aaaa00a0)
  ) CLBLL_R_X73Y125_SLICE_X110Y125_CLUT (
.I0(CLBLL_R_X73Y124_SLICE_X110Y124_A5Q),
.I1(1'b1),
.I2(CLBLL_R_X73Y126_SLICE_X111Y126_AQ),
.I3(CLBLM_L_X72Y124_SLICE_X109Y124_AQ),
.I4(CLBLM_L_X74Y126_SLICE_X112Y126_DQ),
.I5(CLBLL_R_X73Y124_SLICE_X110Y124_BQ),
.O5(CLBLL_R_X73Y125_SLICE_X110Y125_CO5),
.O6(CLBLL_R_X73Y125_SLICE_X110Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ff8800008888)
  ) CLBLL_R_X73Y125_SLICE_X110Y125_BLUT (
.I0(CLBLM_L_X74Y126_SLICE_X112Y126_AQ),
.I1(CLBLL_R_X73Y124_SLICE_X110Y124_BQ),
.I2(1'b1),
.I3(CLBLL_R_X73Y126_SLICE_X111Y126_DQ),
.I4(CLBLL_R_X73Y124_SLICE_X110Y124_A5Q),
.I5(CLBLM_L_X72Y124_SLICE_X109Y124_AQ),
.O5(CLBLL_R_X73Y125_SLICE_X110Y125_BO5),
.O6(CLBLL_R_X73Y125_SLICE_X110Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffeabbeaaa)
  ) CLBLL_R_X73Y125_SLICE_X110Y125_ALUT (
.I0(CLBLL_R_X73Y125_SLICE_X110Y125_BO6),
.I1(CLBLL_R_X73Y124_SLICE_X110Y124_BQ),
.I2(CLBLL_R_X73Y126_SLICE_X111Y126_CQ),
.I3(CLBLM_L_X72Y124_SLICE_X109Y124_AQ),
.I4(CLBLL_R_X73Y126_SLICE_X110Y126_AQ),
.I5(CLBLL_R_X73Y125_SLICE_X110Y125_CO6),
.O5(CLBLL_R_X73Y125_SLICE_X110Y125_AO5),
.O6(CLBLL_R_X73Y125_SLICE_X110Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y125_SLICE_X111Y125_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y125_SLICE_X111Y125_AO5),
.Q(CLBLL_R_X73Y125_SLICE_X111Y125_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y125_SLICE_X111Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y125_SLICE_X111Y125_AO6),
.Q(CLBLL_R_X73Y125_SLICE_X111Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y125_SLICE_X111Y125_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y125_SLICE_X111Y125_BO6),
.Q(CLBLL_R_X73Y125_SLICE_X111Y125_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y125_SLICE_X111Y125_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y125_SLICE_X111Y125_CO6),
.Q(CLBLL_R_X73Y125_SLICE_X111Y125_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y125_SLICE_X111Y125_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y125_SLICE_X111Y125_DO6),
.Q(CLBLL_R_X73Y125_SLICE_X111Y125_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4e4e4e4e44e)
  ) CLBLL_R_X73Y125_SLICE_X111Y125_DLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X73Y125_SLICE_X111Y125_CQ),
.I2(CLBLL_R_X73Y125_SLICE_X111Y125_DQ),
.I3(CLBLM_L_X74Y126_SLICE_X113Y126_AQ),
.I4(CLBLM_L_X74Y126_SLICE_X113Y126_A5Q),
.I5(CLBLL_R_X75Y128_SLICE_X115Y128_AO6),
.O5(CLBLL_R_X73Y125_SLICE_X111Y125_DO5),
.O6(CLBLL_R_X73Y125_SLICE_X111Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd08fd085da85da8)
  ) CLBLL_R_X73Y125_SLICE_X111Y125_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X73Y125_SLICE_X111Y125_CQ),
.I2(CLBLL_R_X73Y126_SLICE_X111Y126_BO5),
.I3(CLBLL_R_X73Y125_SLICE_X111Y125_BQ),
.I4(1'b1),
.I5(CLBLM_L_X72Y125_SLICE_X109Y125_BQ),
.O5(CLBLL_R_X73Y125_SLICE_X111Y125_CO5),
.O6(CLBLL_R_X73Y125_SLICE_X111Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0f0ccd8f0f0)
  ) CLBLL_R_X73Y125_SLICE_X111Y125_BLUT (
.I0(CLBLM_L_X74Y126_SLICE_X113Y126_AQ),
.I1(CLBLL_R_X73Y125_SLICE_X111Y125_BQ),
.I2(CLBLM_L_X72Y125_SLICE_X109Y125_BQ),
.I3(CLBLL_R_X75Y128_SLICE_X115Y128_AO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X74Y126_SLICE_X113Y126_A5Q),
.O5(CLBLL_R_X73Y125_SLICE_X111Y125_BO5),
.O6(CLBLL_R_X73Y125_SLICE_X111Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f0f0ccccaaaa)
  ) CLBLL_R_X73Y125_SLICE_X111Y125_ALUT (
.I0(CLBLM_L_X70Y125_SLICE_X104Y125_BQ),
.I1(CLBLM_L_X70Y125_SLICE_X105Y125_CO6),
.I2(CLBLL_R_X75Y124_SLICE_X114Y124_AQ),
.I3(CLBLM_L_X74Y125_SLICE_X112Y125_AO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLL_R_X73Y125_SLICE_X111Y125_AO5),
.O6(CLBLL_R_X73Y125_SLICE_X111Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y126_SLICE_X110Y126_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y126_SLICE_X110Y126_CO5),
.Q(CLBLL_R_X73Y126_SLICE_X110Y126_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y126_SLICE_X110Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y126_SLICE_X110Y126_AO6),
.Q(CLBLL_R_X73Y126_SLICE_X110Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y126_SLICE_X110Y126_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y126_SLICE_X110Y126_BO6),
.Q(CLBLL_R_X73Y126_SLICE_X110Y126_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y126_SLICE_X110Y126_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y126_SLICE_X110Y126_DO6),
.Q(CLBLL_R_X73Y126_SLICE_X110Y126_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5af0ccccf0f0cccc)
  ) CLBLL_R_X73Y126_SLICE_X110Y126_DLUT (
.I0(CLBLL_R_X71Y126_SLICE_X106Y126_CO6),
.I1(CLBLL_R_X71Y127_SLICE_X107Y127_DQ),
.I2(CLBLL_R_X73Y126_SLICE_X110Y126_DQ),
.I3(CLBLL_R_X73Y126_SLICE_X110Y126_A5Q),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X72Y126_SLICE_X109Y126_AQ),
.O5(CLBLL_R_X73Y126_SLICE_X110Y126_DO5),
.O6(CLBLL_R_X73Y126_SLICE_X110Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33ff33df8fd080)
  ) CLBLL_R_X73Y126_SLICE_X110Y126_CLUT (
.I0(CLBLL_R_X71Y126_SLICE_X106Y126_CO6),
.I1(CLBLL_R_X71Y127_SLICE_X107Y127_AQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLL_R_X73Y126_SLICE_X110Y126_A5Q),
.I4(CLBLM_L_X74Y127_SLICE_X112Y127_AQ),
.I5(1'b1),
.O5(CLBLL_R_X73Y126_SLICE_X110Y126_CO5),
.O6(CLBLL_R_X73Y126_SLICE_X110Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccff005c5cff00)
  ) CLBLL_R_X73Y126_SLICE_X110Y126_BLUT (
.I0(CLBLL_R_X73Y127_SLICE_X110Y127_CO6),
.I1(CLBLL_R_X73Y126_SLICE_X110Y126_BQ),
.I2(CLBLL_R_X71Y126_SLICE_X106Y126_CO6),
.I3(CLBLL_R_X73Y127_SLICE_X110Y127_AQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X73Y126_SLICE_X110Y126_CO6),
.O5(CLBLL_R_X73Y126_SLICE_X110Y126_BO5),
.O6(CLBLL_R_X73Y126_SLICE_X110Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f0aaaac0f0aaaa)
  ) CLBLL_R_X73Y126_SLICE_X110Y126_ALUT (
.I0(CLBLL_R_X73Y126_SLICE_X111Y126_DQ),
.I1(CLBLL_R_X73Y126_SLICE_X111Y126_BO6),
.I2(CLBLL_R_X73Y126_SLICE_X110Y126_AQ),
.I3(CLBLM_L_X74Y126_SLICE_X113Y126_A5Q),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X75Y128_SLICE_X114Y128_AO6),
.O5(CLBLL_R_X73Y126_SLICE_X110Y126_AO5),
.O6(CLBLL_R_X73Y126_SLICE_X110Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y126_SLICE_X111Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y126_SLICE_X111Y126_AO6),
.Q(CLBLL_R_X73Y126_SLICE_X111Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y126_SLICE_X111Y126_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y126_SLICE_X111Y126_CO6),
.Q(CLBLL_R_X73Y126_SLICE_X111Y126_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y126_SLICE_X111Y126_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y126_SLICE_X111Y126_DO6),
.Q(CLBLL_R_X73Y126_SLICE_X111Y126_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7c4f3c0b380f3c0)
  ) CLBLL_R_X73Y126_SLICE_X111Y126_DLUT (
.I0(CLBLL_R_X75Y128_SLICE_X115Y128_AO6),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLL_R_X73Y126_SLICE_X111Y126_DQ),
.I3(CLBLM_L_X74Y126_SLICE_X112Y126_DQ),
.I4(CLBLM_L_X74Y126_SLICE_X112Y126_CO6),
.I5(CLBLL_R_X75Y128_SLICE_X114Y128_AO6),
.O5(CLBLL_R_X73Y126_SLICE_X111Y126_DO5),
.O6(CLBLL_R_X73Y126_SLICE_X111Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50d8d8fa50d8d8)
  ) CLBLL_R_X73Y126_SLICE_X111Y126_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X73Y126_SLICE_X111Y126_CQ),
.I2(CLBLM_L_X74Y126_SLICE_X113Y126_CQ),
.I3(CLBLL_R_X75Y128_SLICE_X114Y128_AO6),
.I4(CLBLL_R_X73Y126_SLICE_X111Y126_BO5),
.I5(1'b1),
.O5(CLBLL_R_X73Y126_SLICE_X111Y126_CO5),
.O6(CLBLL_R_X73Y126_SLICE_X111Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff555500001111)
  ) CLBLL_R_X73Y126_SLICE_X111Y126_BLUT (
.I0(CLBLM_L_X74Y126_SLICE_X113Y126_AQ),
.I1(CLBLM_L_X74Y126_SLICE_X113Y126_A5Q),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_R_X75Y128_SLICE_X115Y128_AO6),
.I5(1'b1),
.O5(CLBLL_R_X73Y126_SLICE_X111Y126_BO5),
.O6(CLBLL_R_X73Y126_SLICE_X111Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f5ccccf0a0cccc)
  ) CLBLL_R_X73Y126_SLICE_X111Y126_ALUT (
.I0(CLBLM_L_X74Y126_SLICE_X112Y126_A5Q),
.I1(CLBLL_R_X73Y126_SLICE_X111Y126_CQ),
.I2(CLBLL_R_X73Y126_SLICE_X111Y126_AQ),
.I3(CLBLL_R_X73Y126_SLICE_X111Y126_BO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X75Y128_SLICE_X114Y128_AO6),
.O5(CLBLL_R_X73Y126_SLICE_X111Y126_AO5),
.O6(CLBLL_R_X73Y126_SLICE_X111Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y127_SLICE_X110Y127_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y127_SLICE_X110Y127_CO5),
.Q(CLBLL_R_X73Y127_SLICE_X110Y127_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y127_SLICE_X110Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y127_SLICE_X110Y127_AO6),
.Q(CLBLL_R_X73Y127_SLICE_X110Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y127_SLICE_X110Y127_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y127_SLICE_X110Y127_BO6),
.Q(CLBLL_R_X73Y127_SLICE_X110Y127_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y127_SLICE_X110Y127_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y127_SLICE_X110Y127_DO6),
.Q(CLBLL_R_X73Y127_SLICE_X110Y127_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4e4e4e4ee44)
  ) CLBLL_R_X73Y127_SLICE_X110Y127_DLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X75Y127_SLICE_X114Y127_BQ),
.I2(CLBLL_R_X73Y127_SLICE_X110Y127_DQ),
.I3(CLBLL_R_X75Y128_SLICE_X114Y128_BO6),
.I4(CLBLL_R_X75Y128_SLICE_X115Y128_CO6),
.I5(CLBLL_R_X75Y127_SLICE_X114Y127_CO5),
.O5(CLBLL_R_X73Y127_SLICE_X110Y127_DO5),
.O6(CLBLL_R_X73Y127_SLICE_X110Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f000f00fd75a820)
  ) CLBLL_R_X73Y127_SLICE_X110Y127_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X75Y128_SLICE_X115Y128_CO6),
.I2(CLBLL_R_X75Y127_SLICE_X114Y127_AQ),
.I3(CLBLL_R_X73Y127_SLICE_X110Y127_A5Q),
.I4(CLBLM_L_X72Y127_SLICE_X109Y127_AQ),
.I5(1'b1),
.O5(CLBLL_R_X73Y127_SLICE_X110Y127_CO5),
.O6(CLBLL_R_X73Y127_SLICE_X110Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88f0f0ccccf0f0)
  ) CLBLL_R_X73Y127_SLICE_X110Y127_BLUT (
.I0(CLBLL_R_X75Y128_SLICE_X115Y128_CO6),
.I1(CLBLL_R_X73Y127_SLICE_X110Y127_BQ),
.I2(CLBLL_R_X73Y127_SLICE_X110Y127_DQ),
.I3(CLBLL_R_X75Y128_SLICE_X114Y128_BO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X73Y127_SLICE_X110Y127_CO6),
.O5(CLBLL_R_X73Y127_SLICE_X110Y127_BO5),
.O6(CLBLL_R_X73Y127_SLICE_X110Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf2d0f2d0ffff0000)
  ) CLBLL_R_X73Y127_SLICE_X110Y127_ALUT (
.I0(CLBLL_R_X75Y127_SLICE_X114Y127_A5Q),
.I1(CLBLL_R_X73Y127_SLICE_X111Y127_BO6),
.I2(CLBLL_R_X73Y127_SLICE_X110Y127_AQ),
.I3(CLBLL_R_X75Y128_SLICE_X114Y128_BO6),
.I4(CLBLL_R_X73Y127_SLICE_X110Y127_BQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLL_R_X73Y127_SLICE_X110Y127_AO5),
.O6(CLBLL_R_X73Y127_SLICE_X110Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y127_SLICE_X111Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y127_SLICE_X111Y127_AO6),
.Q(CLBLL_R_X73Y127_SLICE_X111Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y127_SLICE_X111Y127_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y127_SLICE_X111Y127_CO6),
.Q(CLBLL_R_X73Y127_SLICE_X111Y127_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y127_SLICE_X111Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y127_SLICE_X111Y127_DO5),
.O6(CLBLL_R_X73Y127_SLICE_X111Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50d8d8fa50d8d8)
  ) CLBLL_R_X73Y127_SLICE_X111Y127_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X73Y127_SLICE_X111Y127_CQ),
.I2(CLBLL_R_X75Y127_SLICE_X114Y127_DQ),
.I3(CLBLL_R_X75Y128_SLICE_X114Y128_BO6),
.I4(CLBLL_R_X73Y127_SLICE_X111Y127_BO5),
.I5(1'b1),
.O5(CLBLL_R_X73Y127_SLICE_X111Y127_CO5),
.O6(CLBLL_R_X73Y127_SLICE_X111Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccffff00001111)
  ) CLBLL_R_X73Y127_SLICE_X111Y127_BLUT (
.I0(CLBLL_R_X75Y127_SLICE_X114Y127_A5Q),
.I1(CLBLL_R_X75Y128_SLICE_X115Y128_CO6),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_R_X75Y127_SLICE_X114Y127_AQ),
.I5(1'b1),
.O5(CLBLL_R_X73Y127_SLICE_X111Y127_BO5),
.O6(CLBLL_R_X73Y127_SLICE_X111Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0e4f0e4ffff0000)
  ) CLBLL_R_X73Y127_SLICE_X111Y127_ALUT (
.I0(CLBLL_R_X73Y127_SLICE_X110Y127_A5Q),
.I1(CLBLL_R_X75Y128_SLICE_X114Y128_BO6),
.I2(CLBLL_R_X73Y127_SLICE_X111Y127_AQ),
.I3(CLBLL_R_X73Y127_SLICE_X111Y127_BO6),
.I4(CLBLL_R_X73Y127_SLICE_X111Y127_CQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLL_R_X73Y127_SLICE_X111Y127_AO5),
.O6(CLBLL_R_X73Y127_SLICE_X111Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y128_SLICE_X110Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y128_SLICE_X110Y128_AO6),
.Q(CLBLL_R_X73Y128_SLICE_X110Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y128_SLICE_X110Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y128_SLICE_X110Y128_DO5),
.O6(CLBLL_R_X73Y128_SLICE_X110Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y128_SLICE_X110Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y128_SLICE_X110Y128_CO5),
.O6(CLBLL_R_X73Y128_SLICE_X110Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y128_SLICE_X110Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y128_SLICE_X110Y128_BO5),
.O6(CLBLL_R_X73Y128_SLICE_X110Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0f5a0d782)
  ) CLBLL_R_X73Y128_SLICE_X110Y128_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X75Y127_SLICE_X114Y127_A5Q),
.I2(CLBLL_R_X73Y128_SLICE_X110Y128_AQ),
.I3(CLBLL_R_X73Y128_SLICE_X111Y128_BQ),
.I4(CLBLL_R_X75Y127_SLICE_X114Y127_AQ),
.I5(CLBLL_R_X75Y128_SLICE_X115Y128_CO6),
.O5(CLBLL_R_X73Y128_SLICE_X110Y128_AO5),
.O6(CLBLL_R_X73Y128_SLICE_X110Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y128_SLICE_X111Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y128_SLICE_X111Y128_AO6),
.Q(CLBLL_R_X73Y128_SLICE_X111Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y128_SLICE_X111Y128_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y128_SLICE_X111Y128_BO6),
.Q(CLBLL_R_X73Y128_SLICE_X111Y128_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y128_SLICE_X111Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y128_SLICE_X111Y128_DO5),
.O6(CLBLL_R_X73Y128_SLICE_X111Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y128_SLICE_X111Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y128_SLICE_X111Y128_CO5),
.O6(CLBLL_R_X73Y128_SLICE_X111Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4f0f04e4ef0f0)
  ) CLBLL_R_X73Y128_SLICE_X111Y128_BLUT (
.I0(CLBLL_R_X73Y127_SLICE_X111Y127_BO5),
.I1(CLBLL_R_X73Y128_SLICE_X111Y128_BQ),
.I2(CLBLL_R_X73Y128_SLICE_X111Y128_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X73Y126_SLICE_X110Y126_DQ),
.O5(CLBLL_R_X73Y128_SLICE_X111Y128_BO5),
.O6(CLBLL_R_X73Y128_SLICE_X111Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2e2e2e2e2e2aa)
  ) CLBLL_R_X73Y128_SLICE_X111Y128_ALUT (
.I0(CLBLL_R_X73Y126_SLICE_X110Y126_DQ),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLL_R_X73Y128_SLICE_X111Y128_AQ),
.I3(CLBLL_R_X75Y127_SLICE_X114Y127_A5Q),
.I4(CLBLL_R_X75Y127_SLICE_X114Y127_AQ),
.I5(CLBLL_R_X75Y128_SLICE_X115Y128_CO6),
.O5(CLBLL_R_X73Y128_SLICE_X111Y128_AO5),
.O6(CLBLL_R_X73Y128_SLICE_X111Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y131_SLICE_X110Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y136_SLICE_X105Y136_A5Q),
.Q(CLBLL_R_X73Y131_SLICE_X110Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y131_SLICE_X110Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y131_SLICE_X110Y131_DO5),
.O6(CLBLL_R_X73Y131_SLICE_X110Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y131_SLICE_X110Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y131_SLICE_X110Y131_CO5),
.O6(CLBLL_R_X73Y131_SLICE_X110Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y131_SLICE_X110Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y131_SLICE_X110Y131_BO5),
.O6(CLBLL_R_X73Y131_SLICE_X110Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y131_SLICE_X110Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y131_SLICE_X110Y131_AO5),
.O6(CLBLL_R_X73Y131_SLICE_X110Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y131_SLICE_X111Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y131_SLICE_X111Y131_AO6),
.Q(CLBLL_R_X73Y131_SLICE_X111Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y131_SLICE_X111Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y131_SLICE_X111Y131_DO5),
.O6(CLBLL_R_X73Y131_SLICE_X111Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y131_SLICE_X111Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y131_SLICE_X111Y131_CO5),
.O6(CLBLL_R_X73Y131_SLICE_X111Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y131_SLICE_X111Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y131_SLICE_X111Y131_BO5),
.O6(CLBLL_R_X73Y131_SLICE_X111Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbf3bbf388c088c0)
  ) CLBLL_R_X73Y131_SLICE_X111Y131_ALUT (
.I0(CLBLM_L_X70Y136_SLICE_X105Y136_A5Q),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLL_R_X73Y131_SLICE_X111Y131_AQ),
.I3(CLBLM_L_X60Y94_SLICE_X90Y94_AQ),
.I4(1'b1),
.I5(CLBLM_L_X74Y132_SLICE_X112Y132_CQ),
.O5(CLBLL_R_X73Y131_SLICE_X111Y131_AO5),
.O6(CLBLL_R_X73Y131_SLICE_X111Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y132_SLICE_X110Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y132_SLICE_X110Y132_DO5),
.O6(CLBLL_R_X73Y132_SLICE_X110Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y132_SLICE_X110Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y132_SLICE_X110Y132_CO5),
.O6(CLBLL_R_X73Y132_SLICE_X110Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000080f0f0f0f0)
  ) CLBLL_R_X73Y132_SLICE_X110Y132_BLUT (
.I0(CLBLL_R_X73Y133_SLICE_X110Y133_A5Q),
.I1(CLBLM_L_X70Y136_SLICE_X105Y136_CO6),
.I2(CLBLL_R_X73Y132_SLICE_X111Y132_CO6),
.I3(CLBLM_L_X74Y134_SLICE_X113Y134_CQ),
.I4(CLBLM_L_X74Y134_SLICE_X113Y134_A5Q),
.I5(CLBLL_R_X73Y133_SLICE_X111Y133_A5Q),
.O5(CLBLL_R_X73Y132_SLICE_X110Y132_BO5),
.O6(CLBLL_R_X73Y132_SLICE_X110Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0fffffff5fff5)
  ) CLBLL_R_X73Y132_SLICE_X110Y132_ALUT (
.I0(CLBLM_L_X74Y132_SLICE_X112Y132_CQ),
.I1(1'b1),
.I2(CLBLM_L_X74Y132_SLICE_X113Y132_BQ),
.I3(CLBLL_R_X73Y132_SLICE_X111Y132_AO5),
.I4(CLBLL_R_X73Y131_SLICE_X110Y131_AQ),
.I5(1'b1),
.O5(CLBLL_R_X73Y132_SLICE_X110Y132_AO5),
.O6(CLBLL_R_X73Y132_SLICE_X110Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y132_SLICE_X111Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y132_SLICE_X111Y132_DO5),
.O6(CLBLL_R_X73Y132_SLICE_X111Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000050004000)
  ) CLBLL_R_X73Y132_SLICE_X111Y132_CLUT (
.I0(CLBLM_L_X74Y132_SLICE_X113Y132_BQ),
.I1(CLBLM_L_X76Y133_SLICE_X116Y133_BQ),
.I2(CLBLM_L_X76Y125_SLICE_X117Y125_BQ),
.I3(CLBLM_L_X74Y135_SLICE_X113Y135_BQ),
.I4(CLBLL_R_X75Y133_SLICE_X115Y133_AQ),
.I5(CLBLM_L_X76Y130_SLICE_X116Y130_DQ),
.O5(CLBLL_R_X73Y132_SLICE_X111Y132_CO5),
.O6(CLBLL_R_X73Y132_SLICE_X111Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000c0800000000)
  ) CLBLL_R_X73Y132_SLICE_X111Y132_BLUT (
.I0(CLBLL_R_X75Y133_SLICE_X115Y133_AQ),
.I1(CLBLM_L_X76Y125_SLICE_X117Y125_BQ),
.I2(CLBLM_L_X76Y130_SLICE_X116Y130_DQ),
.I3(CLBLM_L_X76Y133_SLICE_X116Y133_BQ),
.I4(CLBLM_L_X74Y133_SLICE_X112Y133_AQ),
.I5(CLBLM_L_X74Y135_SLICE_X113Y135_BQ),
.O5(CLBLL_R_X73Y132_SLICE_X111Y132_BO5),
.O6(CLBLL_R_X73Y132_SLICE_X111Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa8888f5fff7ff)
  ) CLBLL_R_X73Y132_SLICE_X111Y132_ALUT (
.I0(CLBLM_L_X74Y135_SLICE_X113Y135_BQ),
.I1(CLBLM_L_X76Y133_SLICE_X116Y133_BQ),
.I2(CLBLM_L_X76Y130_SLICE_X116Y130_DQ),
.I3(CLBLM_L_X76Y125_SLICE_X117Y125_BQ),
.I4(CLBLL_R_X75Y133_SLICE_X115Y133_AQ),
.I5(1'b1),
.O5(CLBLL_R_X73Y132_SLICE_X111Y132_AO5),
.O6(CLBLL_R_X73Y132_SLICE_X111Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y133_SLICE_X110Y133_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y133_SLICE_X110Y133_AO5),
.Q(CLBLL_R_X73Y133_SLICE_X110Y133_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y133_SLICE_X110Y133_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y133_SLICE_X110Y133_AO6),
.Q(CLBLL_R_X73Y133_SLICE_X110Y133_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y133_SLICE_X110Y133_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y133_SLICE_X110Y133_BO6),
.Q(CLBLL_R_X73Y133_SLICE_X110Y133_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y133_SLICE_X110Y133_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y133_SLICE_X110Y133_CO6),
.Q(CLBLL_R_X73Y133_SLICE_X110Y133_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2222dddd2020dfdf)
  ) CLBLL_R_X73Y133_SLICE_X110Y133_DLUT (
.I0(CLBLM_L_X74Y135_SLICE_X113Y135_BQ),
.I1(CLBLL_R_X73Y133_SLICE_X110Y133_CQ),
.I2(CLBLL_R_X75Y133_SLICE_X115Y133_AQ),
.I3(1'b1),
.I4(CLBLM_L_X74Y134_SLICE_X113Y134_AQ),
.I5(CLBLM_L_X76Y133_SLICE_X116Y133_BQ),
.O5(CLBLL_R_X73Y133_SLICE_X110Y133_DO5),
.O6(CLBLL_R_X73Y133_SLICE_X110Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hef5fef5faaaaaaaa)
  ) CLBLL_R_X73Y133_SLICE_X110Y133_CLUT (
.I0(CLBLL_R_X73Y133_SLICE_X110Y133_A5Q),
.I1(CLBLL_R_X73Y133_SLICE_X110Y133_AQ),
.I2(CLBLL_R_X75Y133_SLICE_X114Y133_AQ),
.I3(CLBLM_L_X70Y136_SLICE_X105Y136_A5Q),
.I4(1'b1),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLL_R_X73Y133_SLICE_X110Y133_CO5),
.O6(CLBLL_R_X73Y133_SLICE_X110Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcaca3a7acacaca8a)
  ) CLBLL_R_X73Y133_SLICE_X110Y133_BLUT (
.I0(CLBLM_L_X72Y133_SLICE_X108Y133_A5Q),
.I1(CLBLL_R_X73Y133_SLICE_X110Y133_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X72Y133_SLICE_X108Y133_AQ),
.I4(CLBLL_R_X73Y132_SLICE_X110Y132_BO6),
.I5(CLBLL_R_X73Y132_SLICE_X110Y132_AO5),
.O5(CLBLL_R_X73Y133_SLICE_X110Y133_BO5),
.O6(CLBLL_R_X73Y133_SLICE_X110Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00280028507a50d0)
  ) CLBLL_R_X73Y133_SLICE_X110Y133_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X75Y133_SLICE_X114Y133_CO5),
.I2(CLBLL_R_X73Y133_SLICE_X110Y133_AQ),
.I3(CLBLL_R_X75Y133_SLICE_X115Y133_BQ),
.I4(CLBLL_R_X73Y133_SLICE_X110Y133_A5Q),
.I5(1'b1),
.O5(CLBLL_R_X73Y133_SLICE_X110Y133_AO5),
.O6(CLBLL_R_X73Y133_SLICE_X110Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y133_SLICE_X111Y133_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X60Y94_SLICE_X90Y94_AQ),
.Q(CLBLL_R_X73Y133_SLICE_X111Y133_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y133_SLICE_X111Y133_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y133_SLICE_X111Y133_AO6),
.Q(CLBLL_R_X73Y133_SLICE_X111Y133_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ff7700aa0088)
  ) CLBLL_R_X73Y133_SLICE_X111Y133_DLUT (
.I0(CLBLM_L_X74Y135_SLICE_X113Y135_BQ),
.I1(CLBLM_L_X76Y133_SLICE_X116Y133_BQ),
.I2(1'b1),
.I3(CLBLL_R_X73Y133_SLICE_X110Y133_CQ),
.I4(CLBLL_R_X75Y133_SLICE_X115Y133_AQ),
.I5(CLBLM_L_X74Y133_SLICE_X112Y133_AQ),
.O5(CLBLL_R_X73Y133_SLICE_X111Y133_DO5),
.O6(CLBLL_R_X73Y133_SLICE_X111Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000c080000)
  ) CLBLL_R_X73Y133_SLICE_X111Y133_CLUT (
.I0(CLBLM_L_X76Y133_SLICE_X116Y133_BQ),
.I1(CLBLM_L_X74Y135_SLICE_X113Y135_BQ),
.I2(CLBLM_L_X74Y133_SLICE_X112Y133_CQ),
.I3(CLBLL_R_X75Y133_SLICE_X115Y133_AQ),
.I4(CLBLM_L_X76Y125_SLICE_X117Y125_BQ),
.I5(CLBLM_L_X76Y130_SLICE_X116Y130_DQ),
.O5(CLBLL_R_X73Y133_SLICE_X111Y133_CO5),
.O6(CLBLL_R_X73Y133_SLICE_X111Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0030000000200000)
  ) CLBLL_R_X73Y133_SLICE_X111Y133_BLUT (
.I0(CLBLL_R_X75Y133_SLICE_X115Y133_AQ),
.I1(CLBLM_L_X76Y130_SLICE_X116Y130_DQ),
.I2(CLBLM_L_X76Y125_SLICE_X117Y125_BQ),
.I3(CLBLM_L_X74Y134_SLICE_X113Y134_AQ),
.I4(CLBLM_L_X74Y135_SLICE_X113Y135_BQ),
.I5(CLBLM_L_X76Y133_SLICE_X116Y133_BQ),
.O5(CLBLL_R_X73Y133_SLICE_X111Y133_BO5),
.O6(CLBLL_R_X73Y133_SLICE_X111Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbb38880f3f3c0c0)
  ) CLBLL_R_X73Y133_SLICE_X111Y133_ALUT (
.I0(CLBLL_R_X73Y133_SLICE_X111Y133_DO6),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLL_R_X73Y133_SLICE_X111Y133_AQ),
.I3(CLBLM_L_X74Y132_SLICE_X112Y132_BO6),
.I4(CLBLM_L_X74Y134_SLICE_X113Y134_AQ),
.I5(CLBLM_L_X74Y134_SLICE_X112Y134_AO5),
.O5(CLBLL_R_X73Y133_SLICE_X111Y133_AO5),
.O6(CLBLL_R_X73Y133_SLICE_X111Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y134_SLICE_X110Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y134_SLICE_X110Y134_DO5),
.O6(CLBLL_R_X73Y134_SLICE_X110Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y134_SLICE_X110Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y134_SLICE_X110Y134_CO5),
.O6(CLBLL_R_X73Y134_SLICE_X110Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y134_SLICE_X110Y134_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y134_SLICE_X110Y134_BO5),
.O6(CLBLL_R_X73Y134_SLICE_X110Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55005500ff7f0000)
  ) CLBLL_R_X73Y134_SLICE_X110Y134_ALUT (
.I0(CLBLM_L_X74Y134_SLICE_X113Y134_CQ),
.I1(CLBLM_L_X70Y136_SLICE_X105Y136_CO6),
.I2(CLBLL_R_X73Y133_SLICE_X110Y133_A5Q),
.I3(CLBLM_L_X74Y134_SLICE_X113Y134_A5Q),
.I4(CLBLL_R_X71Y134_SLICE_X106Y134_AQ),
.I5(1'b1),
.O5(CLBLL_R_X73Y134_SLICE_X110Y134_AO5),
.O6(CLBLL_R_X73Y134_SLICE_X110Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X73Y134_SLICE_X111Y134_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y134_SLICE_X111Y134_AO6),
.Q(CLBLL_R_X73Y134_SLICE_X111Y134_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y134_SLICE_X111Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y134_SLICE_X111Y134_DO5),
.O6(CLBLL_R_X73Y134_SLICE_X111Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y134_SLICE_X111Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y134_SLICE_X111Y134_CO5),
.O6(CLBLL_R_X73Y134_SLICE_X111Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y134_SLICE_X111Y134_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y134_SLICE_X111Y134_BO5),
.O6(CLBLL_R_X73Y134_SLICE_X111Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f30fff00f100f00)
  ) CLBLL_R_X73Y134_SLICE_X111Y134_ALUT (
.I0(CLBLM_L_X74Y132_SLICE_X112Y132_A5Q),
.I1(CLBLL_R_X73Y133_SLICE_X110Y133_DO6),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X74Y132_SLICE_X112Y132_AQ),
.I4(CLBLM_L_X74Y134_SLICE_X112Y134_AO6),
.I5(CLBLL_R_X73Y134_SLICE_X111Y134_AQ),
.O5(CLBLL_R_X73Y134_SLICE_X111Y134_AO5),
.O6(CLBLL_R_X73Y134_SLICE_X111Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y103_SLICE_X114Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y103_SLICE_X114Y103_DO5),
.O6(CLBLL_R_X75Y103_SLICE_X114Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y103_SLICE_X114Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y103_SLICE_X114Y103_CO5),
.O6(CLBLL_R_X75Y103_SLICE_X114Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ff5f0000ffff)
  ) CLBLL_R_X75Y103_SLICE_X114Y103_BLUT (
.I0(CLBLM_L_X72Y104_SLICE_X109Y104_B5Q),
.I1(1'b1),
.I2(CLBLL_R_X73Y103_SLICE_X111Y103_A5Q),
.I3(CLBLM_L_X72Y104_SLICE_X109Y104_BQ),
.I4(CLBLL_R_X75Y103_SLICE_X114Y103_AO6),
.I5(CLBLM_L_X74Y104_SLICE_X112Y104_CQ),
.O5(CLBLL_R_X75Y103_SLICE_X114Y103_BO5),
.O6(CLBLL_R_X75Y103_SLICE_X114Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00400040ffff)
  ) CLBLL_R_X75Y103_SLICE_X114Y103_ALUT (
.I0(CLBLM_L_X72Y104_SLICE_X109Y104_B5Q),
.I1(CLBLM_L_X74Y104_SLICE_X112Y104_BQ),
.I2(CLBLL_R_X79Y104_SLICE_X122Y104_A5Q),
.I3(CLBLM_L_X72Y104_SLICE_X109Y104_BQ),
.I4(CLBLL_R_X75Y103_SLICE_X115Y103_AQ),
.I5(CLBLL_R_X73Y104_SLICE_X110Y104_A5Q),
.O5(CLBLL_R_X75Y103_SLICE_X114Y103_AO5),
.O6(CLBLL_R_X75Y103_SLICE_X114Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y103_SLICE_X115Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y103_SLICE_X115Y103_AO6),
.Q(CLBLL_R_X75Y103_SLICE_X115Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y103_SLICE_X115Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y103_SLICE_X115Y103_DO5),
.O6(CLBLL_R_X75Y103_SLICE_X115Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y103_SLICE_X115Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y103_SLICE_X115Y103_CO5),
.O6(CLBLL_R_X75Y103_SLICE_X115Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8b8b008b00000000)
  ) CLBLL_R_X75Y103_SLICE_X115Y103_BLUT (
.I0(CLBLL_R_X75Y103_SLICE_X115Y103_AQ),
.I1(CLBLL_R_X79Y104_SLICE_X122Y104_A5Q),
.I2(CLBLL_R_X73Y103_SLICE_X111Y103_A5Q),
.I3(CLBLL_R_X73Y103_SLICE_X110Y103_A5Q),
.I4(CLBLM_L_X60Y101_SLICE_X90Y101_AQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLL_R_X75Y103_SLICE_X115Y103_BO5),
.O6(CLBLL_R_X75Y103_SLICE_X115Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h40007300c000f300)
  ) CLBLL_R_X75Y103_SLICE_X115Y103_ALUT (
.I0(CLBLL_R_X75Y103_SLICE_X115Y103_AQ),
.I1(CLBLM_L_X62Y95_SLICE_X92Y95_AQ),
.I2(CLBLL_R_X73Y103_SLICE_X111Y103_A5Q),
.I3(CLBLL_R_X75Y103_SLICE_X115Y103_BO6),
.I4(CLBLM_L_X60Y101_SLICE_X90Y101_AQ),
.I5(CLBLL_R_X79Y104_SLICE_X122Y104_A5Q),
.O5(CLBLL_R_X75Y103_SLICE_X115Y103_AO5),
.O6(CLBLL_R_X75Y103_SLICE_X115Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y107_SLICE_X114Y107_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y107_SLICE_X93Y107_BQ),
.Q(CLBLL_R_X75Y107_SLICE_X114Y107_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y107_SLICE_X114Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y107_SLICE_X114Y107_DO5),
.O6(CLBLL_R_X75Y107_SLICE_X114Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y107_SLICE_X114Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y107_SLICE_X114Y107_CO5),
.O6(CLBLL_R_X75Y107_SLICE_X114Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y107_SLICE_X114Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y107_SLICE_X114Y107_BO5),
.O6(CLBLL_R_X75Y107_SLICE_X114Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y107_SLICE_X114Y107_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y107_SLICE_X114Y107_AO5),
.O6(CLBLL_R_X75Y107_SLICE_X114Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y107_SLICE_X115Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y107_SLICE_X115Y107_DO5),
.O6(CLBLL_R_X75Y107_SLICE_X115Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y107_SLICE_X115Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y107_SLICE_X115Y107_CO5),
.O6(CLBLL_R_X75Y107_SLICE_X115Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y107_SLICE_X115Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y107_SLICE_X115Y107_BO5),
.O6(CLBLL_R_X75Y107_SLICE_X115Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y107_SLICE_X115Y107_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y107_SLICE_X115Y107_AO5),
.O6(CLBLL_R_X75Y107_SLICE_X115Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y113_SLICE_X114Y113_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y109_SLICE_X113Y109_AQ),
.Q(CLBLL_R_X75Y113_SLICE_X114Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y113_SLICE_X114Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y113_SLICE_X114Y113_DO5),
.O6(CLBLL_R_X75Y113_SLICE_X114Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y113_SLICE_X114Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y113_SLICE_X114Y113_CO5),
.O6(CLBLL_R_X75Y113_SLICE_X114Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y113_SLICE_X114Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y113_SLICE_X114Y113_BO5),
.O6(CLBLL_R_X75Y113_SLICE_X114Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y113_SLICE_X114Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y113_SLICE_X114Y113_AO5),
.O6(CLBLL_R_X75Y113_SLICE_X114Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y113_SLICE_X115Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y113_SLICE_X115Y113_DO5),
.O6(CLBLL_R_X75Y113_SLICE_X115Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y113_SLICE_X115Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y113_SLICE_X115Y113_CO5),
.O6(CLBLL_R_X75Y113_SLICE_X115Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y113_SLICE_X115Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y113_SLICE_X115Y113_BO5),
.O6(CLBLL_R_X75Y113_SLICE_X115Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y113_SLICE_X115Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y113_SLICE_X115Y113_AO5),
.O6(CLBLL_R_X75Y113_SLICE_X115Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y121_SLICE_X114Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y121_SLICE_X114Y121_AO6),
.Q(CLBLL_R_X75Y121_SLICE_X114Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y121_SLICE_X114Y121_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y121_SLICE_X114Y121_BO6),
.Q(CLBLL_R_X75Y121_SLICE_X114Y121_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y121_SLICE_X114Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y121_SLICE_X114Y121_DO5),
.O6(CLBLL_R_X75Y121_SLICE_X114Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0707777707077777)
  ) CLBLL_R_X75Y121_SLICE_X114Y121_CLUT (
.I0(CLBLL_R_X75Y123_SLICE_X115Y123_AQ),
.I1(CLBLM_L_X76Y123_SLICE_X116Y123_BQ),
.I2(CLBLM_L_X74Y123_SLICE_X113Y123_DQ),
.I3(1'b1),
.I4(CLBLL_R_X75Y122_SLICE_X114Y122_CQ),
.I5(1'b1),
.O5(CLBLL_R_X75Y121_SLICE_X114Y121_CO5),
.O6(CLBLL_R_X75Y121_SLICE_X114Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hecccff006444ff00)
  ) CLBLL_R_X75Y121_SLICE_X114Y121_BLUT (
.I0(CLBLM_L_X74Y123_SLICE_X113Y123_CO5),
.I1(CLBLL_R_X75Y121_SLICE_X114Y121_BQ),
.I2(CLBLL_R_X75Y123_SLICE_X115Y123_AQ),
.I3(CLBLL_R_X75Y122_SLICE_X114Y122_AQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X75Y121_SLICE_X114Y121_CO6),
.O5(CLBLL_R_X75Y121_SLICE_X114Y121_BO5),
.O6(CLBLL_R_X75Y121_SLICE_X114Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff004f004f00)
  ) CLBLL_R_X75Y121_SLICE_X114Y121_ALUT (
.I0(CLBLM_L_X76Y123_SLICE_X116Y123_BQ),
.I1(CLBLL_R_X75Y121_SLICE_X114Y121_BQ),
.I2(CLBLL_R_X75Y123_SLICE_X115Y123_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X70Y105_SLICE_X105Y105_AQ),
.I5(1'b1),
.O5(CLBLL_R_X75Y121_SLICE_X114Y121_AO5),
.O6(CLBLL_R_X75Y121_SLICE_X114Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y121_SLICE_X115Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y121_SLICE_X115Y121_DO5),
.O6(CLBLL_R_X75Y121_SLICE_X115Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y121_SLICE_X115Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y121_SLICE_X115Y121_CO5),
.O6(CLBLL_R_X75Y121_SLICE_X115Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y121_SLICE_X115Y121_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y121_SLICE_X115Y121_BO5),
.O6(CLBLL_R_X75Y121_SLICE_X115Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y121_SLICE_X115Y121_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y121_SLICE_X115Y121_AO5),
.O6(CLBLL_R_X75Y121_SLICE_X115Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y122_SLICE_X114Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y122_SLICE_X114Y122_AO6),
.Q(CLBLL_R_X75Y122_SLICE_X114Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y122_SLICE_X114Y122_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y122_SLICE_X114Y122_BO6),
.Q(CLBLL_R_X75Y122_SLICE_X114Y122_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y122_SLICE_X114Y122_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y122_SLICE_X114Y122_CO6),
.Q(CLBLL_R_X75Y122_SLICE_X114Y122_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hddfddddddddddddd)
  ) CLBLL_R_X75Y122_SLICE_X114Y122_DLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X75Y122_SLICE_X114Y122_AQ),
.I2(CLBLL_R_X75Y122_SLICE_X114Y122_BQ),
.I3(CLBLL_R_X75Y123_SLICE_X115Y123_AQ),
.I4(CLBLL_R_X75Y123_SLICE_X114Y123_AO5),
.I5(CLBLM_L_X74Y122_SLICE_X113Y122_AQ),
.O5(CLBLL_R_X75Y122_SLICE_X114Y122_DO5),
.O6(CLBLL_R_X75Y122_SLICE_X114Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7d55dd55cc00cc00)
  ) CLBLL_R_X75Y122_SLICE_X114Y122_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X75Y122_SLICE_X114Y122_CQ),
.I2(CLBLM_L_X74Y123_SLICE_X113Y123_DQ),
.I3(CLBLL_R_X75Y121_SLICE_X114Y121_AO5),
.I4(CLBLL_R_X75Y123_SLICE_X114Y123_AO5),
.I5(CLBLM_L_X74Y122_SLICE_X113Y122_AQ),
.O5(CLBLL_R_X75Y122_SLICE_X114Y122_CO5),
.O6(CLBLL_R_X75Y122_SLICE_X114Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h60ffc0c0c0ffc0c0)
  ) CLBLL_R_X75Y122_SLICE_X114Y122_BLUT (
.I0(CLBLL_R_X75Y123_SLICE_X114Y123_CO6),
.I1(CLBLL_R_X75Y122_SLICE_X114Y122_BQ),
.I2(CLBLL_R_X75Y121_SLICE_X114Y121_AO5),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLL_R_X75Y122_SLICE_X114Y122_CQ),
.I5(CLBLM_L_X74Y122_SLICE_X113Y122_AQ),
.O5(CLBLL_R_X75Y122_SLICE_X114Y122_BO5),
.O6(CLBLL_R_X75Y122_SLICE_X114Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4cccccccc0c0c0c0)
  ) CLBLL_R_X75Y122_SLICE_X114Y122_ALUT (
.I0(CLBLM_L_X74Y123_SLICE_X113Y123_CO5),
.I1(CLBLL_R_X75Y122_SLICE_X114Y122_DO6),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X76Y123_SLICE_X116Y123_BQ),
.I4(CLBLL_R_X75Y121_SLICE_X114Y121_BQ),
.I5(CLBLL_R_X75Y123_SLICE_X115Y123_AQ),
.O5(CLBLL_R_X75Y122_SLICE_X114Y122_AO5),
.O6(CLBLL_R_X75Y122_SLICE_X114Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y122_SLICE_X115Y122_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y122_SLICE_X115Y122_AO5),
.Q(CLBLL_R_X75Y122_SLICE_X115Y122_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y122_SLICE_X115Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y122_SLICE_X115Y122_AO6),
.Q(CLBLL_R_X75Y122_SLICE_X115Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y122_SLICE_X115Y122_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y122_SLICE_X115Y122_BO6),
.Q(CLBLL_R_X75Y122_SLICE_X115Y122_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y122_SLICE_X115Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y122_SLICE_X115Y122_DO5),
.O6(CLBLL_R_X75Y122_SLICE_X115Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y122_SLICE_X115Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y122_SLICE_X115Y122_CO5),
.O6(CLBLL_R_X75Y122_SLICE_X115Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hacffac00acffac00)
  ) CLBLL_R_X75Y122_SLICE_X115Y122_BLUT (
.I0(CLBLL_R_X79Y127_SLICE_X122Y127_BQ),
.I1(CLBLL_R_X75Y122_SLICE_X115Y122_BQ),
.I2(CLBLL_R_X75Y123_SLICE_X114Y123_AO6),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X76Y122_SLICE_X116Y122_AQ),
.I5(1'b1),
.O5(CLBLL_R_X75Y122_SLICE_X115Y122_BO5),
.O6(CLBLL_R_X75Y122_SLICE_X115Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h50505050cceecc44)
  ) CLBLL_R_X75Y122_SLICE_X115Y122_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X75Y122_SLICE_X115Y122_BQ),
.I2(CLBLM_L_X74Y121_SLICE_X113Y121_AQ),
.I3(CLBLL_R_X75Y123_SLICE_X114Y123_AO6),
.I4(CLBLL_R_X75Y122_SLICE_X115Y122_A5Q),
.I5(1'b1),
.O5(CLBLL_R_X75Y122_SLICE_X115Y122_AO5),
.O6(CLBLL_R_X75Y122_SLICE_X115Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y123_SLICE_X114Y123_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y123_SLICE_X114Y123_BO6),
.Q(CLBLL_R_X75Y123_SLICE_X114Y123_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y123_SLICE_X114Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y123_SLICE_X114Y123_DO5),
.O6(CLBLL_R_X75Y123_SLICE_X114Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLL_R_X75Y123_SLICE_X114Y123_CLUT (
.I0(CLBLL_R_X75Y113_SLICE_X114Y113_AQ),
.I1(CLBLM_L_X76Y123_SLICE_X117Y123_AQ),
.I2(CLBLM_L_X74Y123_SLICE_X113Y123_BQ),
.I3(CLBLL_R_X75Y123_SLICE_X114Y123_BQ),
.I4(CLBLM_L_X74Y123_SLICE_X113Y123_A5Q),
.I5(CLBLM_L_X74Y123_SLICE_X113Y123_DQ),
.O5(CLBLL_R_X75Y123_SLICE_X114Y123_CO5),
.O6(CLBLL_R_X75Y123_SLICE_X114Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h06006666f0f0f0f0)
  ) CLBLL_R_X75Y123_SLICE_X114Y123_BLUT (
.I0(CLBLM_L_X74Y123_SLICE_X113Y123_CO5),
.I1(CLBLL_R_X75Y123_SLICE_X114Y123_BQ),
.I2(CLBLM_L_X76Y123_SLICE_X116Y123_BQ),
.I3(CLBLL_R_X75Y121_SLICE_X114Y121_BQ),
.I4(CLBLL_R_X75Y123_SLICE_X115Y123_AQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLL_R_X75Y123_SLICE_X114Y123_BO5),
.O6(CLBLL_R_X75Y123_SLICE_X114Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000a00080000000)
  ) CLBLL_R_X75Y123_SLICE_X114Y123_ALUT (
.I0(CLBLM_L_X74Y123_SLICE_X113Y123_A5Q),
.I1(CLBLL_R_X75Y123_SLICE_X114Y123_BQ),
.I2(CLBLL_R_X75Y113_SLICE_X114Y113_AQ),
.I3(CLBLM_L_X76Y123_SLICE_X117Y123_AQ),
.I4(CLBLM_L_X74Y123_SLICE_X113Y123_BQ),
.I5(1'b1),
.O5(CLBLL_R_X75Y123_SLICE_X114Y123_AO5),
.O6(CLBLL_R_X75Y123_SLICE_X114Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y123_SLICE_X115Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y123_SLICE_X116Y123_DO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y124_SLICE_X115Y124_B5Q),
.Q(CLBLL_R_X75Y123_SLICE_X115Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4400440044004400)
  ) CLBLL_R_X75Y123_SLICE_X115Y123_DLUT (
.I0(CLBLL_R_X77Y123_SLICE_X119Y123_AQ),
.I1(CLBLM_L_X78Y124_SLICE_X120Y124_CQ),
.I2(1'b1),
.I3(CLBLM_L_X76Y123_SLICE_X116Y123_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y123_SLICE_X115Y123_DO5),
.O6(CLBLL_R_X75Y123_SLICE_X115Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5050000050400000)
  ) CLBLL_R_X75Y123_SLICE_X115Y123_CLUT (
.I0(CLBLL_R_X77Y123_SLICE_X119Y123_AQ),
.I1(CLBLM_L_X76Y122_SLICE_X116Y122_A5Q),
.I2(CLBLM_L_X78Y124_SLICE_X120Y124_CQ),
.I3(CLBLM_L_X76Y122_SLICE_X116Y122_AQ),
.I4(CLBLM_L_X76Y123_SLICE_X116Y123_A5Q),
.I5(CLBLM_L_X76Y122_SLICE_X116Y122_BQ),
.O5(CLBLL_R_X75Y123_SLICE_X115Y123_CO5),
.O6(CLBLL_R_X75Y123_SLICE_X115Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff7fffffffffff)
  ) CLBLL_R_X75Y123_SLICE_X115Y123_BLUT (
.I0(CLBLM_L_X76Y123_SLICE_X116Y123_A5Q),
.I1(CLBLM_L_X76Y125_SLICE_X117Y125_AQ),
.I2(CLBLL_R_X75Y124_SLICE_X114Y124_AQ),
.I3(CLBLL_R_X75Y124_SLICE_X114Y124_BQ),
.I4(CLBLL_R_X77Y123_SLICE_X119Y123_AQ),
.I5(CLBLM_L_X78Y124_SLICE_X120Y124_CQ),
.O5(CLBLL_R_X75Y123_SLICE_X115Y123_BO5),
.O6(CLBLL_R_X75Y123_SLICE_X115Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800aaaabfffbfff)
  ) CLBLL_R_X75Y123_SLICE_X115Y123_ALUT (
.I0(CLBLM_L_X76Y123_SLICE_X117Y123_AQ),
.I1(CLBLM_L_X74Y109_SLICE_X113Y109_AQ),
.I2(CLBLM_L_X74Y123_SLICE_X113Y123_BQ),
.I3(CLBLM_L_X74Y123_SLICE_X113Y123_A5Q),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLL_R_X75Y123_SLICE_X115Y123_AO5),
.O6(CLBLL_R_X75Y123_SLICE_X115Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y124_SLICE_X114Y124_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y124_SLICE_X114Y124_CO5),
.Q(CLBLL_R_X75Y124_SLICE_X114Y124_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y124_SLICE_X114Y124_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y124_SLICE_X114Y124_DO5),
.Q(CLBLL_R_X75Y124_SLICE_X114Y124_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y124_SLICE_X114Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y124_SLICE_X114Y124_AO6),
.Q(CLBLL_R_X75Y124_SLICE_X114Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y124_SLICE_X114Y124_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y124_SLICE_X114Y124_BO6),
.Q(CLBLL_R_X75Y124_SLICE_X114Y124_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y124_SLICE_X114Y124_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y124_SLICE_X114Y124_CO6),
.Q(CLBLL_R_X75Y124_SLICE_X114Y124_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y124_SLICE_X114Y124_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y124_SLICE_X114Y124_DO6),
.Q(CLBLL_R_X75Y124_SLICE_X114Y124_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff0f0efe0efe0)
  ) CLBLL_R_X75Y124_SLICE_X114Y124_DLUT (
.I0(CLBLM_L_X74Y123_SLICE_X112Y123_BQ),
.I1(CLBLL_R_X75Y124_SLICE_X114Y124_D5Q),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X76Y123_SLICE_X117Y123_CQ),
.I4(CLBLL_R_X75Y121_SLICE_X114Y121_AQ),
.I5(1'b1),
.O5(CLBLL_R_X75Y124_SLICE_X114Y124_DO5),
.O6(CLBLL_R_X75Y124_SLICE_X114Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff0f0aaffcccc)
  ) CLBLL_R_X75Y124_SLICE_X114Y124_CLUT (
.I0(CLBLL_R_X75Y124_SLICE_X114Y124_C5Q),
.I1(CLBLL_R_X75Y124_SLICE_X114Y124_D5Q),
.I2(CLBLL_R_X75Y124_SLICE_X114Y124_DQ),
.I3(CLBLM_L_X76Y118_SLICE_X117Y118_CQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLL_R_X75Y124_SLICE_X114Y124_CO5),
.O6(CLBLL_R_X75Y124_SLICE_X114Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5577008855dd0088)
  ) CLBLL_R_X75Y124_SLICE_X114Y124_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X75Y124_SLICE_X114Y124_BQ),
.I2(1'b1),
.I3(CLBLL_R_X77Y122_SLICE_X118Y122_CO6),
.I4(CLBLM_L_X76Y125_SLICE_X117Y125_AQ),
.I5(CLBLL_R_X75Y123_SLICE_X115Y123_DO6),
.O5(CLBLL_R_X75Y124_SLICE_X114Y124_BO5),
.O6(CLBLL_R_X75Y124_SLICE_X114Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h557d00a055f500a0)
  ) CLBLL_R_X75Y124_SLICE_X114Y124_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X76Y125_SLICE_X117Y125_AQ),
.I2(CLBLL_R_X75Y124_SLICE_X114Y124_AQ),
.I3(CLBLL_R_X77Y122_SLICE_X118Y122_CO6),
.I4(CLBLL_R_X75Y124_SLICE_X114Y124_BQ),
.I5(CLBLL_R_X75Y123_SLICE_X115Y123_DO6),
.O5(CLBLL_R_X75Y124_SLICE_X114Y124_AO5),
.O6(CLBLL_R_X75Y124_SLICE_X114Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y124_SLICE_X115Y124_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y124_SLICE_X115Y124_BO5),
.Q(CLBLL_R_X75Y124_SLICE_X115Y124_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y124_SLICE_X115Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y124_SLICE_X115Y124_AO6),
.Q(CLBLL_R_X75Y124_SLICE_X115Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y124_SLICE_X115Y124_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y124_SLICE_X115Y124_BO6),
.Q(CLBLL_R_X75Y124_SLICE_X115Y124_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y124_SLICE_X115Y124_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y124_SLICE_X115Y124_CO6),
.Q(CLBLL_R_X75Y124_SLICE_X115Y124_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y124_SLICE_X115Y124_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y124_SLICE_X115Y124_DO6),
.Q(CLBLL_R_X75Y124_SLICE_X115Y124_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbfb7373c8c84040)
  ) CLBLL_R_X75Y124_SLICE_X115Y124_DLUT (
.I0(CLBLM_L_X74Y123_SLICE_X113Y123_CO5),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLL_R_X75Y124_SLICE_X115Y124_DQ),
.I3(1'b1),
.I4(CLBLL_R_X79Y127_SLICE_X122Y127_BQ),
.I5(CLBLM_L_X76Y124_SLICE_X116Y124_CQ),
.O5(CLBLL_R_X75Y124_SLICE_X115Y124_DO5),
.O6(CLBLL_R_X75Y124_SLICE_X115Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeef0f04444f0f0)
  ) CLBLL_R_X75Y124_SLICE_X115Y124_CLUT (
.I0(CLBLM_L_X74Y123_SLICE_X113Y123_CO5),
.I1(CLBLL_R_X75Y124_SLICE_X115Y124_CQ),
.I2(CLBLM_L_X76Y124_SLICE_X116Y124_A5Q),
.I3(1'b1),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X79Y127_SLICE_X122Y127_CQ),
.O5(CLBLL_R_X75Y124_SLICE_X115Y124_CO5),
.O6(CLBLL_R_X75Y124_SLICE_X115Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ccccf5550000)
  ) CLBLL_R_X75Y124_SLICE_X115Y124_BLUT (
.I0(CLBLM_L_X76Y124_SLICE_X116Y124_CO6),
.I1(CLBLL_R_X75Y124_SLICE_X114Y124_CQ),
.I2(CLBLL_R_X75Y124_SLICE_X115Y124_B5Q),
.I3(CLBLL_R_X75Y123_SLICE_X115Y123_AO5),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLL_R_X75Y124_SLICE_X115Y124_BO5),
.O6(CLBLL_R_X75Y124_SLICE_X115Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h30ffb8ff3000b800)
  ) CLBLL_R_X75Y124_SLICE_X115Y124_ALUT (
.I0(CLBLL_R_X75Y124_SLICE_X115Y124_B5Q),
.I1(CLBLM_L_X74Y123_SLICE_X113Y123_CO5),
.I2(CLBLL_R_X75Y124_SLICE_X115Y124_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLL_R_X75Y122_SLICE_X114Y122_AQ),
.I5(CLBLM_L_X76Y124_SLICE_X116Y124_AQ),
.O5(CLBLL_R_X75Y124_SLICE_X115Y124_AO5),
.O6(CLBLL_R_X75Y124_SLICE_X115Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y127_SLICE_X114Y127_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y127_SLICE_X114Y127_AO5),
.Q(CLBLL_R_X75Y127_SLICE_X114Y127_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y127_SLICE_X114Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y127_SLICE_X114Y127_AO6),
.Q(CLBLL_R_X75Y127_SLICE_X114Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y127_SLICE_X114Y127_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y127_SLICE_X114Y127_BO6),
.Q(CLBLL_R_X75Y127_SLICE_X114Y127_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y127_SLICE_X114Y127_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y127_SLICE_X114Y127_DO6),
.Q(CLBLL_R_X75Y127_SLICE_X114Y127_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f1f0e0ffff0000)
  ) CLBLL_R_X75Y127_SLICE_X114Y127_DLUT (
.I0(CLBLL_R_X75Y127_SLICE_X114Y127_A5Q),
.I1(CLBLL_R_X75Y127_SLICE_X114Y127_AQ),
.I2(CLBLL_R_X75Y127_SLICE_X114Y127_DQ),
.I3(CLBLL_R_X75Y128_SLICE_X115Y128_CO6),
.I4(CLBLL_R_X75Y128_SLICE_X114Y128_CQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLL_R_X75Y127_SLICE_X114Y127_DO5),
.O6(CLBLL_R_X75Y127_SLICE_X114Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaffaadddddddd)
  ) CLBLL_R_X75Y127_SLICE_X114Y127_CLUT (
.I0(CLBLL_R_X75Y127_SLICE_X114Y127_A5Q),
.I1(CLBLL_R_X73Y127_SLICE_X110Y127_A5Q),
.I2(1'b1),
.I3(CLBLL_R_X75Y128_SLICE_X115Y128_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y127_SLICE_X114Y127_CO5),
.O6(CLBLL_R_X75Y127_SLICE_X114Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8888fd5da808)
  ) CLBLL_R_X75Y127_SLICE_X114Y127_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X75Y127_SLICE_X114Y127_BQ),
.I2(CLBLL_R_X73Y127_SLICE_X110Y127_A5Q),
.I3(CLBLL_R_X75Y128_SLICE_X114Y128_BO6),
.I4(CLBLL_R_X73Y127_SLICE_X111Y127_AQ),
.I5(CLBLL_R_X75Y127_SLICE_X114Y127_CO6),
.O5(CLBLL_R_X75Y127_SLICE_X114Y127_BO5),
.O6(CLBLL_R_X75Y127_SLICE_X114Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a02022dd88ff00)
  ) CLBLL_R_X75Y127_SLICE_X114Y127_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X75Y127_SLICE_X114Y127_A5Q),
.I2(CLBLL_R_X75Y127_SLICE_X114Y127_AQ),
.I3(CLBLL_R_X73Y127_SLICE_X110Y127_A5Q),
.I4(CLBLL_R_X75Y128_SLICE_X115Y128_CO6),
.I5(1'b1),
.O5(CLBLL_R_X75Y127_SLICE_X114Y127_AO5),
.O6(CLBLL_R_X75Y127_SLICE_X114Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y127_SLICE_X115Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y127_SLICE_X115Y127_AO6),
.Q(CLBLL_R_X75Y127_SLICE_X115Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y127_SLICE_X115Y127_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y127_SLICE_X115Y127_BO6),
.Q(CLBLL_R_X75Y127_SLICE_X115Y127_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y127_SLICE_X115Y127_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y127_SLICE_X115Y127_CO6),
.Q(CLBLL_R_X75Y127_SLICE_X115Y127_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y127_SLICE_X115Y127_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y127_SLICE_X115Y127_DO6),
.Q(CLBLL_R_X75Y127_SLICE_X115Y127_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0a5cccccccc)
  ) CLBLL_R_X75Y127_SLICE_X115Y127_DLUT (
.I0(CLBLM_L_X74Y129_SLICE_X112Y129_AQ),
.I1(CLBLL_R_X75Y127_SLICE_X115Y127_CQ),
.I2(CLBLL_R_X75Y127_SLICE_X115Y127_DQ),
.I3(CLBLM_L_X74Y129_SLICE_X112Y129_A5Q),
.I4(CLBLL_R_X75Y128_SLICE_X115Y128_DO6),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLL_R_X75Y127_SLICE_X115Y127_DO5),
.O6(CLBLL_R_X75Y127_SLICE_X115Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa5acacaaa5acaca)
  ) CLBLL_R_X75Y127_SLICE_X115Y127_CLUT (
.I0(CLBLL_R_X75Y127_SLICE_X115Y127_BQ),
.I1(CLBLL_R_X75Y127_SLICE_X115Y127_CQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X72Y127_SLICE_X108Y127_DQ),
.I4(CLBLM_L_X74Y128_SLICE_X113Y128_BO5),
.I5(1'b1),
.O5(CLBLL_R_X75Y127_SLICE_X115Y127_CO5),
.O6(CLBLL_R_X75Y127_SLICE_X115Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccdffffccc80000)
  ) CLBLL_R_X75Y127_SLICE_X115Y127_BLUT (
.I0(CLBLL_R_X75Y128_SLICE_X115Y128_DO6),
.I1(CLBLL_R_X75Y127_SLICE_X115Y127_BQ),
.I2(CLBLM_L_X74Y129_SLICE_X112Y129_AQ),
.I3(CLBLM_L_X74Y129_SLICE_X112Y129_A5Q),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X72Y127_SLICE_X108Y127_DQ),
.O5(CLBLL_R_X75Y127_SLICE_X115Y127_BO5),
.O6(CLBLL_R_X75Y127_SLICE_X115Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0100000001000100)
  ) CLBLL_R_X75Y127_SLICE_X115Y127_ALUT (
.I0(CLBLM_L_X60Y104_SLICE_X90Y104_AQ),
.I1(CLBLM_L_X62Y105_SLICE_X93Y105_A5Q),
.I2(CLBLL_R_X75Y127_SLICE_X115Y127_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLL_R_X77Y130_SLICE_X118Y130_DO5),
.I5(CLBLM_L_X76Y128_SLICE_X117Y128_CO6),
.O5(CLBLL_R_X75Y127_SLICE_X115Y127_AO5),
.O6(CLBLL_R_X75Y127_SLICE_X115Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y128_SLICE_X114Y128_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y128_SLICE_X114Y128_CO6),
.Q(CLBLL_R_X75Y128_SLICE_X114Y128_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfffcfffcfcffff)
  ) CLBLL_R_X75Y128_SLICE_X114Y128_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X74Y129_SLICE_X113Y129_CO6),
.I2(CLBLM_L_X76Y130_SLICE_X116Y130_AQ),
.I3(CLBLM_L_X76Y128_SLICE_X116Y128_A5Q),
.I4(CLBLL_R_X77Y128_SLICE_X118Y128_B5Q),
.I5(1'b1),
.O5(CLBLL_R_X75Y128_SLICE_X114Y128_DO5),
.O6(CLBLL_R_X75Y128_SLICE_X114Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hca3acacaca7aca8a)
  ) CLBLL_R_X75Y128_SLICE_X114Y128_CLUT (
.I0(CLBLL_R_X75Y127_SLICE_X114Y127_A5Q),
.I1(CLBLL_R_X75Y128_SLICE_X114Y128_CQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLL_R_X75Y128_SLICE_X115Y128_CO6),
.I4(CLBLL_R_X75Y128_SLICE_X114Y128_BO5),
.I5(CLBLL_R_X75Y127_SLICE_X114Y127_AQ),
.O5(CLBLL_R_X75Y128_SLICE_X114Y128_CO5),
.O6(CLBLL_R_X75Y128_SLICE_X114Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcfffcfefefefe)
  ) CLBLL_R_X75Y128_SLICE_X114Y128_BLUT (
.I0(CLBLL_R_X77Y128_SLICE_X118Y128_B5Q),
.I1(CLBLL_R_X75Y129_SLICE_X114Y129_BQ),
.I2(CLBLM_L_X74Y129_SLICE_X113Y129_CO6),
.I3(CLBLM_L_X76Y128_SLICE_X116Y128_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y128_SLICE_X114Y128_BO5),
.O6(CLBLL_R_X75Y128_SLICE_X114Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffafffaffddffdd)
  ) CLBLL_R_X75Y128_SLICE_X114Y128_ALUT (
.I0(CLBLM_L_X76Y128_SLICE_X116Y128_A5Q),
.I1(CLBLL_R_X75Y130_SLICE_X115Y130_AQ),
.I2(CLBLL_R_X75Y129_SLICE_X114Y129_DQ),
.I3(CLBLM_L_X74Y129_SLICE_X113Y129_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y128_SLICE_X114Y128_AO5),
.O6(CLBLL_R_X75Y128_SLICE_X114Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h222222222a222222)
  ) CLBLL_R_X75Y128_SLICE_X115Y128_DLUT (
.I0(CLBLL_R_X75Y130_SLICE_X114Y130_BO6),
.I1(CLBLL_R_X77Y126_SLICE_X118Y126_AQ),
.I2(CLBLL_R_X77Y129_SLICE_X118Y129_CQ),
.I3(CLBLM_L_X76Y128_SLICE_X116Y128_DO6),
.I4(CLBLM_L_X76Y128_SLICE_X117Y128_B5Q),
.I5(CLBLL_R_X77Y128_SLICE_X118Y128_CQ),
.O5(CLBLL_R_X75Y128_SLICE_X115Y128_DO5),
.O6(CLBLL_R_X75Y128_SLICE_X115Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb030303030303030)
  ) CLBLL_R_X75Y128_SLICE_X115Y128_CLUT (
.I0(CLBLL_R_X77Y129_SLICE_X118Y129_CQ),
.I1(CLBLM_L_X62Y105_SLICE_X93Y105_A5Q),
.I2(CLBLL_R_X75Y129_SLICE_X115Y129_DO6),
.I3(CLBLM_L_X76Y128_SLICE_X116Y128_DO6),
.I4(CLBLM_L_X76Y128_SLICE_X117Y128_B5Q),
.I5(CLBLL_R_X77Y128_SLICE_X118Y128_CQ),
.O5(CLBLL_R_X75Y128_SLICE_X115Y128_CO5),
.O6(CLBLL_R_X75Y128_SLICE_X115Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0080ffff00000000)
  ) CLBLL_R_X75Y128_SLICE_X115Y128_BLUT (
.I0(CLBLM_L_X76Y128_SLICE_X116Y128_DO6),
.I1(CLBLL_R_X77Y128_SLICE_X118Y128_CQ),
.I2(CLBLM_L_X76Y128_SLICE_X117Y128_B5Q),
.I3(CLBLL_R_X77Y129_SLICE_X118Y129_CQ),
.I4(CLBLM_L_X60Y104_SLICE_X90Y104_AQ),
.I5(CLBLL_R_X75Y129_SLICE_X115Y129_CO6),
.O5(CLBLL_R_X75Y128_SLICE_X115Y128_BO5),
.O6(CLBLL_R_X75Y128_SLICE_X115Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2000aaaa0000aaaa)
  ) CLBLL_R_X75Y128_SLICE_X115Y128_ALUT (
.I0(CLBLL_R_X75Y129_SLICE_X115Y129_BO6),
.I1(CLBLL_R_X77Y128_SLICE_X118Y128_CQ),
.I2(CLBLM_L_X76Y128_SLICE_X117Y128_B5Q),
.I3(CLBLL_R_X77Y129_SLICE_X118Y129_CQ),
.I4(CLBLL_R_X75Y127_SLICE_X115Y127_AQ),
.I5(CLBLM_L_X76Y128_SLICE_X116Y128_DO6),
.O5(CLBLL_R_X75Y128_SLICE_X115Y128_AO5),
.O6(CLBLL_R_X75Y128_SLICE_X115Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y129_SLICE_X114Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y129_SLICE_X114Y129_AO6),
.Q(CLBLL_R_X75Y129_SLICE_X114Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y129_SLICE_X114Y129_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y129_SLICE_X114Y129_BO6),
.Q(CLBLL_R_X75Y129_SLICE_X114Y129_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y129_SLICE_X114Y129_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y129_SLICE_X114Y129_DO6),
.Q(CLBLL_R_X75Y129_SLICE_X114Y129_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0cc78ccf0ccf0cc)
  ) CLBLL_R_X75Y129_SLICE_X114Y129_DLUT (
.I0(CLBLL_R_X75Y129_SLICE_X114Y129_CO5),
.I1(CLBLL_R_X75Y129_SLICE_X114Y129_AQ),
.I2(CLBLL_R_X75Y129_SLICE_X114Y129_DQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLL_R_X75Y130_SLICE_X114Y130_AQ),
.I5(CLBLM_L_X76Y130_SLICE_X116Y130_BQ),
.O5(CLBLL_R_X75Y129_SLICE_X114Y129_DO5),
.O6(CLBLL_R_X75Y129_SLICE_X114Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0000050500000)
  ) CLBLL_R_X75Y129_SLICE_X114Y129_CLUT (
.I0(CLBLL_R_X77Y128_SLICE_X118Y128_CQ),
.I1(1'b1),
.I2(CLBLL_R_X77Y129_SLICE_X118Y129_CQ),
.I3(1'b1),
.I4(CLBLM_L_X76Y127_SLICE_X116Y127_AQ),
.I5(1'b1),
.O5(CLBLL_R_X75Y129_SLICE_X114Y129_CO5),
.O6(CLBLL_R_X75Y129_SLICE_X114Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd7dd8888dddd8888)
  ) CLBLL_R_X75Y129_SLICE_X114Y129_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X75Y129_SLICE_X114Y129_BQ),
.I2(CLBLL_R_X75Y130_SLICE_X114Y130_AQ),
.I3(CLBLM_L_X76Y130_SLICE_X116Y130_BQ),
.I4(CLBLL_R_X75Y129_SLICE_X115Y129_AQ),
.I5(CLBLL_R_X75Y129_SLICE_X114Y129_CO6),
.O5(CLBLL_R_X75Y129_SLICE_X114Y129_BO5),
.O6(CLBLL_R_X75Y129_SLICE_X114Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7373f3f34044c0c0)
  ) CLBLL_R_X75Y129_SLICE_X114Y129_ALUT (
.I0(CLBLL_R_X75Y130_SLICE_X114Y130_CO6),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLL_R_X75Y129_SLICE_X114Y129_AQ),
.I3(CLBLM_L_X76Y130_SLICE_X116Y130_A5Q),
.I4(CLBLL_R_X75Y129_SLICE_X114Y129_CO5),
.I5(CLBLM_L_X76Y130_SLICE_X116Y130_BQ),
.O5(CLBLL_R_X75Y129_SLICE_X114Y129_AO5),
.O6(CLBLL_R_X75Y129_SLICE_X114Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y129_SLICE_X115Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y129_SLICE_X115Y129_AO6),
.Q(CLBLL_R_X75Y129_SLICE_X115Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000c000800)
  ) CLBLL_R_X75Y129_SLICE_X115Y129_DLUT (
.I0(CLBLM_L_X78Y131_SLICE_X120Y131_AQ),
.I1(CLBLM_L_X76Y125_SLICE_X117Y125_BQ),
.I2(CLBLM_L_X76Y130_SLICE_X116Y130_DQ),
.I3(CLBLL_R_X77Y129_SLICE_X119Y129_BQ),
.I4(CLBLL_R_X77Y130_SLICE_X118Y130_AQ),
.I5(CLBLL_R_X75Y129_SLICE_X114Y129_BQ),
.O5(CLBLL_R_X75Y129_SLICE_X115Y129_DO5),
.O6(CLBLL_R_X75Y129_SLICE_X115Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0404040000000000)
  ) CLBLL_R_X75Y129_SLICE_X115Y129_CLUT (
.I0(CLBLL_R_X75Y130_SLICE_X115Y130_AQ),
.I1(CLBLL_R_X77Y129_SLICE_X119Y129_BQ),
.I2(CLBLM_L_X76Y130_SLICE_X116Y130_DQ),
.I3(CLBLM_L_X78Y131_SLICE_X120Y131_AQ),
.I4(CLBLL_R_X77Y130_SLICE_X118Y130_AQ),
.I5(CLBLM_L_X76Y125_SLICE_X117Y125_BQ),
.O5(CLBLL_R_X75Y129_SLICE_X115Y129_CO5),
.O6(CLBLL_R_X75Y129_SLICE_X115Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0030002000000000)
  ) CLBLL_R_X75Y129_SLICE_X115Y129_BLUT (
.I0(CLBLL_R_X77Y130_SLICE_X118Y130_AQ),
.I1(CLBLM_L_X76Y130_SLICE_X116Y130_DQ),
.I2(CLBLM_L_X76Y125_SLICE_X117Y125_BQ),
.I3(CLBLL_R_X75Y129_SLICE_X114Y129_DQ),
.I4(CLBLM_L_X78Y131_SLICE_X120Y131_AQ),
.I5(CLBLL_R_X77Y129_SLICE_X119Y129_BQ),
.O5(CLBLL_R_X75Y129_SLICE_X115Y129_BO5),
.O6(CLBLL_R_X75Y129_SLICE_X115Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50ccccf050cccc)
  ) CLBLL_R_X75Y129_SLICE_X115Y129_ALUT (
.I0(CLBLL_R_X75Y129_SLICE_X114Y129_CO6),
.I1(CLBLL_R_X75Y130_SLICE_X115Y130_AQ),
.I2(CLBLL_R_X75Y129_SLICE_X115Y129_AQ),
.I3(CLBLM_L_X76Y129_SLICE_X116Y129_AO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X76Y130_SLICE_X116Y130_CO6),
.O5(CLBLL_R_X75Y129_SLICE_X115Y129_AO5),
.O6(CLBLL_R_X75Y129_SLICE_X115Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y130_SLICE_X114Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y130_SLICE_X114Y130_AO6),
.Q(CLBLL_R_X75Y130_SLICE_X114Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h99cc99cc99cccccc)
  ) CLBLL_R_X75Y130_SLICE_X114Y130_DLUT (
.I0(CLBLM_L_X76Y128_SLICE_X117Y128_AQ),
.I1(CLBLL_R_X75Y130_SLICE_X115Y130_AQ),
.I2(1'b1),
.I3(CLBLL_R_X77Y129_SLICE_X119Y129_BQ),
.I4(CLBLM_L_X78Y131_SLICE_X120Y131_AQ),
.I5(CLBLL_R_X77Y130_SLICE_X118Y130_AQ),
.O5(CLBLL_R_X75Y130_SLICE_X114Y130_DO5),
.O6(CLBLL_R_X75Y130_SLICE_X114Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a0f5a0f5a0f0f0f)
  ) CLBLL_R_X75Y130_SLICE_X114Y130_CLUT (
.I0(CLBLM_L_X76Y128_SLICE_X117Y128_AQ),
.I1(1'b1),
.I2(CLBLL_R_X75Y129_SLICE_X114Y129_DQ),
.I3(CLBLL_R_X77Y129_SLICE_X119Y129_BQ),
.I4(CLBLM_L_X78Y131_SLICE_X120Y131_AQ),
.I5(CLBLL_R_X77Y130_SLICE_X118Y130_AQ),
.O5(CLBLL_R_X75Y130_SLICE_X114Y130_CO5),
.O6(CLBLL_R_X75Y130_SLICE_X114Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0300020000000000)
  ) CLBLL_R_X75Y130_SLICE_X114Y130_BLUT (
.I0(CLBLM_L_X78Y131_SLICE_X120Y131_AQ),
.I1(CLBLM_L_X76Y130_SLICE_X116Y130_AQ),
.I2(CLBLM_L_X76Y130_SLICE_X116Y130_DQ),
.I3(CLBLM_L_X76Y125_SLICE_X117Y125_BQ),
.I4(CLBLL_R_X77Y130_SLICE_X118Y130_AQ),
.I5(CLBLL_R_X77Y129_SLICE_X119Y129_BQ),
.O5(CLBLL_R_X75Y130_SLICE_X114Y130_BO5),
.O6(CLBLL_R_X75Y130_SLICE_X114Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f780f5a0f5a0)
  ) CLBLL_R_X75Y130_SLICE_X114Y130_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X77Y129_SLICE_X118Y129_CQ),
.I2(CLBLL_R_X75Y130_SLICE_X114Y130_AQ),
.I3(CLBLM_L_X76Y130_SLICE_X116Y130_A5Q),
.I4(CLBLL_R_X77Y128_SLICE_X118Y128_CQ),
.I5(CLBLM_L_X76Y127_SLICE_X116Y127_AQ),
.O5(CLBLL_R_X75Y130_SLICE_X114Y130_AO5),
.O6(CLBLL_R_X75Y130_SLICE_X114Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y130_SLICE_X115Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y130_SLICE_X115Y130_AO6),
.Q(CLBLL_R_X75Y130_SLICE_X115Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y130_SLICE_X115Y130_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y130_SLICE_X115Y130_CO6),
.Q(CLBLL_R_X75Y130_SLICE_X115Y130_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y130_SLICE_X115Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y130_SLICE_X115Y130_DO5),
.O6(CLBLL_R_X75Y130_SLICE_X115Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5d5a080dddd8888)
  ) CLBLL_R_X75Y130_SLICE_X115Y130_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X75Y130_SLICE_X115Y130_CQ),
.I2(CLBLL_R_X75Y130_SLICE_X114Y130_DO6),
.I3(CLBLM_L_X76Y130_SLICE_X116Y130_CO6),
.I4(CLBLL_R_X75Y129_SLICE_X114Y129_DQ),
.I5(CLBLL_R_X75Y130_SLICE_X115Y130_BO6),
.O5(CLBLL_R_X75Y130_SLICE_X115Y130_CO5),
.O6(CLBLL_R_X75Y130_SLICE_X115Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000c0c000003030)
  ) CLBLL_R_X75Y130_SLICE_X115Y130_BLUT (
.I0(1'b1),
.I1(CLBLL_R_X77Y128_SLICE_X118Y128_CQ),
.I2(CLBLM_L_X76Y127_SLICE_X116Y127_AQ),
.I3(1'b1),
.I4(CLBLL_R_X77Y129_SLICE_X118Y129_CQ),
.I5(1'b1),
.O5(CLBLL_R_X75Y130_SLICE_X115Y130_BO5),
.O6(CLBLL_R_X75Y130_SLICE_X115Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e26ae2e2e2e2e2)
  ) CLBLL_R_X75Y130_SLICE_X115Y130_ALUT (
.I0(CLBLL_R_X75Y130_SLICE_X115Y130_CQ),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLL_R_X75Y130_SLICE_X115Y130_AQ),
.I3(CLBLL_R_X75Y130_SLICE_X115Y130_BO6),
.I4(CLBLL_R_X75Y130_SLICE_X114Y130_AQ),
.I5(CLBLM_L_X76Y130_SLICE_X116Y130_BQ),
.O5(CLBLL_R_X75Y130_SLICE_X115Y130_AO5),
.O6(CLBLL_R_X75Y130_SLICE_X115Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y133_SLICE_X114Y133_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y133_SLICE_X114Y133_AO6),
.Q(CLBLL_R_X75Y133_SLICE_X114Y133_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y133_SLICE_X114Y133_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y133_SLICE_X114Y133_BO6),
.Q(CLBLL_R_X75Y133_SLICE_X114Y133_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010100000800)
  ) CLBLL_R_X75Y133_SLICE_X114Y133_DLUT (
.I0(CLBLM_L_X74Y131_SLICE_X112Y131_AQ),
.I1(CLBLM_L_X74Y132_SLICE_X112Y132_C5Q),
.I2(CLBLL_R_X75Y133_SLICE_X115Y133_AQ),
.I3(CLBLL_R_X75Y134_SLICE_X115Y134_AQ),
.I4(CLBLM_L_X76Y133_SLICE_X116Y133_BQ),
.I5(CLBLL_R_X75Y133_SLICE_X115Y133_BQ),
.O5(CLBLL_R_X75Y133_SLICE_X114Y133_DO5),
.O6(CLBLL_R_X75Y133_SLICE_X114Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00050005ccc8ccc8)
  ) CLBLL_R_X75Y133_SLICE_X114Y133_CLUT (
.I0(CLBLL_R_X75Y133_SLICE_X114Y133_BQ),
.I1(CLBLM_L_X70Y136_SLICE_X105Y136_A5Q),
.I2(CLBLL_R_X75Y133_SLICE_X114Y133_AQ),
.I3(CLBLL_R_X75Y134_SLICE_X115Y134_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y133_SLICE_X114Y133_CO5),
.O6(CLBLL_R_X75Y133_SLICE_X114Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa99f0f0aaaaf0f0)
  ) CLBLL_R_X75Y133_SLICE_X114Y133_BLUT (
.I0(CLBLL_R_X75Y133_SLICE_X114Y133_DO6),
.I1(CLBLM_L_X74Y129_SLICE_X112Y129_BQ),
.I2(CLBLM_L_X74Y132_SLICE_X112Y132_C5Q),
.I3(CLBLL_R_X79Y135_SLICE_X122Y135_AQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X75Y133_SLICE_X114Y133_CO6),
.O5(CLBLL_R_X75Y133_SLICE_X114Y133_BO5),
.O6(CLBLL_R_X75Y133_SLICE_X114Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff7fbfff00004000)
  ) CLBLL_R_X75Y133_SLICE_X114Y133_ALUT (
.I0(CLBLM_L_X74Y132_SLICE_X112Y132_C5Q),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLL_R_X75Y133_SLICE_X115Y133_AO6),
.I3(CLBLL_R_X75Y133_SLICE_X115Y133_BQ),
.I4(CLBLM_L_X74Y131_SLICE_X112Y131_AQ),
.I5(CLBLL_R_X75Y134_SLICE_X115Y134_AQ),
.O5(CLBLL_R_X75Y133_SLICE_X114Y133_AO5),
.O6(CLBLL_R_X75Y133_SLICE_X114Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y133_SLICE_X115Y133_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y133_SLICE_X115Y133_AO5),
.Q(CLBLL_R_X75Y133_SLICE_X115Y133_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y133_SLICE_X115Y133_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y129_SLICE_X112Y129_BQ),
.Q(CLBLL_R_X75Y133_SLICE_X115Y133_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y133_SLICE_X115Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y133_SLICE_X115Y133_DO5),
.O6(CLBLL_R_X75Y133_SLICE_X115Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y133_SLICE_X115Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y133_SLICE_X115Y133_CO5),
.O6(CLBLL_R_X75Y133_SLICE_X115Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y133_SLICE_X115Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y133_SLICE_X115Y133_BO5),
.O6(CLBLL_R_X75Y133_SLICE_X115Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000f0ffd55a800)
  ) CLBLL_R_X75Y133_SLICE_X115Y133_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X75Y134_SLICE_X114Y134_CO5),
.I2(CLBLL_R_X75Y133_SLICE_X115Y133_AQ),
.I3(CLBLL_R_X75Y134_SLICE_X115Y134_BO6),
.I4(CLBLM_L_X76Y133_SLICE_X116Y133_BQ),
.I5(1'b1),
.O5(CLBLL_R_X75Y133_SLICE_X115Y133_AO5),
.O6(CLBLL_R_X75Y133_SLICE_X115Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y134_SLICE_X114Y134_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y134_SLICE_X114Y134_BO6),
.Q(CLBLL_R_X75Y134_SLICE_X114Y134_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y134_SLICE_X114Y134_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y134_SLICE_X114Y134_AO6),
.Q(CLBLL_R_X75Y134_SLICE_X114Y134_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f3f3ffffffff)
  ) CLBLL_R_X75Y134_SLICE_X114Y134_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X74Y134_SLICE_X112Y134_BQ),
.I2(CLBLM_L_X74Y134_SLICE_X112Y134_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X74Y132_SLICE_X112Y132_C5Q),
.O5(CLBLL_R_X75Y134_SLICE_X114Y134_DO5),
.O6(CLBLL_R_X75Y134_SLICE_X114Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000040a44aa44aa)
  ) CLBLL_R_X75Y134_SLICE_X114Y134_CLUT (
.I0(CLBLL_R_X75Y133_SLICE_X115Y133_BQ),
.I1(CLBLL_R_X75Y134_SLICE_X115Y134_AQ),
.I2(CLBLM_L_X76Y133_SLICE_X116Y133_BQ),
.I3(CLBLM_L_X74Y132_SLICE_X112Y132_C5Q),
.I4(CLBLL_R_X75Y133_SLICE_X115Y133_AQ),
.I5(1'b1),
.O5(CLBLL_R_X75Y134_SLICE_X114Y134_CO5),
.O6(CLBLL_R_X75Y134_SLICE_X114Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7830b8b855005500)
  ) CLBLL_R_X75Y134_SLICE_X114Y134_BLUT (
.I0(CLBLL_R_X75Y134_SLICE_X114Y134_A5Q),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLL_R_X75Y134_SLICE_X114Y134_AQ),
.I3(CLBLL_R_X75Y133_SLICE_X115Y133_AQ),
.I4(CLBLL_R_X75Y134_SLICE_X114Y134_CO5),
.I5(1'b1),
.O5(CLBLL_R_X75Y134_SLICE_X114Y134_BO5),
.O6(CLBLL_R_X75Y134_SLICE_X114Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f0cf3c03300f3c0)
  ) CLBLL_R_X75Y134_SLICE_X114Y134_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLL_R_X75Y134_SLICE_X114Y134_AQ),
.I3(CLBLM_L_X76Y134_SLICE_X117Y134_BQ),
.I4(CLBLL_R_X75Y134_SLICE_X114Y134_CO5),
.I5(CLBLL_R_X75Y133_SLICE_X115Y133_AQ),
.O5(CLBLL_R_X75Y134_SLICE_X114Y134_AO5),
.O6(CLBLL_R_X75Y134_SLICE_X114Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X75Y134_SLICE_X115Y134_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X79Y135_SLICE_X122Y135_AQ),
.Q(CLBLL_R_X75Y134_SLICE_X115Y134_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0000000ff)
  ) CLBLL_R_X75Y134_SLICE_X115Y134_DLUT (
.I0(CLBLM_L_X76Y134_SLICE_X116Y134_AQ),
.I1(1'b1),
.I2(CLBLM_L_X76Y134_SLICE_X117Y134_AQ),
.I3(CLBLL_R_X75Y133_SLICE_X115Y133_BQ),
.I4(CLBLL_R_X75Y134_SLICE_X115Y134_AQ),
.I5(1'b1),
.O5(CLBLL_R_X75Y134_SLICE_X115Y134_DO5),
.O6(CLBLL_R_X75Y134_SLICE_X115Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a08080a0a080a)
  ) CLBLL_R_X75Y134_SLICE_X115Y134_CLUT (
.I0(CLBLL_R_X75Y133_SLICE_X114Y133_BQ),
.I1(CLBLL_R_X75Y133_SLICE_X115Y133_AQ),
.I2(CLBLL_R_X75Y134_SLICE_X114Y134_DO6),
.I3(CLBLL_R_X75Y134_SLICE_X115Y134_AO5),
.I4(CLBLM_L_X76Y133_SLICE_X116Y133_BQ),
.I5(CLBLL_R_X75Y134_SLICE_X115Y134_DO5),
.O5(CLBLL_R_X75Y134_SLICE_X115Y134_CO5),
.O6(CLBLL_R_X75Y134_SLICE_X115Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5753f7f75707)
  ) CLBLL_R_X75Y134_SLICE_X115Y134_BLUT (
.I0(CLBLL_R_X75Y134_SLICE_X115Y134_DO6),
.I1(CLBLL_R_X75Y134_SLICE_X115Y134_AQ),
.I2(CLBLL_R_X75Y133_SLICE_X115Y133_BQ),
.I3(CLBLL_R_X75Y134_SLICE_X114Y134_BO5),
.I4(CLBLM_L_X76Y133_SLICE_X116Y133_BQ),
.I5(CLBLM_L_X74Y132_SLICE_X112Y132_C5Q),
.O5(CLBLL_R_X75Y134_SLICE_X115Y134_BO5),
.O6(CLBLL_R_X75Y134_SLICE_X115Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555aaaa7fffbfff)
  ) CLBLL_R_X75Y134_SLICE_X115Y134_ALUT (
.I0(CLBLL_R_X75Y133_SLICE_X115Y133_BQ),
.I1(CLBLM_L_X76Y134_SLICE_X117Y134_BQ),
.I2(CLBLM_L_X76Y133_SLICE_X116Y133_AQ),
.I3(CLBLM_L_X76Y134_SLICE_X116Y134_BQ),
.I4(CLBLM_L_X74Y132_SLICE_X112Y132_C5Q),
.I5(1'b1),
.O5(CLBLL_R_X75Y134_SLICE_X115Y134_AO5),
.O6(CLBLL_R_X75Y134_SLICE_X115Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y104_SLICE_X118Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y104_SLICE_X118Y104_BQ),
.Q(CLBLL_R_X77Y104_SLICE_X118Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y104_SLICE_X118Y104_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y104_SLICE_X118Y104_CQ),
.Q(CLBLL_R_X77Y104_SLICE_X118Y104_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y104_SLICE_X118Y104_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y104_SLICE_X119Y104_AQ),
.Q(CLBLL_R_X77Y104_SLICE_X118Y104_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y104_SLICE_X118Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y104_SLICE_X118Y104_DO5),
.O6(CLBLL_R_X77Y104_SLICE_X118Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y104_SLICE_X118Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y104_SLICE_X118Y104_CO5),
.O6(CLBLL_R_X77Y104_SLICE_X118Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y104_SLICE_X118Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y104_SLICE_X118Y104_BO5),
.O6(CLBLL_R_X77Y104_SLICE_X118Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y104_SLICE_X118Y104_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y104_SLICE_X118Y104_AO5),
.O6(CLBLL_R_X77Y104_SLICE_X118Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y104_SLICE_X119Y104_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y104_SLICE_X119Y104_AO5),
.Q(CLBLL_R_X77Y104_SLICE_X119Y104_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y104_SLICE_X119Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y104_SLICE_X119Y104_AO6),
.Q(CLBLL_R_X77Y104_SLICE_X119Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y104_SLICE_X119Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y104_SLICE_X119Y104_DO5),
.O6(CLBLL_R_X77Y104_SLICE_X119Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y104_SLICE_X119Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y104_SLICE_X119Y104_CO5),
.O6(CLBLL_R_X77Y104_SLICE_X119Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y104_SLICE_X119Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y104_SLICE_X119Y104_BO5),
.O6(CLBLL_R_X77Y104_SLICE_X119Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfffc00aa00aa00)
  ) CLBLL_R_X77Y104_SLICE_X119Y104_ALUT (
.I0(CLBLM_L_X64Y106_SLICE_X97Y106_AQ),
.I1(CLBLL_R_X79Y104_SLICE_X122Y104_BQ),
.I2(CLBLL_R_X77Y104_SLICE_X119Y104_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X78Y104_SLICE_X120Y104_BQ),
.I5(1'b1),
.O5(CLBLL_R_X77Y104_SLICE_X119Y104_AO5),
.O6(CLBLL_R_X77Y104_SLICE_X119Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y108_SLICE_X118Y108_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y100_SLICE_X106Y100_BQ),
.Q(CLBLL_R_X77Y108_SLICE_X118Y108_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y108_SLICE_X118Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y108_SLICE_X118Y108_DO5),
.O6(CLBLL_R_X77Y108_SLICE_X118Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y108_SLICE_X118Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y108_SLICE_X118Y108_CO5),
.O6(CLBLL_R_X77Y108_SLICE_X118Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y108_SLICE_X118Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y108_SLICE_X118Y108_BO5),
.O6(CLBLL_R_X77Y108_SLICE_X118Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y108_SLICE_X118Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y108_SLICE_X118Y108_AO5),
.O6(CLBLL_R_X77Y108_SLICE_X118Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y108_SLICE_X119Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y108_SLICE_X119Y108_DO5),
.O6(CLBLL_R_X77Y108_SLICE_X119Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y108_SLICE_X119Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y108_SLICE_X119Y108_CO5),
.O6(CLBLL_R_X77Y108_SLICE_X119Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y108_SLICE_X119Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y108_SLICE_X119Y108_BO5),
.O6(CLBLL_R_X77Y108_SLICE_X119Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y108_SLICE_X119Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y108_SLICE_X119Y108_AO5),
.O6(CLBLL_R_X77Y108_SLICE_X119Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y113_SLICE_X118Y113_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y111_SLICE_X108Y111_C5Q),
.Q(CLBLL_R_X77Y113_SLICE_X118Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y113_SLICE_X118Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y113_SLICE_X118Y113_DO5),
.O6(CLBLL_R_X77Y113_SLICE_X118Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y113_SLICE_X118Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y113_SLICE_X118Y113_CO5),
.O6(CLBLL_R_X77Y113_SLICE_X118Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y113_SLICE_X118Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y113_SLICE_X118Y113_BO5),
.O6(CLBLL_R_X77Y113_SLICE_X118Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y113_SLICE_X118Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y113_SLICE_X118Y113_AO5),
.O6(CLBLL_R_X77Y113_SLICE_X118Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y113_SLICE_X119Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y113_SLICE_X119Y113_DO5),
.O6(CLBLL_R_X77Y113_SLICE_X119Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y113_SLICE_X119Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y113_SLICE_X119Y113_CO5),
.O6(CLBLL_R_X77Y113_SLICE_X119Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y113_SLICE_X119Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y113_SLICE_X119Y113_BO5),
.O6(CLBLL_R_X77Y113_SLICE_X119Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y113_SLICE_X119Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y113_SLICE_X119Y113_AO5),
.O6(CLBLL_R_X77Y113_SLICE_X119Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y121_SLICE_X118Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y121_SLICE_X118Y121_DO5),
.O6(CLBLL_R_X77Y121_SLICE_X118Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y121_SLICE_X118Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y121_SLICE_X118Y121_CO5),
.O6(CLBLL_R_X77Y121_SLICE_X118Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y121_SLICE_X118Y121_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y121_SLICE_X118Y121_BO5),
.O6(CLBLL_R_X77Y121_SLICE_X118Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeaacc00aabb0033)
  ) CLBLL_R_X77Y121_SLICE_X118Y121_ALUT (
.I0(CLBLL_R_X77Y121_SLICE_X119Y121_DQ),
.I1(CLBLM_L_X76Y118_SLICE_X116Y118_DQ),
.I2(1'b1),
.I3(CLBLM_L_X78Y123_SLICE_X121Y123_A5Q),
.I4(CLBLL_R_X77Y121_SLICE_X119Y121_AQ),
.I5(CLBLM_L_X76Y118_SLICE_X116Y118_AQ),
.O5(CLBLL_R_X77Y121_SLICE_X118Y121_AO5),
.O6(CLBLL_R_X77Y121_SLICE_X118Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y121_SLICE_X119Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y121_SLICE_X119Y121_AO6),
.Q(CLBLL_R_X77Y121_SLICE_X119Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y121_SLICE_X119Y121_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y121_SLICE_X119Y121_CO6),
.Q(CLBLL_R_X77Y121_SLICE_X119Y121_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y121_SLICE_X119Y121_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y121_SLICE_X119Y121_DO6),
.Q(CLBLL_R_X77Y121_SLICE_X119Y121_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h50505014cccccccc)
  ) CLBLL_R_X77Y121_SLICE_X119Y121_DLUT (
.I0(CLBLM_L_X78Y123_SLICE_X121Y123_CO6),
.I1(CLBLL_R_X77Y121_SLICE_X119Y121_CQ),
.I2(CLBLL_R_X77Y121_SLICE_X119Y121_DQ),
.I3(CLBLM_L_X78Y122_SLICE_X120Y122_DO6),
.I4(CLBLL_R_X77Y121_SLICE_X119Y121_BO5),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLL_R_X77Y121_SLICE_X119Y121_DO5),
.O6(CLBLL_R_X77Y121_SLICE_X119Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h44441444f0f0f0f0)
  ) CLBLL_R_X77Y121_SLICE_X119Y121_CLUT (
.I0(CLBLM_L_X78Y123_SLICE_X121Y123_CO6),
.I1(CLBLL_R_X77Y121_SLICE_X119Y121_CQ),
.I2(CLBLL_R_X77Y122_SLICE_X119Y122_DQ),
.I3(CLBLL_R_X77Y122_SLICE_X119Y122_CQ),
.I4(CLBLM_L_X78Y122_SLICE_X120Y122_DO6),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLL_R_X77Y121_SLICE_X119Y121_CO5),
.O6(CLBLL_R_X77Y121_SLICE_X119Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0303055ffddff)
  ) CLBLL_R_X77Y121_SLICE_X119Y121_BLUT (
.I0(CLBLL_R_X77Y122_SLICE_X119Y122_DQ),
.I1(CLBLL_R_X77Y113_SLICE_X118Y113_AQ),
.I2(CLBLL_R_X77Y121_SLICE_X119Y121_AQ),
.I3(CLBLL_R_X77Y122_SLICE_X119Y122_CQ),
.I4(CLBLM_L_X76Y122_SLICE_X117Y122_AQ),
.I5(1'b1),
.O5(CLBLL_R_X77Y121_SLICE_X119Y121_BO5),
.O6(CLBLL_R_X77Y121_SLICE_X119Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ff000ff1ff000)
  ) CLBLL_R_X77Y121_SLICE_X119Y121_ALUT (
.I0(CLBLL_R_X77Y121_SLICE_X119Y121_BO5),
.I1(CLBLL_R_X77Y122_SLICE_X119Y122_AO6),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLL_R_X77Y121_SLICE_X119Y121_BO6),
.I4(CLBLL_R_X77Y121_SLICE_X119Y121_DQ),
.I5(CLBLM_L_X78Y122_SLICE_X120Y122_DO6),
.O5(CLBLL_R_X77Y121_SLICE_X119Y121_AO5),
.O6(CLBLL_R_X77Y121_SLICE_X119Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y122_SLICE_X118Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y122_SLICE_X118Y122_AO6),
.Q(CLBLL_R_X77Y122_SLICE_X118Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y122_SLICE_X118Y122_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y122_SLICE_X118Y122_BO6),
.Q(CLBLL_R_X77Y122_SLICE_X118Y122_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y122_SLICE_X118Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y122_SLICE_X118Y122_DO5),
.O6(CLBLL_R_X77Y122_SLICE_X118Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00ff44ff)
  ) CLBLL_R_X77Y122_SLICE_X118Y122_CLUT (
.I0(CLBLL_R_X77Y121_SLICE_X118Y121_AO6),
.I1(CLBLL_R_X75Y123_SLICE_X114Y123_AO6),
.I2(1'b1),
.I3(CLBLM_L_X76Y125_SLICE_X117Y125_BQ),
.I4(CLBLM_L_X78Y123_SLICE_X120Y123_DO6),
.I5(CLBLL_R_X75Y123_SLICE_X115Y123_CO6),
.O5(CLBLL_R_X77Y122_SLICE_X118Y122_CO5),
.O6(CLBLL_R_X77Y122_SLICE_X118Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88cc283cf0f0f0f0)
  ) CLBLL_R_X77Y122_SLICE_X118Y122_BLUT (
.I0(CLBLM_L_X76Y122_SLICE_X117Y122_AQ),
.I1(CLBLL_R_X77Y122_SLICE_X118Y122_BQ),
.I2(CLBLL_R_X77Y122_SLICE_X118Y122_AQ),
.I3(CLBLL_R_X77Y113_SLICE_X118Y113_AQ),
.I4(CLBLM_L_X78Y122_SLICE_X120Y122_BO6),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLL_R_X77Y122_SLICE_X118Y122_BO5),
.O6(CLBLL_R_X77Y122_SLICE_X118Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h83c3ffff83c30000)
  ) CLBLL_R_X77Y122_SLICE_X118Y122_ALUT (
.I0(CLBLM_L_X76Y122_SLICE_X117Y122_AQ),
.I1(CLBLM_L_X78Y122_SLICE_X120Y122_BO6),
.I2(CLBLL_R_X77Y122_SLICE_X118Y122_AQ),
.I3(CLBLL_R_X77Y113_SLICE_X118Y113_AQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X78Y122_SLICE_X121Y122_BQ),
.O5(CLBLL_R_X77Y122_SLICE_X118Y122_AO5),
.O6(CLBLL_R_X77Y122_SLICE_X118Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y122_SLICE_X119Y122_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y122_SLICE_X119Y122_BO6),
.Q(CLBLL_R_X77Y122_SLICE_X119Y122_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y122_SLICE_X119Y122_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y122_SLICE_X119Y122_CO6),
.Q(CLBLL_R_X77Y122_SLICE_X119Y122_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y122_SLICE_X119Y122_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y122_SLICE_X119Y122_DO6),
.Q(CLBLL_R_X77Y122_SLICE_X119Y122_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa006acccccccc)
  ) CLBLL_R_X77Y122_SLICE_X119Y122_DLUT (
.I0(CLBLL_R_X77Y122_SLICE_X119Y122_DQ),
.I1(CLBLL_R_X77Y122_SLICE_X119Y122_CQ),
.I2(CLBLL_R_X77Y122_SLICE_X119Y122_BQ),
.I3(CLBLM_L_X78Y123_SLICE_X121Y123_CO6),
.I4(CLBLM_L_X78Y122_SLICE_X120Y122_CO6),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLL_R_X77Y122_SLICE_X119Y122_DO5),
.O6(CLBLL_R_X77Y122_SLICE_X119Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc4c433c4ff00ff00)
  ) CLBLL_R_X77Y122_SLICE_X119Y122_CLUT (
.I0(CLBLL_R_X77Y113_SLICE_X118Y113_AQ),
.I1(CLBLL_R_X77Y122_SLICE_X119Y122_CQ),
.I2(CLBLM_L_X76Y122_SLICE_X117Y122_AQ),
.I3(CLBLL_R_X77Y122_SLICE_X119Y122_BQ),
.I4(CLBLM_L_X78Y122_SLICE_X120Y122_CO6),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLL_R_X77Y122_SLICE_X119Y122_CO5),
.O6(CLBLL_R_X77Y122_SLICE_X119Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f000f00cfc06fc0)
  ) CLBLL_R_X77Y122_SLICE_X119Y122_BLUT (
.I0(CLBLL_R_X77Y122_SLICE_X118Y122_AQ),
.I1(CLBLL_R_X77Y122_SLICE_X119Y122_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLL_R_X77Y122_SLICE_X118Y122_BQ),
.I4(CLBLM_L_X78Y122_SLICE_X120Y122_BO6),
.I5(CLBLM_L_X78Y123_SLICE_X121Y123_CO6),
.O5(CLBLL_R_X77Y122_SLICE_X119Y122_BO5),
.O6(CLBLL_R_X77Y122_SLICE_X119Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0cffff5dff5dff)
  ) CLBLL_R_X77Y122_SLICE_X119Y122_ALUT (
.I0(CLBLL_R_X77Y122_SLICE_X118Y122_AQ),
.I1(CLBLL_R_X77Y113_SLICE_X118Y113_AQ),
.I2(CLBLM_L_X76Y122_SLICE_X117Y122_AQ),
.I3(CLBLL_R_X77Y122_SLICE_X118Y122_BQ),
.I4(CLBLL_R_X77Y121_SLICE_X119Y121_CQ),
.I5(1'b1),
.O5(CLBLL_R_X77Y122_SLICE_X119Y122_AO5),
.O6(CLBLL_R_X77Y122_SLICE_X119Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y123_SLICE_X118Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y123_SLICE_X118Y123_AO6),
.Q(CLBLL_R_X77Y123_SLICE_X118Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y123_SLICE_X118Y123_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y123_SLICE_X118Y123_CO6),
.Q(CLBLL_R_X77Y123_SLICE_X118Y123_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0200000000000000)
  ) CLBLL_R_X77Y123_SLICE_X118Y123_DLUT (
.I0(CLBLM_L_X78Y124_SLICE_X120Y124_BQ),
.I1(CLBLL_R_X77Y123_SLICE_X118Y123_CQ),
.I2(CLBLL_R_X77Y124_SLICE_X118Y124_BQ),
.I3(CLBLM_L_X78Y124_SLICE_X120Y124_AQ),
.I4(CLBLM_L_X74Y123_SLICE_X113Y123_CO5),
.I5(CLBLL_R_X77Y123_SLICE_X118Y123_AQ),
.O5(CLBLL_R_X77Y123_SLICE_X118Y123_DO5),
.O6(CLBLL_R_X77Y123_SLICE_X118Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8ddd8d8d8d8d8d8)
  ) CLBLL_R_X77Y123_SLICE_X118Y123_CLUT (
.I0(CLBLM_L_X76Y123_SLICE_X117Y123_AO5),
.I1(CLBLL_R_X77Y123_SLICE_X118Y123_CQ),
.I2(CLBLL_R_X77Y123_SLICE_X118Y123_AQ),
.I3(CLBLL_R_X77Y123_SLICE_X119Y123_CQ),
.I4(CLBLM_L_X76Y124_SLICE_X117Y124_BQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLL_R_X77Y123_SLICE_X118Y123_CO5),
.O6(CLBLL_R_X77Y123_SLICE_X118Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2020202000002000)
  ) CLBLL_R_X77Y123_SLICE_X118Y123_BLUT (
.I0(CLBLM_L_X76Y123_SLICE_X117Y123_AQ),
.I1(CLBLM_L_X74Y123_SLICE_X113Y123_A5Q),
.I2(CLBLL_R_X75Y113_SLICE_X114Y113_AQ),
.I3(CLBLM_L_X78Y124_SLICE_X120Y124_CQ),
.I4(CLBLL_R_X77Y123_SLICE_X119Y123_AQ),
.I5(1'b1),
.O5(CLBLL_R_X77Y123_SLICE_X118Y123_BO5),
.O6(CLBLL_R_X77Y123_SLICE_X118Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88c0c8c0ccc0ccc0)
  ) CLBLL_R_X77Y123_SLICE_X118Y123_ALUT (
.I0(CLBLL_R_X77Y124_SLICE_X118Y124_DO6),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLL_R_X77Y123_SLICE_X118Y123_AQ),
.I3(CLBLL_R_X77Y123_SLICE_X118Y123_BO6),
.I4(CLBLL_R_X77Y123_SLICE_X119Y123_AQ),
.I5(CLBLM_L_X78Y124_SLICE_X120Y124_CQ),
.O5(CLBLL_R_X77Y123_SLICE_X118Y123_AO5),
.O6(CLBLL_R_X77Y123_SLICE_X118Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y123_SLICE_X119Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y123_SLICE_X119Y123_AO6),
.Q(CLBLL_R_X77Y123_SLICE_X119Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y123_SLICE_X119Y123_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y123_SLICE_X119Y123_CO6),
.Q(CLBLL_R_X77Y123_SLICE_X119Y123_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00ff00fd00)
  ) CLBLL_R_X77Y123_SLICE_X119Y123_DLUT (
.I0(CLBLL_R_X75Y123_SLICE_X114Y123_AO6),
.I1(CLBLL_R_X77Y121_SLICE_X118Y121_AO6),
.I2(CLBLL_R_X77Y124_SLICE_X118Y124_AO5),
.I3(CLBLM_L_X76Y125_SLICE_X117Y125_BQ),
.I4(CLBLL_R_X77Y123_SLICE_X118Y123_AQ),
.I5(CLBLM_L_X78Y124_SLICE_X120Y124_CQ),
.O5(CLBLL_R_X77Y123_SLICE_X119Y123_DO5),
.O6(CLBLL_R_X77Y123_SLICE_X119Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefe5454eefe4454)
  ) CLBLL_R_X77Y123_SLICE_X119Y123_CLUT (
.I0(CLBLM_L_X76Y123_SLICE_X117Y123_AO5),
.I1(CLBLM_L_X76Y125_SLICE_X117Y125_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLL_R_X75Y122_SLICE_X114Y122_AQ),
.I4(CLBLL_R_X77Y123_SLICE_X119Y123_CQ),
.I5(CLBLM_L_X76Y119_SLICE_X116Y119_BO6),
.O5(CLBLL_R_X77Y123_SLICE_X119Y123_CO5),
.O6(CLBLL_R_X77Y123_SLICE_X119Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaaaaffffffef)
  ) CLBLL_R_X77Y123_SLICE_X119Y123_BLUT (
.I0(CLBLM_L_X78Y124_SLICE_X120Y124_CQ),
.I1(CLBLL_R_X77Y124_SLICE_X118Y124_AO5),
.I2(CLBLL_R_X75Y123_SLICE_X114Y123_AO6),
.I3(CLBLL_R_X77Y121_SLICE_X118Y121_AO6),
.I4(CLBLL_R_X77Y123_SLICE_X118Y123_AQ),
.I5(1'b1),
.O5(CLBLL_R_X77Y123_SLICE_X119Y123_BO5),
.O6(CLBLL_R_X77Y123_SLICE_X119Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0bbf0fff000f000)
  ) CLBLL_R_X77Y123_SLICE_X119Y123_ALUT (
.I0(CLBLL_R_X77Y123_SLICE_X119Y123_CQ),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLL_R_X77Y123_SLICE_X119Y123_AQ),
.I3(CLBLM_L_X76Y123_SLICE_X117Y123_AO5),
.I4(CLBLM_L_X76Y124_SLICE_X117Y124_BQ),
.I5(CLBLL_R_X77Y123_SLICE_X118Y123_CQ),
.O5(CLBLL_R_X77Y123_SLICE_X119Y123_AO5),
.O6(CLBLL_R_X77Y123_SLICE_X119Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y124_SLICE_X118Y124_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y124_SLICE_X118Y124_BO6),
.Q(CLBLL_R_X77Y124_SLICE_X118Y124_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00aa00aa00aa)
  ) CLBLL_R_X77Y124_SLICE_X118Y124_DLUT (
.I0(CLBLM_L_X76Y124_SLICE_X117Y124_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_R_X77Y123_SLICE_X119Y123_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y124_SLICE_X118Y124_DO5),
.O6(CLBLL_R_X77Y124_SLICE_X118Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000cc8000000000)
  ) CLBLL_R_X77Y124_SLICE_X118Y124_CLUT (
.I0(CLBLM_L_X78Y124_SLICE_X120Y124_BQ),
.I1(CLBLM_L_X78Y124_SLICE_X120Y124_CQ),
.I2(CLBLM_L_X78Y124_SLICE_X120Y124_AQ),
.I3(CLBLL_R_X77Y124_SLICE_X118Y124_BQ),
.I4(CLBLL_R_X77Y123_SLICE_X119Y123_AQ),
.I5(CLBLL_R_X77Y123_SLICE_X118Y123_BO6),
.O5(CLBLL_R_X77Y124_SLICE_X118Y124_CO5),
.O6(CLBLL_R_X77Y124_SLICE_X118Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33003300f3f0b3a0)
  ) CLBLL_R_X77Y124_SLICE_X118Y124_BLUT (
.I0(CLBLL_R_X77Y123_SLICE_X118Y123_BO5),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLL_R_X77Y126_SLICE_X118Y126_AO5),
.I3(CLBLM_L_X78Y124_SLICE_X120Y124_CQ),
.I4(CLBLL_R_X77Y124_SLICE_X118Y124_BQ),
.I5(CLBLL_R_X77Y124_SLICE_X118Y124_CO6),
.O5(CLBLL_R_X77Y124_SLICE_X118Y124_BO5),
.O6(CLBLL_R_X77Y124_SLICE_X118Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaa8affffffcc)
  ) CLBLL_R_X77Y124_SLICE_X118Y124_ALUT (
.I0(CLBLL_R_X77Y125_SLICE_X118Y125_CQ),
.I1(CLBLL_R_X77Y124_SLICE_X118Y124_BQ),
.I2(CLBLM_L_X76Y123_SLICE_X116Y123_AQ),
.I3(CLBLM_L_X78Y124_SLICE_X120Y124_AQ),
.I4(CLBLM_L_X78Y124_SLICE_X120Y124_BQ),
.I5(1'b1),
.O5(CLBLL_R_X77Y124_SLICE_X118Y124_AO5),
.O6(CLBLL_R_X77Y124_SLICE_X118Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y124_SLICE_X119Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y124_SLICE_X119Y124_AO6),
.Q(CLBLL_R_X77Y124_SLICE_X119Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y124_SLICE_X119Y124_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y124_SLICE_X119Y124_BO6),
.Q(CLBLL_R_X77Y124_SLICE_X119Y124_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y124_SLICE_X119Y124_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y124_SLICE_X119Y124_CO6),
.Q(CLBLL_R_X77Y124_SLICE_X119Y124_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha2a2a2a2a2a2a2a2)
  ) CLBLL_R_X77Y124_SLICE_X119Y124_DLUT (
.I0(CLBLL_R_X75Y122_SLICE_X114Y122_AQ),
.I1(CLBLL_R_X77Y123_SLICE_X118Y123_DO6),
.I2(CLBLM_L_X76Y119_SLICE_X116Y119_BO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y124_SLICE_X119Y124_DO5),
.O6(CLBLL_R_X77Y124_SLICE_X119Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6ccc0000f0f0f0f0)
  ) CLBLL_R_X77Y124_SLICE_X119Y124_CLUT (
.I0(CLBLL_R_X77Y123_SLICE_X118Y123_DO6),
.I1(CLBLL_R_X77Y124_SLICE_X119Y124_CQ),
.I2(CLBLL_R_X77Y124_SLICE_X119Y124_BQ),
.I3(CLBLL_R_X77Y124_SLICE_X119Y124_AQ),
.I4(CLBLL_R_X77Y124_SLICE_X119Y124_DO6),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLL_R_X77Y124_SLICE_X119Y124_CO5),
.O6(CLBLL_R_X77Y124_SLICE_X119Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h73aa00aa80aa00aa)
  ) CLBLL_R_X77Y124_SLICE_X119Y124_BLUT (
.I0(CLBLL_R_X77Y124_SLICE_X119Y124_AQ),
.I1(CLBLL_R_X77Y123_SLICE_X118Y123_DO6),
.I2(CLBLM_L_X76Y119_SLICE_X116Y119_BO6),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLL_R_X75Y122_SLICE_X114Y122_AQ),
.I5(CLBLL_R_X77Y124_SLICE_X119Y124_BQ),
.O5(CLBLL_R_X77Y124_SLICE_X119Y124_BO5),
.O6(CLBLL_R_X77Y124_SLICE_X119Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h66f022f000f000f0)
  ) CLBLL_R_X77Y124_SLICE_X119Y124_ALUT (
.I0(CLBLL_R_X77Y124_SLICE_X119Y124_AQ),
.I1(CLBLL_R_X77Y123_SLICE_X118Y123_DO6),
.I2(CLBLM_L_X76Y124_SLICE_X117Y124_BQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X76Y119_SLICE_X116Y119_BO6),
.I5(CLBLL_R_X75Y122_SLICE_X114Y122_AQ),
.O5(CLBLL_R_X77Y124_SLICE_X119Y124_AO5),
.O6(CLBLL_R_X77Y124_SLICE_X119Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y125_SLICE_X118Y125_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y125_SLICE_X118Y125_AO5),
.Q(CLBLL_R_X77Y125_SLICE_X118Y125_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y125_SLICE_X118Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y125_SLICE_X118Y125_AO6),
.Q(CLBLL_R_X77Y125_SLICE_X118Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y125_SLICE_X118Y125_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y125_SLICE_X118Y125_BO6),
.Q(CLBLL_R_X77Y125_SLICE_X118Y125_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y125_SLICE_X118Y125_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y125_SLICE_X118Y125_CO6),
.Q(CLBLL_R_X77Y125_SLICE_X118Y125_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y125_SLICE_X118Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y125_SLICE_X118Y125_DO5),
.O6(CLBLL_R_X77Y125_SLICE_X118Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ffffaaaaaaaa)
  ) CLBLL_R_X77Y125_SLICE_X118Y125_CLUT (
.I0(CLBLL_R_X77Y127_SLICE_X118Y127_AQ),
.I1(CLBLL_R_X77Y125_SLICE_X118Y125_CQ),
.I2(CLBLL_R_X77Y125_SLICE_X118Y125_BQ),
.I3(CLBLL_R_X77Y125_SLICE_X118Y125_A5Q),
.I4(CLBLM_L_X76Y125_SLICE_X117Y125_CO6),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLL_R_X77Y125_SLICE_X118Y125_CO5),
.O6(CLBLL_R_X77Y125_SLICE_X118Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aaccaaffffdddd)
  ) CLBLL_R_X77Y125_SLICE_X118Y125_BLUT (
.I0(CLBLL_R_X77Y125_SLICE_X118Y125_CQ),
.I1(CLBLL_R_X77Y125_SLICE_X118Y125_BQ),
.I2(1'b1),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLL_R_X77Y125_SLICE_X118Y125_A5Q),
.I5(1'b1),
.O5(CLBLL_R_X77Y125_SLICE_X118Y125_BO5),
.O6(CLBLL_R_X77Y125_SLICE_X118Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00000099cc99cc)
  ) CLBLL_R_X77Y125_SLICE_X118Y125_ALUT (
.I0(CLBLL_R_X77Y125_SLICE_X118Y125_CQ),
.I1(CLBLL_R_X77Y125_SLICE_X118Y125_BQ),
.I2(1'b1),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_R_X67Y116_SLICE_X100Y116_AQ),
.I5(1'b1),
.O5(CLBLL_R_X77Y125_SLICE_X118Y125_AO5),
.O6(CLBLL_R_X77Y125_SLICE_X118Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y125_SLICE_X119Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y125_SLICE_X119Y125_DO5),
.O6(CLBLL_R_X77Y125_SLICE_X119Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y125_SLICE_X119Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y125_SLICE_X119Y125_CO5),
.O6(CLBLL_R_X77Y125_SLICE_X119Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y125_SLICE_X119Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y125_SLICE_X119Y125_BO5),
.O6(CLBLL_R_X77Y125_SLICE_X119Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y125_SLICE_X119Y125_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y125_SLICE_X119Y125_AO5),
.O6(CLBLL_R_X77Y125_SLICE_X119Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y126_SLICE_X118Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y105_SLICE_X93Y105_A5Q),
.Q(CLBLL_R_X77Y126_SLICE_X118Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y126_SLICE_X118Y126_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y126_SLICE_X118Y126_AO6),
.Q(CLBLL_R_X77Y126_SLICE_X118Y126_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y126_SLICE_X118Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y126_SLICE_X118Y126_DO5),
.O6(CLBLL_R_X77Y126_SLICE_X118Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y126_SLICE_X118Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y126_SLICE_X118Y126_CO5),
.O6(CLBLL_R_X77Y126_SLICE_X118Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y126_SLICE_X118Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y126_SLICE_X118Y126_BO5),
.O6(CLBLL_R_X77Y126_SLICE_X118Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cf03cf0aa00ff00)
  ) CLBLL_R_X77Y126_SLICE_X118Y126_ALUT (
.I0(CLBLL_R_X77Y123_SLICE_X119Y123_CQ),
.I1(CLBLL_R_X77Y126_SLICE_X118Y126_BQ),
.I2(CLBLL_R_X77Y126_SLICE_X118Y126_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X76Y124_SLICE_X117Y124_BQ),
.I5(1'b1),
.O5(CLBLL_R_X77Y126_SLICE_X118Y126_AO5),
.O6(CLBLL_R_X77Y126_SLICE_X118Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y126_SLICE_X119Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y126_SLICE_X119Y126_DO5),
.O6(CLBLL_R_X77Y126_SLICE_X119Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y126_SLICE_X119Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y126_SLICE_X119Y126_CO5),
.O6(CLBLL_R_X77Y126_SLICE_X119Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y126_SLICE_X119Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y126_SLICE_X119Y126_BO5),
.O6(CLBLL_R_X77Y126_SLICE_X119Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y126_SLICE_X119Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y126_SLICE_X119Y126_AO5),
.O6(CLBLL_R_X77Y126_SLICE_X119Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y127_SLICE_X118Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y127_SLICE_X118Y127_AO6),
.Q(CLBLL_R_X77Y127_SLICE_X118Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y127_SLICE_X118Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y127_SLICE_X118Y127_DO5),
.O6(CLBLL_R_X77Y127_SLICE_X118Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y127_SLICE_X118Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y127_SLICE_X118Y127_CO5),
.O6(CLBLL_R_X77Y127_SLICE_X118Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y127_SLICE_X118Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y127_SLICE_X118Y127_BO5),
.O6(CLBLL_R_X77Y127_SLICE_X118Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5fff500a0ffa000)
  ) CLBLL_R_X77Y127_SLICE_X118Y127_ALUT (
.I0(CLBLL_R_X77Y125_SLICE_X118Y125_BO5),
.I1(1'b1),
.I2(CLBLL_R_X77Y127_SLICE_X118Y127_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLL_R_X79Y127_SLICE_X122Y127_BQ),
.I5(CLBLL_R_X79Y127_SLICE_X122Y127_A5Q),
.O5(CLBLL_R_X77Y127_SLICE_X118Y127_AO5),
.O6(CLBLL_R_X77Y127_SLICE_X118Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y127_SLICE_X119Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y127_SLICE_X119Y127_AO6),
.Q(CLBLL_R_X77Y127_SLICE_X119Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y127_SLICE_X119Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y127_SLICE_X119Y127_DO5),
.O6(CLBLL_R_X77Y127_SLICE_X119Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y127_SLICE_X119Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y127_SLICE_X119Y127_CO5),
.O6(CLBLL_R_X77Y127_SLICE_X119Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y127_SLICE_X119Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y127_SLICE_X119Y127_BO5),
.O6(CLBLL_R_X77Y127_SLICE_X119Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000550000008c00)
  ) CLBLL_R_X77Y127_SLICE_X119Y127_ALUT (
.I0(CLBLM_L_X78Y127_SLICE_X121Y127_CO6),
.I1(CLBLL_R_X77Y123_SLICE_X119Y123_DO6),
.I2(CLBLL_R_X77Y127_SLICE_X119Y127_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X78Y127_SLICE_X121Y127_BO6),
.I5(1'b1),
.O5(CLBLL_R_X77Y127_SLICE_X119Y127_AO5),
.O6(CLBLL_R_X77Y127_SLICE_X119Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y128_SLICE_X118Y128_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y128_SLICE_X118Y128_BO5),
.Q(CLBLL_R_X77Y128_SLICE_X118Y128_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y128_SLICE_X118Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y127_SLICE_X116Y127_AQ),
.Q(CLBLL_R_X77Y128_SLICE_X118Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y128_SLICE_X118Y128_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y128_SLICE_X118Y128_BO6),
.Q(CLBLL_R_X77Y128_SLICE_X118Y128_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y128_SLICE_X118Y128_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y128_SLICE_X118Y128_AO5),
.Q(CLBLL_R_X77Y128_SLICE_X118Y128_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y128_SLICE_X118Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y128_SLICE_X118Y128_DO5),
.O6(CLBLL_R_X77Y128_SLICE_X118Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0e0f0e000110011)
  ) CLBLL_R_X77Y128_SLICE_X118Y128_CLUT (
.I0(CLBLL_R_X77Y129_SLICE_X118Y129_AQ),
.I1(CLBLL_R_X77Y128_SLICE_X119Y128_BQ),
.I2(CLBLM_L_X76Y128_SLICE_X116Y128_CQ),
.I3(CLBLL_R_X77Y130_SLICE_X119Y130_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y128_SLICE_X118Y128_CO5),
.O6(CLBLL_R_X77Y128_SLICE_X118Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccf0ccaaccaa)
  ) CLBLL_R_X77Y128_SLICE_X118Y128_BLUT (
.I0(CLBLM_L_X76Y128_SLICE_X116Y128_A5Q),
.I1(CLBLM_L_X76Y128_SLICE_X116Y128_CQ),
.I2(CLBLL_R_X77Y128_SLICE_X119Y128_A5Q),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y128_SLICE_X118Y128_BO5),
.O6(CLBLL_R_X77Y128_SLICE_X118Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a05cfca0fc)
  ) CLBLL_R_X77Y128_SLICE_X118Y128_ALUT (
.I0(CLBLL_R_X77Y128_SLICE_X119Y128_BQ),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLL_R_X77Y129_SLICE_X118Y129_CQ),
.I3(CLBLL_R_X77Y129_SLICE_X119Y129_AO6),
.I4(CLBLL_R_X77Y128_SLICE_X118Y128_CQ),
.I5(1'b1),
.O5(CLBLL_R_X77Y128_SLICE_X118Y128_AO5),
.O6(CLBLL_R_X77Y128_SLICE_X118Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y128_SLICE_X119Y128_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y128_SLICE_X119Y128_DQ),
.Q(CLBLL_R_X77Y128_SLICE_X119Y128_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y128_SLICE_X119Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y128_SLICE_X119Y128_AO6),
.Q(CLBLL_R_X77Y128_SLICE_X119Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y128_SLICE_X119Y128_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y128_SLICE_X119Y128_BO6),
.Q(CLBLL_R_X77Y128_SLICE_X119Y128_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y128_SLICE_X119Y128_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y128_SLICE_X119Y128_CO6),
.Q(CLBLL_R_X77Y128_SLICE_X119Y128_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y128_SLICE_X119Y128_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y128_SLICE_X119Y128_DO6),
.Q(CLBLL_R_X77Y128_SLICE_X119Y128_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ee22f0f0f0f0)
  ) CLBLL_R_X77Y128_SLICE_X119Y128_DLUT (
.I0(CLBLL_R_X77Y128_SLICE_X119Y128_DQ),
.I1(CLBLM_L_X62Y105_SLICE_X93Y105_A5Q),
.I2(CLBLL_R_X77Y128_SLICE_X118Y128_B5Q),
.I3(CLBLM_L_X76Y128_SLICE_X116Y128_CQ),
.I4(1'b1),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLL_R_X77Y128_SLICE_X119Y128_DO5),
.O6(CLBLL_R_X77Y128_SLICE_X119Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacacacffff0000)
  ) CLBLL_R_X77Y128_SLICE_X119Y128_CLUT (
.I0(CLBLM_L_X78Y128_SLICE_X120Y128_AQ),
.I1(CLBLL_R_X77Y128_SLICE_X119Y128_CQ),
.I2(CLBLL_R_X77Y128_SLICE_X119Y128_BQ),
.I3(1'b1),
.I4(CLBLL_R_X77Y128_SLICE_X119Y128_AQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLL_R_X77Y128_SLICE_X119Y128_CO5),
.O6(CLBLL_R_X77Y128_SLICE_X119Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc3300bf8c7340)
  ) CLBLL_R_X77Y128_SLICE_X119Y128_BLUT (
.I0(CLBLM_L_X76Y127_SLICE_X116Y127_AQ),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLL_R_X77Y128_SLICE_X118Y128_CO5),
.I3(CLBLL_R_X77Y128_SLICE_X118Y128_BQ),
.I4(CLBLM_L_X78Y129_SLICE_X120Y129_AO6),
.I5(CLBLM_L_X80Y132_SLICE_X124Y132_AQ),
.O5(CLBLL_R_X77Y128_SLICE_X119Y128_BO5),
.O6(CLBLL_R_X77Y128_SLICE_X119Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0accccaaaacccc)
  ) CLBLL_R_X77Y128_SLICE_X119Y128_ALUT (
.I0(CLBLL_R_X77Y128_SLICE_X119Y128_AQ),
.I1(CLBLM_L_X78Y128_SLICE_X120Y128_AQ),
.I2(CLBLL_R_X77Y128_SLICE_X118Y128_AO6),
.I3(CLBLL_R_X77Y128_SLICE_X118Y128_BQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X77Y128_SLICE_X118Y128_CQ),
.O5(CLBLL_R_X77Y128_SLICE_X119Y128_AO5),
.O6(CLBLL_R_X77Y128_SLICE_X119Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y129_SLICE_X118Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y129_SLICE_X118Y129_AO6),
.Q(CLBLL_R_X77Y129_SLICE_X118Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y129_SLICE_X118Y129_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y129_SLICE_X118Y129_BO6),
.Q(CLBLL_R_X77Y129_SLICE_X118Y129_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y129_SLICE_X118Y129_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y129_SLICE_X118Y129_CO6),
.Q(CLBLL_R_X77Y129_SLICE_X118Y129_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y129_SLICE_X118Y129_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y129_SLICE_X118Y129_DO6),
.Q(CLBLL_R_X77Y129_SLICE_X118Y129_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5dd55dd50cc00cc0)
  ) CLBLL_R_X77Y129_SLICE_X118Y129_DLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X77Y129_SLICE_X119Y129_AO6),
.I2(CLBLL_R_X77Y129_SLICE_X118Y129_DQ),
.I3(CLBLL_R_X77Y129_SLICE_X119Y129_DO6),
.I4(1'b1),
.I5(CLBLL_R_X77Y129_SLICE_X119Y129_BQ),
.O5(CLBLL_R_X77Y129_SLICE_X118Y129_DO5),
.O6(CLBLL_R_X77Y129_SLICE_X118Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h76660000ff660000)
  ) CLBLL_R_X77Y129_SLICE_X118Y129_CLUT (
.I0(CLBLL_R_X77Y128_SLICE_X119Y128_BQ),
.I1(CLBLL_R_X77Y129_SLICE_X118Y129_CQ),
.I2(CLBLL_R_X77Y128_SLICE_X118Y128_CQ),
.I3(CLBLL_R_X77Y130_SLICE_X119Y130_CO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X77Y129_SLICE_X119Y129_BQ),
.O5(CLBLL_R_X77Y129_SLICE_X118Y129_CO5),
.O6(CLBLL_R_X77Y129_SLICE_X118Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2828f8f88888f8f8)
  ) CLBLL_R_X77Y129_SLICE_X118Y129_BLUT (
.I0(CLBLL_R_X77Y129_SLICE_X119Y129_AO6),
.I1(CLBLL_R_X77Y129_SLICE_X118Y129_BQ),
.I2(CLBLL_R_X77Y129_SLICE_X118Y129_DQ),
.I3(1'b1),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X77Y129_SLICE_X119Y129_DO6),
.O5(CLBLL_R_X77Y129_SLICE_X118Y129_BO5),
.O6(CLBLL_R_X77Y129_SLICE_X118Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7dfffff00200000)
  ) CLBLL_R_X77Y129_SLICE_X118Y129_ALUT (
.I0(CLBLL_R_X77Y130_SLICE_X118Y130_AO5),
.I1(CLBLL_R_X77Y128_SLICE_X119Y128_A5Q),
.I2(CLBLL_R_X77Y128_SLICE_X118Y128_AQ),
.I3(CLBLL_R_X77Y128_SLICE_X118Y128_BQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X77Y130_SLICE_X119Y130_AQ),
.O5(CLBLL_R_X77Y129_SLICE_X118Y129_AO5),
.O6(CLBLL_R_X77Y129_SLICE_X118Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y129_SLICE_X119Y129_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y129_SLICE_X119Y129_BO6),
.Q(CLBLL_R_X77Y129_SLICE_X119Y129_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h008a000000aa0000)
  ) CLBLL_R_X77Y129_SLICE_X119Y129_DLUT (
.I0(CLBLL_R_X77Y128_SLICE_X119Y128_BQ),
.I1(CLBLL_R_X77Y128_SLICE_X119Y128_CQ),
.I2(CLBLL_R_X77Y128_SLICE_X118Y128_BQ),
.I3(CLBLL_R_X77Y129_SLICE_X118Y129_CQ),
.I4(CLBLL_R_X77Y128_SLICE_X118Y128_CQ),
.I5(CLBLM_L_X78Y128_SLICE_X120Y128_AQ),
.O5(CLBLL_R_X77Y129_SLICE_X119Y129_DO5),
.O6(CLBLL_R_X77Y129_SLICE_X119Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd0000000f0000000)
  ) CLBLL_R_X77Y129_SLICE_X119Y129_CLUT (
.I0(CLBLM_L_X78Y128_SLICE_X120Y128_AQ),
.I1(CLBLL_R_X77Y128_SLICE_X119Y128_CQ),
.I2(CLBLL_R_X77Y128_SLICE_X119Y128_BQ),
.I3(CLBLL_R_X77Y129_SLICE_X119Y129_AO5),
.I4(CLBLL_R_X77Y129_SLICE_X118Y129_DQ),
.I5(CLBLL_R_X77Y128_SLICE_X118Y128_BQ),
.O5(CLBLL_R_X77Y129_SLICE_X119Y129_CO5),
.O6(CLBLL_R_X77Y129_SLICE_X119Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2fefefef20e0e0e0)
  ) CLBLL_R_X77Y129_SLICE_X119Y129_BLUT (
.I0(CLBLL_R_X77Y130_SLICE_X119Y130_CO6),
.I1(CLBLL_R_X77Y129_SLICE_X119Y129_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLL_R_X77Y129_SLICE_X118Y129_BQ),
.I4(CLBLL_R_X77Y129_SLICE_X119Y129_CO6),
.I5(CLBLL_R_X77Y128_SLICE_X119Y128_CQ),
.O5(CLBLL_R_X77Y129_SLICE_X119Y129_BO5),
.O6(CLBLL_R_X77Y129_SLICE_X119Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd0d050d00000ff00)
  ) CLBLL_R_X77Y129_SLICE_X119Y129_ALUT (
.I0(CLBLL_R_X77Y130_SLICE_X119Y130_CO6),
.I1(CLBLL_R_X77Y129_SLICE_X119Y129_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLL_R_X77Y128_SLICE_X118Y128_CQ),
.I4(CLBLL_R_X77Y129_SLICE_X118Y129_CQ),
.I5(1'b1),
.O5(CLBLL_R_X77Y129_SLICE_X119Y129_AO5),
.O6(CLBLL_R_X77Y129_SLICE_X119Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y130_SLICE_X118Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y130_SLICE_X118Y130_AO6),
.Q(CLBLL_R_X77Y130_SLICE_X118Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y130_SLICE_X118Y130_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y130_SLICE_X118Y130_BO5),
.Q(CLBLL_R_X77Y130_SLICE_X118Y130_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y130_SLICE_X118Y130_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y130_SLICE_X118Y130_CO6),
.Q(CLBLL_R_X77Y130_SLICE_X118Y130_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555888800050008)
  ) CLBLL_R_X77Y130_SLICE_X118Y130_DLUT (
.I0(CLBLL_R_X77Y128_SLICE_X118Y128_BQ),
.I1(CLBLL_R_X77Y130_SLICE_X119Y130_AQ),
.I2(CLBLM_L_X78Y131_SLICE_X120Y131_AQ),
.I3(CLBLL_R_X77Y130_SLICE_X118Y130_AQ),
.I4(CLBLL_R_X77Y128_SLICE_X118Y128_AQ),
.I5(1'b1),
.O5(CLBLL_R_X77Y130_SLICE_X118Y130_DO5),
.O6(CLBLL_R_X77Y130_SLICE_X118Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7272d8d85050d8d8)
  ) CLBLL_R_X77Y130_SLICE_X118Y130_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X77Y130_SLICE_X118Y130_CQ),
.I2(CLBLL_R_X77Y131_SLICE_X119Y131_BQ),
.I3(1'b1),
.I4(CLBLL_R_X77Y130_SLICE_X118Y130_DO6),
.I5(CLBLL_R_X77Y130_SLICE_X118Y130_AQ),
.O5(CLBLL_R_X77Y130_SLICE_X118Y130_CO5),
.O6(CLBLL_R_X77Y130_SLICE_X118Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3030303064c4ff00)
  ) CLBLL_R_X77Y130_SLICE_X118Y130_BLUT (
.I0(CLBLL_R_X77Y130_SLICE_X118Y130_DO6),
.I1(CLBLL_R_X77Y130_SLICE_X118Y130_BQ),
.I2(CLBLL_R_X77Y130_SLICE_X118Y130_AQ),
.I3(CLBLL_R_X77Y130_SLICE_X118Y130_CQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLL_R_X77Y130_SLICE_X118Y130_BO5),
.O6(CLBLL_R_X77Y130_SLICE_X118Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa00cccc03030303)
  ) CLBLL_R_X77Y130_SLICE_X118Y130_ALUT (
.I0(CLBLL_R_X77Y130_SLICE_X118Y130_DO6),
.I1(CLBLM_L_X78Y131_SLICE_X120Y131_AQ),
.I2(CLBLL_R_X77Y130_SLICE_X118Y130_AQ),
.I3(CLBLL_R_X77Y131_SLICE_X118Y131_AO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLL_R_X77Y130_SLICE_X118Y130_AO5),
.O6(CLBLL_R_X77Y130_SLICE_X118Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y130_SLICE_X119Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X80Y132_SLICE_X124Y132_AQ),
.Q(CLBLL_R_X77Y130_SLICE_X119Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y130_SLICE_X119Y130_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y130_SLICE_X119Y130_BO6),
.Q(CLBLL_R_X77Y130_SLICE_X119Y130_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0055005500550055)
  ) CLBLL_R_X77Y130_SLICE_X119Y130_DLUT (
.I0(CLBLL_R_X77Y128_SLICE_X118Y128_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_R_X77Y130_SLICE_X119Y130_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y130_SLICE_X119Y130_DO5),
.O6(CLBLL_R_X77Y130_SLICE_X119Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000a8a8a8aa)
  ) CLBLL_R_X77Y130_SLICE_X119Y130_CLUT (
.I0(CLBLL_R_X77Y128_SLICE_X119Y128_BQ),
.I1(CLBLL_R_X77Y130_SLICE_X118Y130_AQ),
.I2(CLBLM_L_X78Y131_SLICE_X120Y131_AQ),
.I3(CLBLL_R_X77Y130_SLICE_X119Y130_AO5),
.I4(CLBLL_R_X77Y130_SLICE_X119Y130_DO6),
.I5(CLBLM_L_X78Y129_SLICE_X120Y129_BO6),
.O5(CLBLL_R_X77Y130_SLICE_X119Y130_CO5),
.O6(CLBLL_R_X77Y130_SLICE_X119Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcf2fcf8fc080c080)
  ) CLBLL_R_X77Y130_SLICE_X119Y130_BLUT (
.I0(CLBLM_L_X78Y130_SLICE_X120Y130_DO6),
.I1(CLBLL_R_X77Y130_SLICE_X119Y130_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLL_R_X77Y130_SLICE_X119Y130_DO6),
.I4(CLBLM_L_X78Y130_SLICE_X120Y130_AQ),
.I5(CLBLM_L_X78Y130_SLICE_X120Y130_BQ),
.O5(CLBLL_R_X77Y130_SLICE_X119Y130_BO5),
.O6(CLBLL_R_X77Y130_SLICE_X119Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0ff0f07ffff7ff)
  ) CLBLL_R_X77Y130_SLICE_X119Y130_ALUT (
.I0(CLBLL_R_X77Y131_SLICE_X119Y131_BQ),
.I1(CLBLL_R_X77Y130_SLICE_X119Y130_BQ),
.I2(CLBLL_R_X77Y128_SLICE_X118Y128_BQ),
.I3(CLBLM_L_X78Y130_SLICE_X120Y130_AQ),
.I4(CLBLL_R_X77Y128_SLICE_X118Y128_AQ),
.I5(1'b1),
.O5(CLBLL_R_X77Y130_SLICE_X119Y130_AO5),
.O6(CLBLL_R_X77Y130_SLICE_X119Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y131_SLICE_X118Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y131_SLICE_X118Y131_DO5),
.O6(CLBLL_R_X77Y131_SLICE_X118Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y131_SLICE_X118Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y131_SLICE_X118Y131_CO5),
.O6(CLBLL_R_X77Y131_SLICE_X118Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y131_SLICE_X118Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y131_SLICE_X118Y131_BO5),
.O6(CLBLL_R_X77Y131_SLICE_X118Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3d053d05ffffffc7)
  ) CLBLL_R_X77Y131_SLICE_X118Y131_ALUT (
.I0(CLBLL_R_X77Y130_SLICE_X119Y130_AQ),
.I1(CLBLL_R_X77Y128_SLICE_X118Y128_BQ),
.I2(CLBLL_R_X77Y128_SLICE_X118Y128_AQ),
.I3(CLBLM_L_X78Y131_SLICE_X120Y131_AQ),
.I4(CLBLL_R_X77Y130_SLICE_X118Y130_BO6),
.I5(CLBLL_R_X77Y131_SLICE_X119Y131_DO6),
.O5(CLBLL_R_X77Y131_SLICE_X118Y131_AO5),
.O6(CLBLL_R_X77Y131_SLICE_X118Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y131_SLICE_X119Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y131_SLICE_X119Y131_AO6),
.Q(CLBLL_R_X77Y131_SLICE_X119Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X77Y131_SLICE_X119Y131_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y131_SLICE_X119Y131_BO6),
.Q(CLBLL_R_X77Y131_SLICE_X119Y131_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888888888888888)
  ) CLBLL_R_X77Y131_SLICE_X119Y131_DLUT (
.I0(CLBLM_L_X78Y130_SLICE_X120Y130_BQ),
.I1(CLBLL_R_X77Y131_SLICE_X119Y131_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y131_SLICE_X119Y131_DO5),
.O6(CLBLL_R_X77Y131_SLICE_X119Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1f11ff11ff11ff11)
  ) CLBLL_R_X77Y131_SLICE_X119Y131_CLUT (
.I0(CLBLL_R_X77Y128_SLICE_X118Y128_AQ),
.I1(CLBLL_R_X77Y130_SLICE_X119Y130_AQ),
.I2(CLBLM_L_X78Y130_SLICE_X120Y130_AQ),
.I3(CLBLM_L_X78Y130_SLICE_X120Y130_DO6),
.I4(CLBLL_R_X77Y130_SLICE_X119Y130_BQ),
.I5(CLBLM_L_X78Y130_SLICE_X120Y130_BQ),
.O5(CLBLL_R_X77Y131_SLICE_X119Y131_CO5),
.O6(CLBLL_R_X77Y131_SLICE_X119Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccff002288ff00)
  ) CLBLL_R_X77Y131_SLICE_X119Y131_BLUT (
.I0(CLBLM_L_X78Y130_SLICE_X120Y130_DO6),
.I1(CLBLL_R_X77Y131_SLICE_X119Y131_BQ),
.I2(1'b1),
.I3(CLBLL_R_X77Y131_SLICE_X119Y131_AQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X77Y131_SLICE_X119Y131_CO6),
.O5(CLBLL_R_X77Y131_SLICE_X119Y131_BO5),
.O6(CLBLL_R_X77Y131_SLICE_X119Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3c0f3c03b083b08)
  ) CLBLL_R_X77Y131_SLICE_X119Y131_ALUT (
.I0(CLBLM_L_X78Y130_SLICE_X120Y130_DO6),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLL_R_X77Y131_SLICE_X119Y131_AQ),
.I3(CLBLL_R_X77Y130_SLICE_X119Y130_BQ),
.I4(1'b1),
.I5(CLBLL_R_X77Y131_SLICE_X119Y131_CO6),
.O5(CLBLL_R_X77Y131_SLICE_X119Y131_AO5),
.O6(CLBLL_R_X77Y131_SLICE_X119Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y96_SLICE_X122Y96_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y96_SLICE_X122Y96_DO5),
.O6(CLBLL_R_X79Y96_SLICE_X122Y96_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y96_SLICE_X122Y96_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y96_SLICE_X122Y96_CO5),
.O6(CLBLL_R_X79Y96_SLICE_X122Y96_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y96_SLICE_X122Y96_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y96_SLICE_X122Y96_BO5),
.O6(CLBLL_R_X79Y96_SLICE_X122Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fff0fff0fff0f)
  ) CLBLL_R_X79Y96_SLICE_X122Y96_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X103Y69_SLICE_X162Y69_A5Q),
.I3(CLBLM_L_X82Y98_SLICE_X128Y98_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y96_SLICE_X122Y96_AO5),
.O6(CLBLL_R_X79Y96_SLICE_X122Y96_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y96_SLICE_X123Y96_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y96_SLICE_X123Y96_DO5),
.O6(CLBLL_R_X79Y96_SLICE_X123Y96_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y96_SLICE_X123Y96_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y96_SLICE_X123Y96_CO5),
.O6(CLBLL_R_X79Y96_SLICE_X123Y96_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y96_SLICE_X123Y96_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y96_SLICE_X123Y96_BO5),
.O6(CLBLL_R_X79Y96_SLICE_X123Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y96_SLICE_X123Y96_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y96_SLICE_X123Y96_AO5),
.O6(CLBLL_R_X79Y96_SLICE_X123Y96_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y99_SLICE_X122Y99_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y99_SLICE_X122Y99_DO5),
.O6(CLBLL_R_X79Y99_SLICE_X122Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y99_SLICE_X122Y99_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y99_SLICE_X122Y99_CO5),
.O6(CLBLL_R_X79Y99_SLICE_X122Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y99_SLICE_X122Y99_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y99_SLICE_X122Y99_BO5),
.O6(CLBLL_R_X79Y99_SLICE_X122Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f000f000f000f0)
  ) CLBLL_R_X79Y99_SLICE_X122Y99_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X103Y69_SLICE_X162Y69_A5Q),
.I3(CLBLM_L_X82Y98_SLICE_X128Y98_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y99_SLICE_X122Y99_AO5),
.O6(CLBLL_R_X79Y99_SLICE_X122Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y99_SLICE_X123Y99_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y99_SLICE_X123Y99_DO5),
.O6(CLBLL_R_X79Y99_SLICE_X123Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y99_SLICE_X123Y99_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y99_SLICE_X123Y99_CO5),
.O6(CLBLL_R_X79Y99_SLICE_X123Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y99_SLICE_X123Y99_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y99_SLICE_X123Y99_BO5),
.O6(CLBLL_R_X79Y99_SLICE_X123Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y99_SLICE_X123Y99_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y99_SLICE_X123Y99_AO5),
.O6(CLBLL_R_X79Y99_SLICE_X123Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X79Y104_SLICE_X122Y104_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y103_SLICE_X115Y103_AQ),
.Q(CLBLL_R_X79Y104_SLICE_X122Y104_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X79Y104_SLICE_X122Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X79Y104_SLICE_X122Y104_AO6),
.Q(CLBLL_R_X79Y104_SLICE_X122Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X79Y104_SLICE_X122Y104_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X79Y104_SLICE_X122Y104_BO6),
.Q(CLBLL_R_X79Y104_SLICE_X122Y104_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y104_SLICE_X122Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y104_SLICE_X122Y104_DO5),
.O6(CLBLL_R_X79Y104_SLICE_X122Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y104_SLICE_X122Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y104_SLICE_X122Y104_CO5),
.O6(CLBLL_R_X79Y104_SLICE_X122Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5faf50a03fcf30c0)
  ) CLBLL_R_X79Y104_SLICE_X122Y104_BLUT (
.I0(CLBLM_L_X72Y118_SLICE_X108Y118_A5Q),
.I1(CLBLL_R_X75Y124_SLICE_X115Y124_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_R_X103Y76_SLICE_X162Y76_AO6),
.I4(CLBLM_R_X103Y76_SLICE_X162Y76_BQ),
.I5(CLBLL_R_X77Y104_SLICE_X118Y104_CQ),
.O5(CLBLL_R_X79Y104_SLICE_X122Y104_BO5),
.O6(CLBLL_R_X79Y104_SLICE_X122Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f50500fff00f0)
  ) CLBLL_R_X79Y104_SLICE_X122Y104_ALUT (
.I0(CLBLM_L_X72Y118_SLICE_X108Y118_A5Q),
.I1(1'b1),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLL_R_X75Y124_SLICE_X115Y124_BQ),
.I4(CLBLM_R_X103Y69_SLICE_X162Y69_A5Q),
.I5(CLBLL_R_X77Y104_SLICE_X118Y104_CQ),
.O5(CLBLL_R_X79Y104_SLICE_X122Y104_AO5),
.O6(CLBLL_R_X79Y104_SLICE_X122Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y104_SLICE_X123Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y104_SLICE_X123Y104_DO5),
.O6(CLBLL_R_X79Y104_SLICE_X123Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y104_SLICE_X123Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y104_SLICE_X123Y104_CO5),
.O6(CLBLL_R_X79Y104_SLICE_X123Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y104_SLICE_X123Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y104_SLICE_X123Y104_BO5),
.O6(CLBLL_R_X79Y104_SLICE_X123Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y104_SLICE_X123Y104_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y104_SLICE_X123Y104_AO5),
.O6(CLBLL_R_X79Y104_SLICE_X123Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X79Y127_SLICE_X122Y127_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X83Y130_SLICE_X130Y130_DQ),
.Q(CLBLL_R_X79Y127_SLICE_X122Y127_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X79Y127_SLICE_X122Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X79Y127_SLICE_X122Y127_AO6),
.Q(CLBLL_R_X79Y127_SLICE_X122Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X79Y127_SLICE_X122Y127_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X79Y127_SLICE_X122Y127_BO6),
.Q(CLBLL_R_X79Y127_SLICE_X122Y127_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X79Y127_SLICE_X122Y127_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X79Y127_SLICE_X122Y127_CO6),
.Q(CLBLL_R_X79Y127_SLICE_X122Y127_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699996666999966)
  ) CLBLL_R_X79Y127_SLICE_X122Y127_DLUT (
.I0(CLBLL_R_X79Y128_SLICE_X122Y128_AQ),
.I1(CLBLL_R_X79Y127_SLICE_X122Y127_CQ),
.I2(1'b1),
.I3(CLBLL_R_X79Y128_SLICE_X122Y128_CQ),
.I4(CLBLL_R_X79Y128_SLICE_X122Y128_DQ),
.I5(1'b1),
.O5(CLBLL_R_X79Y127_SLICE_X122Y127_DO5),
.O6(CLBLL_R_X79Y127_SLICE_X122Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccff00f0f0f0f0)
  ) CLBLL_R_X79Y127_SLICE_X122Y127_CLUT (
.I0(1'b1),
.I1(CLBLL_R_X79Y127_SLICE_X122Y127_CQ),
.I2(CLBLL_R_X79Y128_SLICE_X122Y128_BQ),
.I3(CLBLL_R_X83Y130_SLICE_X130Y130_CQ),
.I4(CLBLL_R_X77Y125_SLICE_X118Y125_BO5),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLL_R_X79Y127_SLICE_X122Y127_CO5),
.O6(CLBLL_R_X79Y127_SLICE_X122Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8ff00d8d8ff00)
  ) CLBLL_R_X79Y127_SLICE_X122Y127_BLUT (
.I0(CLBLL_R_X77Y125_SLICE_X118Y125_BO5),
.I1(CLBLL_R_X79Y127_SLICE_X122Y127_BQ),
.I2(CLBLL_R_X83Y130_SLICE_X130Y130_DQ),
.I3(CLBLL_R_X79Y127_SLICE_X122Y127_CQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLL_R_X79Y127_SLICE_X122Y127_BO5),
.O6(CLBLL_R_X79Y127_SLICE_X122Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5ffa0fff500a000)
  ) CLBLL_R_X79Y127_SLICE_X122Y127_ALUT (
.I0(CLBLL_R_X77Y125_SLICE_X118Y125_BO5),
.I1(1'b1),
.I2(CLBLL_R_X79Y127_SLICE_X122Y127_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLL_R_X77Y125_SLICE_X118Y125_AQ),
.I5(CLBLL_R_X79Y127_SLICE_X122Y127_A5Q),
.O5(CLBLL_R_X79Y127_SLICE_X122Y127_AO5),
.O6(CLBLL_R_X79Y127_SLICE_X122Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y127_SLICE_X123Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y127_SLICE_X123Y127_DO5),
.O6(CLBLL_R_X79Y127_SLICE_X123Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y127_SLICE_X123Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y127_SLICE_X123Y127_CO5),
.O6(CLBLL_R_X79Y127_SLICE_X123Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y127_SLICE_X123Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y127_SLICE_X123Y127_BO5),
.O6(CLBLL_R_X79Y127_SLICE_X123Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y127_SLICE_X123Y127_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y127_SLICE_X123Y127_AO5),
.O6(CLBLL_R_X79Y127_SLICE_X123Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X79Y128_SLICE_X122Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X79Y128_SLICE_X122Y128_AO6),
.Q(CLBLL_R_X79Y128_SLICE_X122Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X79Y128_SLICE_X122Y128_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X79Y128_SLICE_X122Y128_BO6),
.Q(CLBLL_R_X79Y128_SLICE_X122Y128_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X79Y128_SLICE_X122Y128_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X79Y128_SLICE_X122Y128_CO6),
.Q(CLBLL_R_X79Y128_SLICE_X122Y128_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X79Y128_SLICE_X122Y128_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X79Y128_SLICE_X122Y128_DO6),
.Q(CLBLL_R_X79Y128_SLICE_X122Y128_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aaaacccccccc)
  ) CLBLL_R_X79Y128_SLICE_X122Y128_DLUT (
.I0(CLBLL_R_X83Y130_SLICE_X130Y130_AQ),
.I1(CLBLL_R_X79Y128_SLICE_X122Y128_AQ),
.I2(CLBLL_R_X79Y128_SLICE_X122Y128_DQ),
.I3(1'b1),
.I4(CLBLL_R_X77Y125_SLICE_X118Y125_BO5),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLL_R_X79Y128_SLICE_X122Y128_DO5),
.O6(CLBLL_R_X79Y128_SLICE_X122Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cfc0aaaaaaaa)
  ) CLBLL_R_X79Y128_SLICE_X122Y128_CLUT (
.I0(CLBLL_R_X79Y127_SLICE_X122Y127_AQ),
.I1(CLBLL_R_X79Y128_SLICE_X122Y128_CQ),
.I2(CLBLL_R_X77Y125_SLICE_X118Y125_BO5),
.I3(CLBLM_L_X82Y130_SLICE_X128Y130_AQ),
.I4(1'b1),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLL_R_X79Y128_SLICE_X122Y128_CO5),
.O6(CLBLL_R_X79Y128_SLICE_X122Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8888f0f0f0f0)
  ) CLBLL_R_X79Y128_SLICE_X122Y128_BLUT (
.I0(CLBLL_R_X77Y125_SLICE_X118Y125_BO5),
.I1(CLBLL_R_X79Y128_SLICE_X122Y128_BQ),
.I2(CLBLL_R_X79Y128_SLICE_X122Y128_DQ),
.I3(1'b1),
.I4(CLBLL_R_X83Y130_SLICE_X130Y130_BQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLL_R_X79Y128_SLICE_X122Y128_BO5),
.O6(CLBLL_R_X79Y128_SLICE_X122Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he4ffe400e4ffe400)
  ) CLBLL_R_X79Y128_SLICE_X122Y128_ALUT (
.I0(CLBLL_R_X77Y125_SLICE_X118Y125_BO5),
.I1(CLBLL_R_X83Y132_SLICE_X130Y132_AQ),
.I2(CLBLL_R_X79Y128_SLICE_X122Y128_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLL_R_X79Y128_SLICE_X122Y128_CQ),
.I5(1'b1),
.O5(CLBLL_R_X79Y128_SLICE_X122Y128_AO5),
.O6(CLBLL_R_X79Y128_SLICE_X122Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y128_SLICE_X123Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y128_SLICE_X123Y128_DO5),
.O6(CLBLL_R_X79Y128_SLICE_X123Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y128_SLICE_X123Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y128_SLICE_X123Y128_CO5),
.O6(CLBLL_R_X79Y128_SLICE_X123Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y128_SLICE_X123Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y128_SLICE_X123Y128_BO5),
.O6(CLBLL_R_X79Y128_SLICE_X123Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y128_SLICE_X123Y128_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y128_SLICE_X123Y128_AO5),
.O6(CLBLL_R_X79Y128_SLICE_X123Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X79Y135_SLICE_X122Y135_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y133_SLICE_X114Y133_BQ),
.Q(CLBLL_R_X79Y135_SLICE_X122Y135_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y135_SLICE_X122Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y135_SLICE_X122Y135_DO5),
.O6(CLBLL_R_X79Y135_SLICE_X122Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y135_SLICE_X122Y135_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y135_SLICE_X122Y135_CO5),
.O6(CLBLL_R_X79Y135_SLICE_X122Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y135_SLICE_X122Y135_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y135_SLICE_X122Y135_BO5),
.O6(CLBLL_R_X79Y135_SLICE_X122Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y135_SLICE_X122Y135_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y135_SLICE_X122Y135_AO5),
.O6(CLBLL_R_X79Y135_SLICE_X122Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y135_SLICE_X123Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y135_SLICE_X123Y135_DO5),
.O6(CLBLL_R_X79Y135_SLICE_X123Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y135_SLICE_X123Y135_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y135_SLICE_X123Y135_CO5),
.O6(CLBLL_R_X79Y135_SLICE_X123Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y135_SLICE_X123Y135_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y135_SLICE_X123Y135_BO5),
.O6(CLBLL_R_X79Y135_SLICE_X123Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y135_SLICE_X123Y135_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y135_SLICE_X123Y135_AO5),
.O6(CLBLL_R_X79Y135_SLICE_X123Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X83Y94_SLICE_X130Y94_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X83Y94_SLICE_X130Y94_AO5),
.Q(CLBLL_R_X83Y94_SLICE_X130Y94_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X83Y94_SLICE_X130Y94_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X83Y94_SLICE_X130Y94_AO6),
.Q(CLBLL_R_X83Y94_SLICE_X130Y94_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X83Y94_SLICE_X130Y94_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X83Y94_SLICE_X130Y94_A5Q),
.Q(CLBLL_R_X83Y94_SLICE_X130Y94_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X83Y94_SLICE_X130Y94_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X83Y94_SLICE_X130Y94_DO5),
.O6(CLBLL_R_X83Y94_SLICE_X130Y94_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X83Y94_SLICE_X130Y94_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X83Y94_SLICE_X130Y94_CO5),
.O6(CLBLL_R_X83Y94_SLICE_X130Y94_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X83Y94_SLICE_X130Y94_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X83Y94_SLICE_X130Y94_BO5),
.O6(CLBLL_R_X83Y94_SLICE_X130Y94_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6666cccc77227722)
  ) CLBLL_R_X83Y94_SLICE_X130Y94_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X83Y94_SLICE_X130Y94_BQ),
.I2(1'b1),
.I3(CLBLM_L_X82Y98_SLICE_X128Y98_A5Q),
.I4(CLBLL_R_X83Y94_SLICE_X130Y94_A5Q),
.I5(1'b1),
.O5(CLBLL_R_X83Y94_SLICE_X130Y94_AO5),
.O6(CLBLL_R_X83Y94_SLICE_X130Y94_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X83Y94_SLICE_X131Y94_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X83Y94_SLICE_X131Y94_DO5),
.O6(CLBLL_R_X83Y94_SLICE_X131Y94_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X83Y94_SLICE_X131Y94_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X83Y94_SLICE_X131Y94_CO5),
.O6(CLBLL_R_X83Y94_SLICE_X131Y94_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X83Y94_SLICE_X131Y94_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X83Y94_SLICE_X131Y94_BO5),
.O6(CLBLL_R_X83Y94_SLICE_X131Y94_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X83Y94_SLICE_X131Y94_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X83Y94_SLICE_X131Y94_AO5),
.O6(CLBLL_R_X83Y94_SLICE_X131Y94_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X83Y130_SLICE_X130Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X83Y132_SLICE_X130Y132_AQ),
.Q(CLBLL_R_X83Y130_SLICE_X130Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X83Y130_SLICE_X130Y130_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X83Y130_SLICE_X130Y130_AQ),
.Q(CLBLL_R_X83Y130_SLICE_X130Y130_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X83Y130_SLICE_X130Y130_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X83Y130_SLICE_X130Y130_BQ),
.Q(CLBLL_R_X83Y130_SLICE_X130Y130_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X83Y130_SLICE_X130Y130_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X83Y130_SLICE_X130Y130_CQ),
.Q(CLBLL_R_X83Y130_SLICE_X130Y130_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X83Y130_SLICE_X130Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X83Y130_SLICE_X130Y130_DO5),
.O6(CLBLL_R_X83Y130_SLICE_X130Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X83Y130_SLICE_X130Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X83Y130_SLICE_X130Y130_CO5),
.O6(CLBLL_R_X83Y130_SLICE_X130Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X83Y130_SLICE_X130Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X83Y130_SLICE_X130Y130_BO5),
.O6(CLBLL_R_X83Y130_SLICE_X130Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X83Y130_SLICE_X130Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X83Y130_SLICE_X130Y130_AO5),
.O6(CLBLL_R_X83Y130_SLICE_X130Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X83Y130_SLICE_X131Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X83Y130_SLICE_X131Y130_DO5),
.O6(CLBLL_R_X83Y130_SLICE_X131Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X83Y130_SLICE_X131Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X83Y130_SLICE_X131Y130_CO5),
.O6(CLBLL_R_X83Y130_SLICE_X131Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X83Y130_SLICE_X131Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X83Y130_SLICE_X131Y130_BO5),
.O6(CLBLL_R_X83Y130_SLICE_X131Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X83Y130_SLICE_X131Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X83Y130_SLICE_X131Y130_AO5),
.O6(CLBLL_R_X83Y130_SLICE_X131Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X83Y132_SLICE_X130Y132_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X82Y130_SLICE_X128Y130_AQ),
.Q(CLBLL_R_X83Y132_SLICE_X130Y132_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X83Y132_SLICE_X130Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X83Y132_SLICE_X130Y132_DO5),
.O6(CLBLL_R_X83Y132_SLICE_X130Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X83Y132_SLICE_X130Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X83Y132_SLICE_X130Y132_CO5),
.O6(CLBLL_R_X83Y132_SLICE_X130Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X83Y132_SLICE_X130Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X83Y132_SLICE_X130Y132_BO5),
.O6(CLBLL_R_X83Y132_SLICE_X130Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X83Y132_SLICE_X130Y132_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X83Y132_SLICE_X130Y132_AO5),
.O6(CLBLL_R_X83Y132_SLICE_X130Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X83Y132_SLICE_X131Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X83Y132_SLICE_X131Y132_DO5),
.O6(CLBLL_R_X83Y132_SLICE_X131Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X83Y132_SLICE_X131Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X83Y132_SLICE_X131Y132_CO5),
.O6(CLBLL_R_X83Y132_SLICE_X131Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X83Y132_SLICE_X131Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X83Y132_SLICE_X131Y132_BO5),
.O6(CLBLL_R_X83Y132_SLICE_X131Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X83Y132_SLICE_X131Y132_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X83Y132_SLICE_X131Y132_AO5),
.O6(CLBLL_R_X83Y132_SLICE_X131Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y92_SLICE_X90Y92_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y134_SLICE_X106Y134_AQ),
.Q(CLBLM_L_X60Y92_SLICE_X90Y92_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y92_SLICE_X90Y92_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.Q(CLBLM_L_X60Y92_SLICE_X90Y92_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y92_SLICE_X90Y92_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y92_SLICE_X90Y92_DO5),
.O6(CLBLM_L_X60Y92_SLICE_X90Y92_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y92_SLICE_X90Y92_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y92_SLICE_X90Y92_CO5),
.O6(CLBLM_L_X60Y92_SLICE_X90Y92_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y92_SLICE_X90Y92_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y92_SLICE_X90Y92_BO5),
.O6(CLBLM_L_X60Y92_SLICE_X90Y92_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y92_SLICE_X90Y92_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y92_SLICE_X90Y92_AO5),
.O6(CLBLM_L_X60Y92_SLICE_X90Y92_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y92_SLICE_X91Y92_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y92_SLICE_X91Y92_DO5),
.O6(CLBLM_L_X60Y92_SLICE_X91Y92_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y92_SLICE_X91Y92_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y92_SLICE_X91Y92_CO5),
.O6(CLBLM_L_X60Y92_SLICE_X91Y92_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y92_SLICE_X91Y92_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y92_SLICE_X91Y92_BO5),
.O6(CLBLM_L_X60Y92_SLICE_X91Y92_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y92_SLICE_X91Y92_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y92_SLICE_X91Y92_AO5),
.O6(CLBLM_L_X60Y92_SLICE_X91Y92_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y94_SLICE_X90Y94_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X60Y92_SLICE_X90Y92_AQ),
.Q(CLBLM_L_X60Y94_SLICE_X90Y94_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y94_SLICE_X90Y94_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y95_SLICE_X92Y95_BQ),
.Q(CLBLM_L_X60Y94_SLICE_X90Y94_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y94_SLICE_X90Y94_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X60Y94_SLICE_X90Y94_BQ),
.Q(CLBLM_L_X60Y94_SLICE_X90Y94_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y94_SLICE_X90Y94_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y94_SLICE_X90Y94_DO5),
.O6(CLBLM_L_X60Y94_SLICE_X90Y94_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y94_SLICE_X90Y94_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y94_SLICE_X90Y94_CO5),
.O6(CLBLM_L_X60Y94_SLICE_X90Y94_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y94_SLICE_X90Y94_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y94_SLICE_X90Y94_BO5),
.O6(CLBLM_L_X60Y94_SLICE_X90Y94_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y94_SLICE_X90Y94_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y94_SLICE_X90Y94_AO5),
.O6(CLBLM_L_X60Y94_SLICE_X90Y94_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y94_SLICE_X91Y94_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y94_SLICE_X91Y94_DO5),
.O6(CLBLM_L_X60Y94_SLICE_X91Y94_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y94_SLICE_X91Y94_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y94_SLICE_X91Y94_CO5),
.O6(CLBLM_L_X60Y94_SLICE_X91Y94_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y94_SLICE_X91Y94_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y94_SLICE_X91Y94_BO5),
.O6(CLBLM_L_X60Y94_SLICE_X91Y94_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y94_SLICE_X91Y94_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y94_SLICE_X91Y94_AO5),
.O6(CLBLM_L_X60Y94_SLICE_X91Y94_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y97_SLICE_X90Y97_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y107_SLICE_X93Y107_A5Q),
.Q(CLBLM_L_X60Y97_SLICE_X90Y97_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y97_SLICE_X90Y97_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X60Y99_SLICE_X90Y99_AQ),
.Q(CLBLM_L_X60Y97_SLICE_X90Y97_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y97_SLICE_X90Y97_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y98_SLICE_X94Y98_BQ),
.Q(CLBLM_L_X60Y97_SLICE_X90Y97_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y97_SLICE_X90Y97_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y97_SLICE_X103Y97_AQ),
.Q(CLBLM_L_X60Y97_SLICE_X90Y97_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y97_SLICE_X90Y97_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y97_SLICE_X90Y97_DO5),
.O6(CLBLM_L_X60Y97_SLICE_X90Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y97_SLICE_X90Y97_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y97_SLICE_X90Y97_CO5),
.O6(CLBLM_L_X60Y97_SLICE_X90Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y97_SLICE_X90Y97_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y97_SLICE_X90Y97_BO5),
.O6(CLBLM_L_X60Y97_SLICE_X90Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y97_SLICE_X90Y97_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y97_SLICE_X90Y97_AO5),
.O6(CLBLM_L_X60Y97_SLICE_X90Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y97_SLICE_X91Y97_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y110_SLICE_X99Y110_B5Q),
.Q(CLBLM_L_X60Y97_SLICE_X91Y97_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y97_SLICE_X91Y97_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y97_SLICE_X91Y97_DO5),
.O6(CLBLM_L_X60Y97_SLICE_X91Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y97_SLICE_X91Y97_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y97_SLICE_X91Y97_CO5),
.O6(CLBLM_L_X60Y97_SLICE_X91Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y97_SLICE_X91Y97_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y97_SLICE_X91Y97_BO5),
.O6(CLBLM_L_X60Y97_SLICE_X91Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y97_SLICE_X91Y97_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y97_SLICE_X91Y97_AO5),
.O6(CLBLM_L_X60Y97_SLICE_X91Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y99_SLICE_X90Y99_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y100_SLICE_X105Y100_CQ),
.Q(CLBLM_L_X60Y99_SLICE_X90Y99_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y99_SLICE_X90Y99_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X60Y99_SLICE_X90Y99_DQ),
.Q(CLBLM_L_X60Y99_SLICE_X90Y99_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y99_SLICE_X90Y99_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X60Y99_SLICE_X90Y99_BQ),
.Q(CLBLM_L_X60Y99_SLICE_X90Y99_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y99_SLICE_X90Y99_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y101_SLICE_X92Y101_AQ),
.Q(CLBLM_L_X60Y99_SLICE_X90Y99_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y99_SLICE_X90Y99_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y99_SLICE_X90Y99_DO5),
.O6(CLBLM_L_X60Y99_SLICE_X90Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y99_SLICE_X90Y99_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y99_SLICE_X90Y99_CO5),
.O6(CLBLM_L_X60Y99_SLICE_X90Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y99_SLICE_X90Y99_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y99_SLICE_X90Y99_BO5),
.O6(CLBLM_L_X60Y99_SLICE_X90Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y99_SLICE_X90Y99_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y99_SLICE_X90Y99_AO5),
.O6(CLBLM_L_X60Y99_SLICE_X90Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y99_SLICE_X91Y99_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y99_SLICE_X91Y99_DO5),
.O6(CLBLM_L_X60Y99_SLICE_X91Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y99_SLICE_X91Y99_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y99_SLICE_X91Y99_CO5),
.O6(CLBLM_L_X60Y99_SLICE_X91Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y99_SLICE_X91Y99_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y99_SLICE_X91Y99_BO5),
.O6(CLBLM_L_X60Y99_SLICE_X91Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y99_SLICE_X91Y99_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y99_SLICE_X91Y99_AO5),
.O6(CLBLM_L_X60Y99_SLICE_X91Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y101_SLICE_X90Y101_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y95_SLICE_X92Y95_AQ),
.Q(CLBLM_L_X60Y101_SLICE_X90Y101_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y101_SLICE_X90Y101_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.Q(CLBLM_L_X60Y101_SLICE_X90Y101_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y101_SLICE_X90Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y101_SLICE_X90Y101_DO5),
.O6(CLBLM_L_X60Y101_SLICE_X90Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y101_SLICE_X90Y101_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y101_SLICE_X90Y101_CO5),
.O6(CLBLM_L_X60Y101_SLICE_X90Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y101_SLICE_X90Y101_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y101_SLICE_X90Y101_BO5),
.O6(CLBLM_L_X60Y101_SLICE_X90Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y101_SLICE_X90Y101_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y101_SLICE_X90Y101_AO5),
.O6(CLBLM_L_X60Y101_SLICE_X90Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y101_SLICE_X91Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y101_SLICE_X91Y101_DO5),
.O6(CLBLM_L_X60Y101_SLICE_X91Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y101_SLICE_X91Y101_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y101_SLICE_X91Y101_CO5),
.O6(CLBLM_L_X60Y101_SLICE_X91Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y101_SLICE_X91Y101_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y101_SLICE_X91Y101_BO5),
.O6(CLBLM_L_X60Y101_SLICE_X91Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y101_SLICE_X91Y101_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y101_SLICE_X91Y101_AO5),
.O6(CLBLM_L_X60Y101_SLICE_X91Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y104_SLICE_X90Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y127_SLICE_X115Y127_AQ),
.Q(CLBLM_L_X60Y104_SLICE_X90Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y104_SLICE_X90Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y104_SLICE_X90Y104_DO5),
.O6(CLBLM_L_X60Y104_SLICE_X90Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y104_SLICE_X90Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y104_SLICE_X90Y104_CO5),
.O6(CLBLM_L_X60Y104_SLICE_X90Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y104_SLICE_X90Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y104_SLICE_X90Y104_BO5),
.O6(CLBLM_L_X60Y104_SLICE_X90Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y104_SLICE_X90Y104_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y104_SLICE_X90Y104_AO5),
.O6(CLBLM_L_X60Y104_SLICE_X90Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y104_SLICE_X91Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y104_SLICE_X91Y104_DO5),
.O6(CLBLM_L_X60Y104_SLICE_X91Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y104_SLICE_X91Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y104_SLICE_X91Y104_CO5),
.O6(CLBLM_L_X60Y104_SLICE_X91Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y104_SLICE_X91Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y104_SLICE_X91Y104_BO5),
.O6(CLBLM_L_X60Y104_SLICE_X91Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y104_SLICE_X91Y104_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y104_SLICE_X91Y104_AO5),
.O6(CLBLM_L_X60Y104_SLICE_X91Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y90_SLICE_X92Y90_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y106_SLICE_X108Y106_A5Q),
.Q(CLBLM_L_X62Y90_SLICE_X92Y90_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y90_SLICE_X92Y90_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y90_SLICE_X92Y90_DO5),
.O6(CLBLM_L_X62Y90_SLICE_X92Y90_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y90_SLICE_X92Y90_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y90_SLICE_X92Y90_CO5),
.O6(CLBLM_L_X62Y90_SLICE_X92Y90_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y90_SLICE_X92Y90_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y90_SLICE_X92Y90_BO5),
.O6(CLBLM_L_X62Y90_SLICE_X92Y90_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y90_SLICE_X92Y90_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y90_SLICE_X92Y90_AO5),
.O6(CLBLM_L_X62Y90_SLICE_X92Y90_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y90_SLICE_X93Y90_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y90_SLICE_X93Y90_DO5),
.O6(CLBLM_L_X62Y90_SLICE_X93Y90_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y90_SLICE_X93Y90_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y90_SLICE_X93Y90_CO5),
.O6(CLBLM_L_X62Y90_SLICE_X93Y90_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y90_SLICE_X93Y90_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y90_SLICE_X93Y90_BO5),
.O6(CLBLM_L_X62Y90_SLICE_X93Y90_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y90_SLICE_X93Y90_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y90_SLICE_X93Y90_AO5),
.O6(CLBLM_L_X62Y90_SLICE_X93Y90_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y92_SLICE_X92Y92_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y90_SLICE_X92Y90_AQ),
.Q(CLBLM_L_X62Y92_SLICE_X92Y92_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y92_SLICE_X92Y92_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X60Y97_SLICE_X91Y97_AQ),
.Q(CLBLM_L_X62Y92_SLICE_X92Y92_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y92_SLICE_X92Y92_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y92_SLICE_X92Y92_DO5),
.O6(CLBLM_L_X62Y92_SLICE_X92Y92_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y92_SLICE_X92Y92_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y92_SLICE_X92Y92_CO5),
.O6(CLBLM_L_X62Y92_SLICE_X92Y92_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y92_SLICE_X92Y92_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y92_SLICE_X92Y92_BO5),
.O6(CLBLM_L_X62Y92_SLICE_X92Y92_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y92_SLICE_X92Y92_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y92_SLICE_X92Y92_AO5),
.O6(CLBLM_L_X62Y92_SLICE_X92Y92_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y92_SLICE_X93Y92_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y92_SLICE_X93Y92_DO5),
.O6(CLBLM_L_X62Y92_SLICE_X93Y92_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y92_SLICE_X93Y92_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y92_SLICE_X93Y92_CO5),
.O6(CLBLM_L_X62Y92_SLICE_X93Y92_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y92_SLICE_X93Y92_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y92_SLICE_X93Y92_BO5),
.O6(CLBLM_L_X62Y92_SLICE_X93Y92_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y92_SLICE_X93Y92_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y92_SLICE_X93Y92_AO5),
.O6(CLBLM_L_X62Y92_SLICE_X93Y92_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y95_SLICE_X92Y95_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y103_SLICE_X111Y103_A5Q),
.Q(CLBLM_L_X62Y95_SLICE_X92Y95_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y95_SLICE_X92Y95_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y95_SLICE_X102Y95_A5Q),
.Q(CLBLM_L_X62Y95_SLICE_X92Y95_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y95_SLICE_X92Y95_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X60Y97_SLICE_X90Y97_DQ),
.Q(CLBLM_L_X62Y95_SLICE_X92Y95_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y95_SLICE_X92Y95_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y95_SLICE_X92Y95_DO5),
.O6(CLBLM_L_X62Y95_SLICE_X92Y95_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y95_SLICE_X92Y95_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y95_SLICE_X92Y95_CO5),
.O6(CLBLM_L_X62Y95_SLICE_X92Y95_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y95_SLICE_X92Y95_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y95_SLICE_X92Y95_BO5),
.O6(CLBLM_L_X62Y95_SLICE_X92Y95_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y95_SLICE_X92Y95_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y95_SLICE_X92Y95_AO5),
.O6(CLBLM_L_X62Y95_SLICE_X92Y95_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y95_SLICE_X93Y95_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y95_SLICE_X93Y95_DO5),
.O6(CLBLM_L_X62Y95_SLICE_X93Y95_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y95_SLICE_X93Y95_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y95_SLICE_X93Y95_CO5),
.O6(CLBLM_L_X62Y95_SLICE_X93Y95_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y95_SLICE_X93Y95_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y95_SLICE_X93Y95_BO5),
.O6(CLBLM_L_X62Y95_SLICE_X93Y95_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y95_SLICE_X93Y95_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y95_SLICE_X93Y95_AO5),
.O6(CLBLM_L_X62Y95_SLICE_X93Y95_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y97_SLICE_X92Y97_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y97_SLICE_X92Y97_DO5),
.O6(CLBLM_L_X62Y97_SLICE_X92Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y97_SLICE_X92Y97_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y97_SLICE_X92Y97_CO5),
.O6(CLBLM_L_X62Y97_SLICE_X92Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y97_SLICE_X92Y97_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y97_SLICE_X92Y97_BO5),
.O6(CLBLM_L_X62Y97_SLICE_X92Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y97_SLICE_X92Y97_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y97_SLICE_X92Y97_AO5),
.O6(CLBLM_L_X62Y97_SLICE_X92Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y97_SLICE_X93Y97_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y97_SLICE_X93Y97_AO6),
.Q(CLBLM_L_X62Y97_SLICE_X93Y97_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y97_SLICE_X93Y97_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y97_SLICE_X93Y97_BO6),
.Q(CLBLM_L_X62Y97_SLICE_X93Y97_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y97_SLICE_X93Y97_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y97_SLICE_X93Y97_DO5),
.O6(CLBLM_L_X62Y97_SLICE_X93Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y97_SLICE_X93Y97_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y97_SLICE_X93Y97_CO5),
.O6(CLBLM_L_X62Y97_SLICE_X93Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0f0ccaaf0f0)
  ) CLBLM_L_X62Y97_SLICE_X93Y97_BLUT (
.I0(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I1(CLBLM_L_X62Y97_SLICE_X93Y97_BQ),
.I2(CLBLM_L_X62Y97_SLICE_X93Y97_AQ),
.I3(CLBLM_R_X63Y99_SLICE_X94Y99_CO5),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X64Y97_SLICE_X97Y97_BO6),
.O5(CLBLM_L_X62Y97_SLICE_X93Y97_BO5),
.O6(CLBLM_L_X62Y97_SLICE_X93Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000e2ffe200)
  ) CLBLM_L_X62Y97_SLICE_X93Y97_ALUT (
.I0(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I1(CLBLM_R_X63Y99_SLICE_X94Y99_CO6),
.I2(CLBLM_L_X62Y97_SLICE_X93Y97_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_R_X63Y96_SLICE_X94Y96_BQ),
.I5(CLBLM_L_X64Y97_SLICE_X97Y97_BO6),
.O5(CLBLM_L_X62Y97_SLICE_X93Y97_AO5),
.O6(CLBLM_L_X62Y97_SLICE_X93Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y98_SLICE_X92Y98_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y98_SLICE_X92Y98_DO5),
.O6(CLBLM_L_X62Y98_SLICE_X92Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y98_SLICE_X92Y98_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y98_SLICE_X92Y98_CO5),
.O6(CLBLM_L_X62Y98_SLICE_X92Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y98_SLICE_X92Y98_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y98_SLICE_X92Y98_BO5),
.O6(CLBLM_L_X62Y98_SLICE_X92Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y98_SLICE_X92Y98_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y98_SLICE_X92Y98_AO5),
.O6(CLBLM_L_X62Y98_SLICE_X92Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y98_SLICE_X93Y98_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y98_SLICE_X93Y98_AO6),
.Q(CLBLM_L_X62Y98_SLICE_X93Y98_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y98_SLICE_X93Y98_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y98_SLICE_X93Y98_BO6),
.Q(CLBLM_L_X62Y98_SLICE_X93Y98_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y98_SLICE_X93Y98_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y98_SLICE_X93Y98_CO6),
.Q(CLBLM_L_X62Y98_SLICE_X93Y98_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y98_SLICE_X93Y98_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y98_SLICE_X93Y98_DO5),
.O6(CLBLM_L_X62Y98_SLICE_X93Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaacfaaccaac0aa)
  ) CLBLM_L_X62Y98_SLICE_X93Y98_CLUT (
.I0(CLBLM_L_X62Y98_SLICE_X93Y98_BQ),
.I1(CLBLM_L_X62Y98_SLICE_X93Y98_CQ),
.I2(CLBLM_R_X63Y99_SLICE_X94Y99_CO5),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X64Y98_SLICE_X96Y98_AO5),
.I5(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.O5(CLBLM_L_X62Y98_SLICE_X93Y98_CO5),
.O6(CLBLM_L_X62Y98_SLICE_X93Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa5050fad850d8)
  ) CLBLM_L_X62Y98_SLICE_X93Y98_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I2(CLBLM_L_X62Y98_SLICE_X93Y98_AQ),
.I3(CLBLM_R_X63Y99_SLICE_X94Y99_CO6),
.I4(CLBLM_L_X62Y98_SLICE_X93Y98_BQ),
.I5(CLBLM_L_X64Y98_SLICE_X96Y98_AO5),
.O5(CLBLM_L_X62Y98_SLICE_X93Y98_BO5),
.O6(CLBLM_L_X62Y98_SLICE_X93Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f5a0cccccccc)
  ) CLBLM_L_X62Y98_SLICE_X93Y98_ALUT (
.I0(CLBLM_L_X64Y98_SLICE_X96Y98_AO5),
.I1(CLBLM_L_X64Y98_SLICE_X96Y98_BQ),
.I2(CLBLM_L_X62Y98_SLICE_X93Y98_AQ),
.I3(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I4(CLBLM_R_X63Y99_SLICE_X94Y99_BO5),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X62Y98_SLICE_X93Y98_AO5),
.O6(CLBLM_L_X62Y98_SLICE_X93Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y99_SLICE_X92Y99_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y99_SLICE_X92Y99_DO5),
.O6(CLBLM_L_X62Y99_SLICE_X92Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y99_SLICE_X92Y99_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y99_SLICE_X92Y99_CO5),
.O6(CLBLM_L_X62Y99_SLICE_X92Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y99_SLICE_X92Y99_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y99_SLICE_X92Y99_BO5),
.O6(CLBLM_L_X62Y99_SLICE_X92Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y99_SLICE_X92Y99_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y99_SLICE_X92Y99_AO5),
.O6(CLBLM_L_X62Y99_SLICE_X92Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y99_SLICE_X93Y99_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y99_SLICE_X93Y99_AO6),
.Q(CLBLM_L_X62Y99_SLICE_X93Y99_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y99_SLICE_X93Y99_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y99_SLICE_X93Y99_DO5),
.O6(CLBLM_L_X62Y99_SLICE_X93Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y99_SLICE_X93Y99_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y99_SLICE_X93Y99_CO5),
.O6(CLBLM_L_X62Y99_SLICE_X93Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h80c0a2f300000000)
  ) CLBLM_L_X62Y99_SLICE_X93Y99_BLUT (
.I0(CLBLM_L_X60Y92_SLICE_X90Y92_BQ),
.I1(CLBLM_L_X76Y111_SLICE_X116Y111_BQ),
.I2(CLBLM_L_X62Y99_SLICE_X93Y99_AQ),
.I3(CLBLM_R_X63Y98_SLICE_X94Y98_AQ),
.I4(CLBLM_R_X63Y98_SLICE_X94Y98_BQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X62Y99_SLICE_X93Y99_BO5),
.O6(CLBLM_L_X62Y99_SLICE_X93Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f00000055005500)
  ) CLBLM_L_X62Y99_SLICE_X93Y99_ALUT (
.I0(CLBLM_L_X60Y92_SLICE_X90Y92_BQ),
.I1(CLBLM_L_X76Y111_SLICE_X116Y111_BQ),
.I2(CLBLM_L_X62Y99_SLICE_X93Y99_AQ),
.I3(CLBLM_L_X62Y99_SLICE_X93Y99_BO6),
.I4(CLBLM_R_X63Y98_SLICE_X94Y98_BQ),
.I5(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.O5(CLBLM_L_X62Y99_SLICE_X93Y99_AO5),
.O6(CLBLM_L_X62Y99_SLICE_X93Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y100_SLICE_X92Y100_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y100_SLICE_X92Y100_AO6),
.Q(CLBLM_L_X62Y100_SLICE_X92Y100_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y100_SLICE_X92Y100_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y100_SLICE_X92Y100_DO5),
.O6(CLBLM_L_X62Y100_SLICE_X92Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y100_SLICE_X92Y100_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y100_SLICE_X92Y100_CO5),
.O6(CLBLM_L_X62Y100_SLICE_X92Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y100_SLICE_X92Y100_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y100_SLICE_X92Y100_BO5),
.O6(CLBLM_L_X62Y100_SLICE_X92Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4c4c00cc000000cc)
  ) CLBLM_L_X62Y100_SLICE_X92Y100_ALUT (
.I0(CLBLM_L_X62Y101_SLICE_X92Y101_AQ),
.I1(CLBLM_L_X62Y101_SLICE_X92Y101_BO6),
.I2(CLBLM_L_X62Y100_SLICE_X92Y100_AQ),
.I3(CLBLM_L_X60Y99_SLICE_X90Y99_CQ),
.I4(CLBLM_L_X60Y99_SLICE_X90Y99_BQ),
.I5(CLBLM_L_X60Y99_SLICE_X90Y99_DQ),
.O5(CLBLM_L_X62Y100_SLICE_X92Y100_AO5),
.O6(CLBLM_L_X62Y100_SLICE_X92Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y100_SLICE_X93Y100_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y100_SLICE_X93Y100_DO5),
.O6(CLBLM_L_X62Y100_SLICE_X93Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y100_SLICE_X93Y100_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y100_SLICE_X93Y100_CO5),
.O6(CLBLM_L_X62Y100_SLICE_X93Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y100_SLICE_X93Y100_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y100_SLICE_X93Y100_BO5),
.O6(CLBLM_L_X62Y100_SLICE_X93Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0000000000000)
  ) CLBLM_L_X62Y100_SLICE_X93Y100_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X60Y99_SLICE_X90Y99_DQ),
.I2(CLBLM_L_X60Y99_SLICE_X90Y99_BQ),
.I3(1'b1),
.I4(CLBLM_L_X62Y100_SLICE_X92Y100_AQ),
.I5(CLBLM_L_X62Y101_SLICE_X92Y101_AQ),
.O5(CLBLM_L_X62Y100_SLICE_X93Y100_AO5),
.O6(CLBLM_L_X62Y100_SLICE_X93Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y101_SLICE_X92Y101_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y100_SLICE_X92Y100_AQ),
.Q(CLBLM_L_X62Y101_SLICE_X92Y101_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y101_SLICE_X92Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y101_SLICE_X92Y101_DO5),
.O6(CLBLM_L_X62Y101_SLICE_X92Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y101_SLICE_X92Y101_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y101_SLICE_X92Y101_CO5),
.O6(CLBLM_L_X62Y101_SLICE_X92Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0400000cc440c04)
  ) CLBLM_L_X62Y101_SLICE_X92Y101_BLUT (
.I0(CLBLM_R_X63Y101_SLICE_X94Y101_AQ),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_L_X62Y101_SLICE_X92Y101_AQ),
.I3(CLBLM_L_X60Y99_SLICE_X90Y99_CQ),
.I4(CLBLM_L_X62Y100_SLICE_X92Y100_AQ),
.I5(CLBLM_L_X60Y99_SLICE_X90Y99_DQ),
.O5(CLBLM_L_X62Y101_SLICE_X92Y101_BO5),
.O6(CLBLM_L_X62Y101_SLICE_X92Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00a000a0cc000000)
  ) CLBLM_L_X62Y101_SLICE_X92Y101_ALUT (
.I0(CLBLM_L_X60Y99_SLICE_X90Y99_BQ),
.I1(CLBLM_L_X62Y102_SLICE_X92Y102_BQ),
.I2(CLBLM_L_X62Y102_SLICE_X92Y102_CQ),
.I3(CLBLM_L_X64Y101_SLICE_X96Y101_B5Q),
.I4(CLBLM_L_X60Y99_SLICE_X90Y99_DQ),
.I5(CLBLM_L_X64Y101_SLICE_X96Y101_BQ),
.O5(CLBLM_L_X62Y101_SLICE_X92Y101_AO5),
.O6(CLBLM_L_X62Y101_SLICE_X92Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeaffaaffaaffaa)
  ) CLBLM_L_X62Y101_SLICE_X93Y101_DLUT (
.I0(CLBLM_R_X63Y101_SLICE_X94Y101_AO6),
.I1(CLBLM_R_X63Y101_SLICE_X94Y101_BQ),
.I2(CLBLM_R_X63Y101_SLICE_X94Y101_BO6),
.I3(CLBLM_L_X62Y101_SLICE_X93Y101_AO5),
.I4(CLBLM_L_X64Y101_SLICE_X96Y101_A5Q),
.I5(CLBLM_L_X62Y103_SLICE_X93Y103_BQ),
.O5(CLBLM_L_X62Y101_SLICE_X93Y101_DO5),
.O6(CLBLM_L_X62Y101_SLICE_X93Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffd555aaaa8000)
  ) CLBLM_L_X62Y101_SLICE_X93Y101_CLUT (
.I0(CLBLM_L_X62Y101_SLICE_X93Y101_AO6),
.I1(CLBLM_L_X62Y102_SLICE_X92Y102_AQ),
.I2(CLBLM_L_X62Y101_SLICE_X92Y101_AQ),
.I3(CLBLM_R_X63Y101_SLICE_X94Y101_BO6),
.I4(CLBLM_L_X62Y101_SLICE_X92Y101_AO6),
.I5(CLBLM_L_X62Y101_SLICE_X93Y101_BO6),
.O5(CLBLM_L_X62Y101_SLICE_X93Y101_CO5),
.O6(CLBLM_L_X62Y101_SLICE_X93Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc022c00000220000)
  ) CLBLM_L_X62Y101_SLICE_X93Y101_BLUT (
.I0(CLBLM_L_X60Y99_SLICE_X90Y99_BQ),
.I1(CLBLM_L_X64Y101_SLICE_X96Y101_BQ),
.I2(CLBLM_L_X60Y99_SLICE_X90Y99_DQ),
.I3(CLBLM_L_X64Y101_SLICE_X96Y101_B5Q),
.I4(CLBLM_L_X62Y102_SLICE_X93Y102_DQ),
.I5(CLBLM_L_X62Y102_SLICE_X93Y102_CQ),
.O5(CLBLM_L_X62Y101_SLICE_X93Y101_BO5),
.O6(CLBLM_L_X62Y101_SLICE_X93Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5a20000000)
  ) CLBLM_L_X62Y101_SLICE_X93Y101_ALUT (
.I0(CLBLM_L_X64Y101_SLICE_X96Y101_A5Q),
.I1(CLBLM_L_X64Y101_SLICE_X96Y101_BQ),
.I2(CLBLM_L_X62Y100_SLICE_X92Y100_AQ),
.I3(CLBLM_L_X62Y103_SLICE_X93Y103_AQ),
.I4(CLBLM_L_X64Y101_SLICE_X96Y101_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X62Y101_SLICE_X93Y101_AO5),
.O6(CLBLM_L_X62Y101_SLICE_X93Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y102_SLICE_X92Y102_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y102_SLICE_X92Y102_AO6),
.Q(CLBLM_L_X62Y102_SLICE_X92Y102_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y102_SLICE_X92Y102_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y102_SLICE_X92Y102_BO6),
.Q(CLBLM_L_X62Y102_SLICE_X92Y102_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y102_SLICE_X92Y102_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y102_SLICE_X92Y102_CO6),
.Q(CLBLM_L_X62Y102_SLICE_X92Y102_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he000a000c0000000)
  ) CLBLM_L_X62Y102_SLICE_X92Y102_DLUT (
.I0(CLBLM_L_X62Y100_SLICE_X92Y100_AQ),
.I1(CLBLM_R_X63Y102_SLICE_X94Y102_BQ),
.I2(CLBLM_L_X64Y101_SLICE_X96Y101_BQ),
.I3(CLBLM_L_X64Y101_SLICE_X96Y101_B5Q),
.I4(CLBLM_L_X62Y103_SLICE_X92Y103_A5Q),
.I5(CLBLM_L_X62Y102_SLICE_X93Y102_BQ),
.O5(CLBLM_L_X62Y102_SLICE_X92Y102_DO5),
.O6(CLBLM_L_X62Y102_SLICE_X92Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaacfaaccaac0aa)
  ) CLBLM_L_X62Y102_SLICE_X92Y102_CLUT (
.I0(CLBLM_L_X62Y102_SLICE_X92Y102_BQ),
.I1(CLBLM_L_X62Y102_SLICE_X92Y102_CQ),
.I2(CLBLM_R_X63Y103_SLICE_X94Y103_AO5),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_R_X63Y102_SLICE_X94Y102_DO6),
.I5(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.O5(CLBLM_L_X62Y102_SLICE_X92Y102_CO5),
.O6(CLBLM_L_X62Y102_SLICE_X92Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccddf0f0cc88f0f0)
  ) CLBLM_L_X62Y102_SLICE_X92Y102_BLUT (
.I0(CLBLM_R_X63Y102_SLICE_X94Y102_DO6),
.I1(CLBLM_L_X62Y102_SLICE_X92Y102_BQ),
.I2(CLBLM_L_X62Y102_SLICE_X92Y102_AQ),
.I3(CLBLM_R_X63Y102_SLICE_X94Y102_DO5),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.O5(CLBLM_L_X62Y102_SLICE_X92Y102_BO5),
.O6(CLBLM_L_X62Y102_SLICE_X92Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f1ff00e0e0ff00)
  ) CLBLM_L_X62Y102_SLICE_X92Y102_ALUT (
.I0(CLBLM_R_X63Y102_SLICE_X94Y102_DO6),
.I1(CLBLM_R_X63Y103_SLICE_X94Y103_AO6),
.I2(CLBLM_L_X62Y102_SLICE_X92Y102_AQ),
.I3(CLBLM_L_X62Y102_SLICE_X93Y102_BQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.O5(CLBLM_L_X62Y102_SLICE_X92Y102_AO5),
.O6(CLBLM_L_X62Y102_SLICE_X92Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y102_SLICE_X93Y102_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y102_SLICE_X93Y102_AO6),
.Q(CLBLM_L_X62Y102_SLICE_X93Y102_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y102_SLICE_X93Y102_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y102_SLICE_X93Y102_BO6),
.Q(CLBLM_L_X62Y102_SLICE_X93Y102_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y102_SLICE_X93Y102_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y102_SLICE_X93Y102_CO6),
.Q(CLBLM_L_X62Y102_SLICE_X93Y102_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y102_SLICE_X93Y102_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y102_SLICE_X93Y102_DO6),
.Q(CLBLM_L_X62Y102_SLICE_X93Y102_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4eee4e4e444)
  ) CLBLM_L_X62Y102_SLICE_X93Y102_DLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X62Y102_SLICE_X93Y102_CQ),
.I2(CLBLM_L_X62Y102_SLICE_X93Y102_DQ),
.I3(CLBLM_R_X63Y103_SLICE_X94Y103_AO5),
.I4(CLBLM_L_X64Y102_SLICE_X96Y102_BO6),
.I5(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.O5(CLBLM_L_X62Y102_SLICE_X93Y102_DO5),
.O6(CLBLM_L_X62Y102_SLICE_X93Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88dd88f5a0)
  ) CLBLM_L_X62Y102_SLICE_X93Y102_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X62Y102_SLICE_X93Y102_CQ),
.I2(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I3(CLBLM_L_X62Y103_SLICE_X93Y103_CQ),
.I4(CLBLM_L_X64Y102_SLICE_X96Y102_BO6),
.I5(CLBLM_R_X63Y102_SLICE_X94Y102_DO5),
.O5(CLBLM_L_X62Y102_SLICE_X93Y102_CO5),
.O6(CLBLM_L_X62Y102_SLICE_X93Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0df8fd080)
  ) CLBLM_L_X62Y102_SLICE_X93Y102_BLUT (
.I0(CLBLM_R_X63Y102_SLICE_X95Y102_AO5),
.I1(CLBLM_L_X62Y102_SLICE_X93Y102_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I4(CLBLM_R_X63Y102_SLICE_X95Y102_BQ),
.I5(CLBLM_R_X63Y102_SLICE_X94Y102_DO6),
.O5(CLBLM_L_X62Y102_SLICE_X93Y102_BO5),
.O6(CLBLM_L_X62Y102_SLICE_X93Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf2f2ff00d0d0ff00)
  ) CLBLM_L_X62Y102_SLICE_X93Y102_ALUT (
.I0(CLBLM_L_X64Y102_SLICE_X96Y102_A5Q),
.I1(CLBLM_L_X64Y102_SLICE_X96Y102_BO6),
.I2(CLBLM_L_X62Y102_SLICE_X93Y102_AQ),
.I3(CLBLM_L_X62Y102_SLICE_X93Y102_DQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.O5(CLBLM_L_X62Y102_SLICE_X93Y102_AO5),
.O6(CLBLM_L_X62Y102_SLICE_X93Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y103_SLICE_X92Y103_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y101_SLICE_X94Y101_AQ),
.Q(CLBLM_L_X62Y103_SLICE_X92Y103_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y103_SLICE_X92Y103_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y103_SLICE_X92Y103_A5Q),
.Q(CLBLM_L_X62Y103_SLICE_X92Y103_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y103_SLICE_X92Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y103_SLICE_X92Y103_AO6),
.Q(CLBLM_L_X62Y103_SLICE_X92Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y103_SLICE_X92Y103_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y103_SLICE_X92Y103_BO6),
.Q(CLBLM_L_X62Y103_SLICE_X92Y103_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y103_SLICE_X92Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y103_SLICE_X92Y103_DO5),
.O6(CLBLM_L_X62Y103_SLICE_X92Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f070f070f0)
  ) CLBLM_L_X62Y103_SLICE_X92Y103_CLUT (
.I0(CLBLM_L_X64Y101_SLICE_X96Y101_B5Q),
.I1(CLBLM_L_X62Y103_SLICE_X92Y103_AQ),
.I2(CLBLM_L_X64Y101_SLICE_X96Y101_A5Q),
.I3(CLBLM_L_X62Y103_SLICE_X92Y103_A5Q),
.I4(1'b1),
.I5(CLBLM_L_X64Y101_SLICE_X96Y101_BQ),
.O5(CLBLM_L_X62Y103_SLICE_X92Y103_CO5),
.O6(CLBLM_L_X62Y103_SLICE_X92Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccfaaaaccc0aaaa)
  ) CLBLM_L_X62Y103_SLICE_X92Y103_BLUT (
.I0(CLBLM_L_X62Y103_SLICE_X92Y103_AQ),
.I1(CLBLM_L_X62Y103_SLICE_X92Y103_BQ),
.I2(CLBLM_R_X63Y102_SLICE_X94Y102_DO5),
.I3(CLBLM_R_X63Y103_SLICE_X95Y103_BO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.O5(CLBLM_L_X62Y103_SLICE_X92Y103_BO5),
.O6(CLBLM_L_X62Y103_SLICE_X92Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aaaaf3c0aaaa)
  ) CLBLM_L_X62Y103_SLICE_X92Y103_ALUT (
.I0(CLBLM_R_X63Y103_SLICE_X95Y103_AQ),
.I1(CLBLM_R_X63Y103_SLICE_X94Y103_AO6),
.I2(CLBLM_L_X62Y103_SLICE_X92Y103_AQ),
.I3(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_R_X63Y103_SLICE_X95Y103_BO6),
.O5(CLBLM_L_X62Y103_SLICE_X92Y103_AO5),
.O6(CLBLM_L_X62Y103_SLICE_X92Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y103_SLICE_X93Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y103_SLICE_X93Y103_AO6),
.Q(CLBLM_L_X62Y103_SLICE_X93Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y103_SLICE_X93Y103_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y103_SLICE_X93Y103_BO6),
.Q(CLBLM_L_X62Y103_SLICE_X93Y103_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y103_SLICE_X93Y103_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y103_SLICE_X93Y103_CO6),
.Q(CLBLM_L_X62Y103_SLICE_X93Y103_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y103_SLICE_X93Y103_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y103_SLICE_X93Y103_DO6),
.Q(CLBLM_L_X62Y103_SLICE_X93Y103_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f7f5d5a0a2a080)
  ) CLBLM_L_X62Y103_SLICE_X93Y103_DLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_R_X63Y103_SLICE_X95Y103_BO6),
.I2(CLBLM_L_X62Y103_SLICE_X93Y103_DQ),
.I3(CLBLM_R_X63Y103_SLICE_X94Y103_AO5),
.I4(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I5(CLBLM_L_X62Y103_SLICE_X92Y103_BQ),
.O5(CLBLM_L_X62Y103_SLICE_X93Y103_DO5),
.O6(CLBLM_L_X62Y103_SLICE_X93Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0df8fd080)
  ) CLBLM_L_X62Y103_SLICE_X93Y103_CLUT (
.I0(CLBLM_L_X64Y102_SLICE_X96Y102_BO6),
.I1(CLBLM_L_X62Y103_SLICE_X93Y103_CQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I4(CLBLM_L_X62Y103_SLICE_X93Y103_AQ),
.I5(CLBLM_R_X63Y103_SLICE_X94Y103_AO6),
.O5(CLBLM_L_X62Y103_SLICE_X93Y103_CO5),
.O6(CLBLM_L_X62Y103_SLICE_X93Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccff00e4e4ff00)
  ) CLBLM_L_X62Y103_SLICE_X93Y103_BLUT (
.I0(CLBLM_L_X64Y102_SLICE_X96Y102_A5Q),
.I1(CLBLM_L_X62Y103_SLICE_X93Y103_BQ),
.I2(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I3(CLBLM_L_X62Y103_SLICE_X93Y103_DQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_R_X63Y103_SLICE_X95Y103_BO6),
.O5(CLBLM_L_X62Y103_SLICE_X93Y103_BO5),
.O6(CLBLM_L_X62Y103_SLICE_X93Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaafccccaaa0cccc)
  ) CLBLM_L_X62Y103_SLICE_X93Y103_ALUT (
.I0(CLBLM_L_X62Y103_SLICE_X93Y103_AQ),
.I1(CLBLM_L_X62Y103_SLICE_X93Y103_BQ),
.I2(CLBLM_L_X64Y102_SLICE_X96Y102_BO6),
.I3(CLBLM_R_X63Y102_SLICE_X95Y102_AO5),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.O5(CLBLM_L_X62Y103_SLICE_X93Y103_AO5),
.O6(CLBLM_L_X62Y103_SLICE_X93Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y105_SLICE_X92Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y105_SLICE_X92Y105_DO5),
.O6(CLBLM_L_X62Y105_SLICE_X92Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y105_SLICE_X92Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y105_SLICE_X92Y105_CO5),
.O6(CLBLM_L_X62Y105_SLICE_X92Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y105_SLICE_X92Y105_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y105_SLICE_X92Y105_BO5),
.O6(CLBLM_L_X62Y105_SLICE_X92Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y105_SLICE_X92Y105_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y105_SLICE_X92Y105_AO5),
.O6(CLBLM_L_X62Y105_SLICE_X92Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y105_SLICE_X93Y105_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X60Y104_SLICE_X90Y104_AQ),
.Q(CLBLM_L_X62Y105_SLICE_X93Y105_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y105_SLICE_X93Y105_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y105_SLICE_X93Y105_AO6),
.Q(CLBLM_L_X62Y105_SLICE_X93Y105_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y105_SLICE_X93Y105_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y105_SLICE_X93Y105_BO6),
.Q(CLBLM_L_X62Y105_SLICE_X93Y105_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y105_SLICE_X93Y105_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y105_SLICE_X93Y105_CO6),
.Q(CLBLM_L_X62Y105_SLICE_X93Y105_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0880088f8008800)
  ) CLBLM_L_X62Y105_SLICE_X93Y105_DLUT (
.I0(CLBLM_R_X63Y105_SLICE_X95Y105_BQ),
.I1(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I2(CLBLM_L_X62Y106_SLICE_X92Y106_BQ),
.I3(CLBLM_R_X63Y105_SLICE_X95Y105_A5Q),
.I4(CLBLM_L_X62Y105_SLICE_X93Y105_AQ),
.I5(CLBLM_L_X62Y107_SLICE_X93Y107_BQ),
.O5(CLBLM_L_X62Y105_SLICE_X93Y105_DO5),
.O6(CLBLM_L_X62Y105_SLICE_X93Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcdc8cdc8ffff0000)
  ) CLBLM_L_X62Y105_SLICE_X93Y105_CLUT (
.I0(CLBLM_L_X64Y106_SLICE_X96Y106_DO5),
.I1(CLBLM_L_X62Y105_SLICE_X93Y105_CQ),
.I2(CLBLM_L_X64Y105_SLICE_X96Y105_BO5),
.I3(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I4(CLBLM_L_X62Y105_SLICE_X93Y105_AQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X62Y105_SLICE_X93Y105_CO5),
.O6(CLBLM_L_X62Y105_SLICE_X93Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00d8ffd800)
  ) CLBLM_L_X62Y105_SLICE_X93Y105_BLUT (
.I0(CLBLM_L_X64Y106_SLICE_X96Y106_DO6),
.I1(CLBLM_L_X62Y105_SLICE_X93Y105_BQ),
.I2(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X62Y107_SLICE_X93Y107_AQ),
.I5(CLBLM_L_X64Y105_SLICE_X96Y105_AO6),
.O5(CLBLM_L_X62Y105_SLICE_X93Y105_BO5),
.O6(CLBLM_L_X62Y105_SLICE_X93Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1e0fffff1e00000)
  ) CLBLM_L_X62Y105_SLICE_X93Y105_ALUT (
.I0(CLBLM_L_X64Y106_SLICE_X96Y106_DO6),
.I1(CLBLM_L_X64Y105_SLICE_X96Y105_BO5),
.I2(CLBLM_L_X62Y105_SLICE_X93Y105_AQ),
.I3(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X62Y106_SLICE_X93Y106_CQ),
.O5(CLBLM_L_X62Y105_SLICE_X93Y105_AO5),
.O6(CLBLM_L_X62Y105_SLICE_X93Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y106_SLICE_X92Y106_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y106_SLICE_X93Y106_AQ),
.Q(CLBLM_L_X62Y106_SLICE_X92Y106_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y106_SLICE_X92Y106_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y106_SLICE_X92Y106_AQ),
.Q(CLBLM_L_X62Y106_SLICE_X92Y106_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8f0f8f0f0f0f0f0f)
  ) CLBLM_L_X62Y106_SLICE_X92Y106_DLUT (
.I0(CLBLM_R_X63Y105_SLICE_X94Y105_C5Q),
.I1(CLBLM_L_X64Y106_SLICE_X96Y106_A5Q),
.I2(CLBLM_R_X63Y105_SLICE_X95Y105_A5Q),
.I3(CLBLM_L_X62Y105_SLICE_X93Y105_CQ),
.I4(1'b1),
.I5(CLBLM_R_X63Y105_SLICE_X94Y105_CQ),
.O5(CLBLM_L_X62Y106_SLICE_X92Y106_DO5),
.O6(CLBLM_L_X62Y106_SLICE_X92Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aaaa000caaae)
  ) CLBLM_L_X62Y106_SLICE_X92Y106_CLUT (
.I0(CLBLM_L_X62Y106_SLICE_X92Y106_AO6),
.I1(CLBLM_R_X63Y106_SLICE_X94Y106_CO6),
.I2(CLBLM_R_X63Y106_SLICE_X95Y106_DO6),
.I3(CLBLM_L_X62Y107_SLICE_X92Y107_AO6),
.I4(CLBLM_L_X62Y106_SLICE_X92Y106_DO6),
.I5(CLBLM_L_X62Y106_SLICE_X92Y106_BO6),
.O5(CLBLM_L_X62Y106_SLICE_X92Y106_CO5),
.O6(CLBLM_L_X62Y106_SLICE_X92Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf800000088000000)
  ) CLBLM_L_X62Y106_SLICE_X92Y106_BLUT (
.I0(CLBLM_L_X64Y106_SLICE_X96Y106_CQ),
.I1(CLBLM_L_X62Y107_SLICE_X93Y107_BQ),
.I2(CLBLM_L_X62Y106_SLICE_X92Y106_AQ),
.I3(CLBLM_R_X63Y105_SLICE_X94Y105_CQ),
.I4(CLBLM_R_X63Y105_SLICE_X94Y105_C5Q),
.I5(CLBLM_R_X63Y107_SLICE_X95Y107_BQ),
.O5(CLBLM_L_X62Y106_SLICE_X92Y106_BO5),
.O6(CLBLM_L_X62Y106_SLICE_X92Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafbbffffffbbff)
  ) CLBLM_L_X62Y106_SLICE_X92Y106_ALUT (
.I0(CLBLM_R_X63Y105_SLICE_X94Y105_CQ),
.I1(CLBLM_L_X64Y106_SLICE_X96Y106_AQ),
.I2(CLBLM_L_X62Y106_SLICE_X92Y106_AQ),
.I3(CLBLM_L_X62Y106_SLICE_X93Y106_AQ),
.I4(CLBLM_R_X63Y105_SLICE_X94Y105_C5Q),
.I5(CLBLM_L_X62Y106_SLICE_X93Y106_CQ),
.O5(CLBLM_L_X62Y106_SLICE_X92Y106_AO5),
.O6(CLBLM_L_X62Y106_SLICE_X92Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y106_SLICE_X93Y106_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X60Y101_SLICE_X90Y101_BQ),
.Q(CLBLM_L_X62Y106_SLICE_X93Y106_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y106_SLICE_X93Y106_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y106_SLICE_X93Y106_BO6),
.Q(CLBLM_L_X62Y106_SLICE_X93Y106_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y106_SLICE_X93Y106_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y106_SLICE_X93Y106_CO6),
.Q(CLBLM_L_X62Y106_SLICE_X93Y106_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaa8aaaaaaaa)
  ) CLBLM_L_X62Y106_SLICE_X93Y106_DLUT (
.I0(CLBLM_L_X64Y105_SLICE_X97Y105_DO6),
.I1(CLBLM_R_X63Y106_SLICE_X94Y106_DO6),
.I2(CLBLM_L_X62Y107_SLICE_X93Y107_DO6),
.I3(CLBLM_L_X62Y106_SLICE_X93Y106_AO5),
.I4(CLBLM_R_X63Y107_SLICE_X94Y107_CO6),
.I5(CLBLM_L_X62Y106_SLICE_X92Y106_CO6),
.O5(CLBLM_L_X62Y106_SLICE_X93Y106_DO5),
.O6(CLBLM_L_X62Y106_SLICE_X93Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccfc0aaaaaaaa)
  ) CLBLM_L_X62Y106_SLICE_X93Y106_CLUT (
.I0(CLBLM_L_X64Y106_SLICE_X96Y106_AQ),
.I1(CLBLM_L_X62Y106_SLICE_X93Y106_CQ),
.I2(CLBLM_L_X64Y106_SLICE_X96Y106_BO5),
.I3(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I4(CLBLM_L_X64Y105_SLICE_X96Y105_BO5),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X62Y106_SLICE_X93Y106_CO5),
.O6(CLBLM_L_X62Y106_SLICE_X93Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdcffdc008cff8c00)
  ) CLBLM_L_X62Y106_SLICE_X93Y106_BLUT (
.I0(CLBLM_L_X64Y105_SLICE_X96Y105_BO5),
.I1(CLBLM_L_X62Y106_SLICE_X93Y106_BQ),
.I2(CLBLM_L_X64Y106_SLICE_X97Y106_C5Q),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X62Y105_SLICE_X93Y105_CQ),
.I5(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.O5(CLBLM_L_X62Y106_SLICE_X93Y106_BO5),
.O6(CLBLM_L_X62Y106_SLICE_X93Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0303030320000000)
  ) CLBLM_L_X62Y106_SLICE_X93Y106_ALUT (
.I0(CLBLM_R_X63Y105_SLICE_X95Y105_A5Q),
.I1(CLBLM_R_X63Y105_SLICE_X94Y105_CQ),
.I2(CLBLM_R_X63Y105_SLICE_X94Y105_C5Q),
.I3(CLBLM_L_X62Y107_SLICE_X93Y107_BQ),
.I4(CLBLM_R_X63Y106_SLICE_X95Y106_BQ),
.I5(1'b1),
.O5(CLBLM_L_X62Y106_SLICE_X93Y106_AO5),
.O6(CLBLM_L_X62Y106_SLICE_X93Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y107_SLICE_X92Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y107_SLICE_X92Y107_DO5),
.O6(CLBLM_L_X62Y107_SLICE_X92Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y107_SLICE_X92Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y107_SLICE_X92Y107_CO5),
.O6(CLBLM_L_X62Y107_SLICE_X92Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd000d0000000d0d0)
  ) CLBLM_L_X62Y107_SLICE_X92Y107_BLUT (
.I0(CLBLM_L_X62Y106_SLICE_X93Y106_AQ),
.I1(CLBLM_L_X60Y101_SLICE_X90Y101_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X62Y107_SLICE_X93Y107_BQ),
.I4(CLBLM_L_X62Y107_SLICE_X93Y107_A5Q),
.I5(CLBLL_R_X75Y107_SLICE_X114Y107_AQ),
.O5(CLBLM_L_X62Y107_SLICE_X92Y107_BO5),
.O6(CLBLM_L_X62Y107_SLICE_X92Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0040aa00aa00)
  ) CLBLM_L_X62Y107_SLICE_X92Y107_ALUT (
.I0(CLBLM_R_X63Y105_SLICE_X94Y105_C5Q),
.I1(CLBLM_R_X63Y107_SLICE_X94Y107_AQ),
.I2(CLBLM_L_X62Y106_SLICE_X92Y106_BQ),
.I3(CLBLM_R_X63Y105_SLICE_X94Y105_CQ),
.I4(CLBLM_R_X63Y105_SLICE_X95Y105_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X62Y107_SLICE_X92Y107_AO5),
.O6(CLBLM_L_X62Y107_SLICE_X92Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y107_SLICE_X93Y107_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y107_SLICE_X114Y107_AQ),
.Q(CLBLM_L_X62Y107_SLICE_X93Y107_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y107_SLICE_X93Y107_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.Q(CLBLM_L_X62Y107_SLICE_X93Y107_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y107_SLICE_X93Y107_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.Q(CLBLM_L_X62Y107_SLICE_X93Y107_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c040c000c000c00)
  ) CLBLM_L_X62Y107_SLICE_X93Y107_DLUT (
.I0(CLBLM_L_X62Y107_SLICE_X93Y107_CO5),
.I1(CLBLM_R_X63Y105_SLICE_X94Y105_CQ),
.I2(CLBLM_R_X63Y105_SLICE_X94Y105_C5Q),
.I3(CLBLM_L_X62Y105_SLICE_X93Y105_DO6),
.I4(CLBLM_L_X62Y107_SLICE_X93Y107_AQ),
.I5(CLBLL_R_X75Y107_SLICE_X114Y107_AQ),
.O5(CLBLM_L_X62Y107_SLICE_X93Y107_DO5),
.O6(CLBLM_L_X62Y107_SLICE_X93Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc00000005a5a5a5a)
  ) CLBLM_L_X62Y107_SLICE_X93Y107_CLUT (
.I0(CLBLM_R_X63Y105_SLICE_X95Y105_A5Q),
.I1(CLBLL_R_X75Y107_SLICE_X114Y107_AQ),
.I2(CLBLM_L_X62Y107_SLICE_X93Y107_BQ),
.I3(CLBLM_L_X62Y107_SLICE_X93Y107_A5Q),
.I4(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I5(1'b1),
.O5(CLBLM_L_X62Y107_SLICE_X93Y107_CO5),
.O6(CLBLM_L_X62Y107_SLICE_X93Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h008044c48080c4c4)
  ) CLBLM_L_X62Y107_SLICE_X93Y107_BLUT (
.I0(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I1(CLBLM_L_X62Y107_SLICE_X92Y107_BO6),
.I2(CLBLM_L_X62Y107_SLICE_X93Y107_A5Q),
.I3(CLBLL_R_X75Y107_SLICE_X114Y107_AQ),
.I4(CLBLM_L_X60Y101_SLICE_X90Y101_BQ),
.I5(CLBLM_L_X62Y107_SLICE_X93Y107_BQ),
.O5(CLBLM_L_X62Y107_SLICE_X93Y107_BO5),
.O6(CLBLM_L_X62Y107_SLICE_X93Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaafccccaaa0cccc)
  ) CLBLM_L_X62Y107_SLICE_X93Y107_ALUT (
.I0(CLBLM_L_X62Y107_SLICE_X93Y107_AQ),
.I1(CLBLM_R_X63Y106_SLICE_X95Y106_BQ),
.I2(CLBLM_L_X64Y106_SLICE_X96Y106_BO5),
.I3(CLBLM_L_X64Y105_SLICE_X96Y105_AO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.O5(CLBLM_L_X62Y107_SLICE_X93Y107_AO5),
.O6(CLBLM_L_X62Y107_SLICE_X93Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y96_SLICE_X96Y96_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y96_SLICE_X96Y96_DO5),
.O6(CLBLM_L_X64Y96_SLICE_X96Y96_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y96_SLICE_X96Y96_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y96_SLICE_X96Y96_CO5),
.O6(CLBLM_L_X64Y96_SLICE_X96Y96_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y96_SLICE_X96Y96_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y96_SLICE_X96Y96_BO5),
.O6(CLBLM_L_X64Y96_SLICE_X96Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y96_SLICE_X96Y96_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y96_SLICE_X96Y96_AO5),
.O6(CLBLM_L_X64Y96_SLICE_X96Y96_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y96_SLICE_X97Y96_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y99_SLICE_X97Y99_A5Q),
.Q(CLBLM_L_X64Y96_SLICE_X97Y96_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y96_SLICE_X97Y96_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y96_SLICE_X97Y96_AO6),
.Q(CLBLM_L_X64Y96_SLICE_X97Y96_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y96_SLICE_X97Y96_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y96_SLICE_X97Y96_DO5),
.O6(CLBLM_L_X64Y96_SLICE_X97Y96_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y96_SLICE_X97Y96_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y96_SLICE_X97Y96_CO5),
.O6(CLBLM_L_X64Y96_SLICE_X97Y96_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y96_SLICE_X97Y96_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y96_SLICE_X97Y96_BO5),
.O6(CLBLM_L_X64Y96_SLICE_X97Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7575757522202220)
  ) CLBLM_L_X64Y96_SLICE_X97Y96_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X64Y97_SLICE_X97Y97_AQ),
.I2(CLBLM_L_X64Y96_SLICE_X97Y96_AQ),
.I3(CLBLM_L_X64Y99_SLICE_X97Y99_A5Q),
.I4(1'b1),
.I5(CLBLM_L_X64Y96_SLICE_X97Y96_A5Q),
.O5(CLBLM_L_X64Y96_SLICE_X97Y96_AO5),
.O6(CLBLM_L_X64Y96_SLICE_X97Y96_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y97_SLICE_X96Y97_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y97_SLICE_X96Y97_AO6),
.Q(CLBLM_L_X64Y97_SLICE_X96Y97_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y97_SLICE_X96Y97_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y97_SLICE_X96Y97_BO6),
.Q(CLBLM_L_X64Y97_SLICE_X96Y97_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y97_SLICE_X96Y97_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y97_SLICE_X96Y97_CO6),
.Q(CLBLM_L_X64Y97_SLICE_X96Y97_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y97_SLICE_X96Y97_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y97_SLICE_X96Y97_DO6),
.Q(CLBLM_L_X64Y97_SLICE_X96Y97_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55fd5daa00a808)
  ) CLBLM_L_X64Y97_SLICE_X96Y97_DLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I2(CLBLM_L_X64Y97_SLICE_X97Y97_BO5),
.I3(CLBLM_L_X64Y97_SLICE_X96Y97_DQ),
.I4(CLBLM_R_X63Y99_SLICE_X94Y99_CO5),
.I5(CLBLM_R_X63Y96_SLICE_X95Y96_CQ),
.O5(CLBLM_L_X64Y97_SLICE_X96Y97_DO5),
.O6(CLBLM_L_X64Y97_SLICE_X96Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccf0ddf088f0)
  ) CLBLM_L_X64Y97_SLICE_X96Y97_CLUT (
.I0(CLBLM_R_X63Y99_SLICE_X94Y99_BO6),
.I1(CLBLM_L_X64Y97_SLICE_X96Y97_CQ),
.I2(CLBLM_R_X63Y97_SLICE_X94Y97_BQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I5(CLBLM_L_X64Y98_SLICE_X96Y98_AO6),
.O5(CLBLM_L_X64Y97_SLICE_X96Y97_CO5),
.O6(CLBLM_L_X64Y97_SLICE_X96Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcecec4c4ff00ff00)
  ) CLBLM_L_X64Y97_SLICE_X96Y97_BLUT (
.I0(CLBLM_R_X63Y99_SLICE_X94Y99_A5Q),
.I1(CLBLM_L_X64Y97_SLICE_X96Y97_BQ),
.I2(CLBLM_L_X64Y97_SLICE_X97Y97_BO5),
.I3(CLBLM_L_X64Y97_SLICE_X96Y97_DQ),
.I4(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X64Y97_SLICE_X96Y97_BO5),
.O6(CLBLM_L_X64Y97_SLICE_X96Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0e2ff00ff00)
  ) CLBLM_L_X64Y97_SLICE_X96Y97_ALUT (
.I0(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I1(CLBLM_R_X63Y99_SLICE_X94Y99_BO6),
.I2(CLBLM_L_X64Y97_SLICE_X96Y97_AQ),
.I3(CLBLM_L_X64Y99_SLICE_X96Y99_BQ),
.I4(CLBLM_L_X64Y99_SLICE_X96Y99_A5Q),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X64Y97_SLICE_X96Y97_AO5),
.O6(CLBLM_L_X64Y97_SLICE_X96Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y97_SLICE_X97Y97_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y97_SLICE_X97Y97_AO5),
.Q(CLBLM_L_X64Y97_SLICE_X97Y97_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y97_SLICE_X97Y97_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y97_SLICE_X97Y97_AO6),
.Q(CLBLM_L_X64Y97_SLICE_X97Y97_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y97_SLICE_X97Y97_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y97_SLICE_X97Y97_CO6),
.Q(CLBLM_L_X64Y97_SLICE_X97Y97_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y97_SLICE_X97Y97_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y97_SLICE_X97Y97_DO6),
.Q(CLBLM_L_X64Y97_SLICE_X97Y97_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0e2e2ff00ff00)
  ) CLBLM_L_X64Y97_SLICE_X97Y97_DLUT (
.I0(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I1(CLBLM_L_X64Y98_SLICE_X96Y98_AO6),
.I2(CLBLM_L_X64Y97_SLICE_X97Y97_DQ),
.I3(CLBLM_R_X63Y96_SLICE_X95Y96_DQ),
.I4(CLBLM_R_X63Y99_SLICE_X94Y99_CO5),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X64Y97_SLICE_X97Y97_DO5),
.O6(CLBLM_L_X64Y97_SLICE_X97Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88ccccf0f0f0f0)
  ) CLBLM_L_X64Y97_SLICE_X97Y97_CLUT (
.I0(CLBLM_L_X64Y98_SLICE_X96Y98_AO6),
.I1(CLBLM_L_X64Y97_SLICE_X97Y97_CQ),
.I2(CLBLM_L_X64Y97_SLICE_X97Y97_DQ),
.I3(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I4(CLBLM_R_X63Y99_SLICE_X94Y99_A5Q),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X64Y97_SLICE_X97Y97_CO5),
.O6(CLBLM_L_X64Y97_SLICE_X97Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddddddeeeeeeee)
  ) CLBLM_L_X64Y97_SLICE_X97Y97_BLUT (
.I0(CLBLM_L_X64Y99_SLICE_X96Y99_A5Q),
.I1(CLBLM_L_X64Y99_SLICE_X96Y99_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y97_SLICE_X97Y97_BO5),
.O6(CLBLM_L_X64Y97_SLICE_X97Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc30307744bb88)
  ) CLBLM_L_X64Y97_SLICE_X97Y97_ALUT (
.I0(CLBLM_R_X63Y98_SLICE_X94Y98_AO5),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_L_X64Y96_SLICE_X97Y96_AQ),
.I3(CLBLM_R_X63Y97_SLICE_X94Y97_CQ),
.I4(CLBLM_L_X64Y97_SLICE_X97Y97_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X64Y97_SLICE_X97Y97_AO5),
.O6(CLBLM_L_X64Y97_SLICE_X97Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y98_SLICE_X96Y98_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y98_SLICE_X96Y98_BO6),
.Q(CLBLM_L_X64Y98_SLICE_X96Y98_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y98_SLICE_X96Y98_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y98_SLICE_X96Y98_DO5),
.O6(CLBLM_L_X64Y98_SLICE_X96Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h153faaff3f3fffff)
  ) CLBLM_L_X64Y98_SLICE_X96Y98_CLUT (
.I0(CLBLM_L_X62Y99_SLICE_X93Y99_AQ),
.I1(CLBLM_R_X63Y97_SLICE_X94Y97_AQ),
.I2(CLBLM_R_X63Y96_SLICE_X95Y96_CQ),
.I3(CLBLM_L_X76Y111_SLICE_X116Y111_BQ),
.I4(CLBLM_L_X64Y97_SLICE_X97Y97_A5Q),
.I5(CLBLM_R_X63Y96_SLICE_X94Y96_BQ),
.O5(CLBLM_L_X64Y98_SLICE_X96Y98_CO5),
.O6(CLBLM_L_X64Y98_SLICE_X96Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8d8d8d8fad850)
  ) CLBLM_L_X64Y98_SLICE_X96Y98_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X64Y98_SLICE_X96Y98_BQ),
.I2(CLBLM_L_X64Y97_SLICE_X97Y97_CQ),
.I3(CLBLM_R_X63Y99_SLICE_X94Y99_BO6),
.I4(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I5(CLBLM_L_X64Y98_SLICE_X96Y98_AO5),
.O5(CLBLM_L_X64Y98_SLICE_X96Y98_BO5),
.O6(CLBLM_L_X64Y98_SLICE_X96Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbbbbb77777777)
  ) CLBLM_L_X64Y98_SLICE_X96Y98_ALUT (
.I0(CLBLM_L_X64Y99_SLICE_X96Y99_A5Q),
.I1(CLBLM_L_X64Y99_SLICE_X96Y99_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y98_SLICE_X96Y98_AO5),
.O6(CLBLM_L_X64Y98_SLICE_X96Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y98_SLICE_X97Y98_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y98_SLICE_X97Y98_DO5),
.O6(CLBLM_L_X64Y98_SLICE_X97Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y98_SLICE_X97Y98_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y98_SLICE_X97Y98_CO5),
.O6(CLBLM_L_X64Y98_SLICE_X97Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y98_SLICE_X97Y98_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y98_SLICE_X97Y98_BO5),
.O6(CLBLM_L_X64Y98_SLICE_X97Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y98_SLICE_X97Y98_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y98_SLICE_X97Y98_AO5),
.O6(CLBLM_L_X64Y98_SLICE_X97Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y99_SLICE_X96Y99_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y99_SLICE_X96Y99_AO5),
.Q(CLBLM_L_X64Y99_SLICE_X96Y99_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y99_SLICE_X96Y99_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y99_SLICE_X96Y99_AO6),
.Q(CLBLM_L_X64Y99_SLICE_X96Y99_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y99_SLICE_X96Y99_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y99_SLICE_X96Y99_BO6),
.Q(CLBLM_L_X64Y99_SLICE_X96Y99_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y99_SLICE_X96Y99_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y99_SLICE_X96Y99_CO6),
.Q(CLBLM_L_X64Y99_SLICE_X96Y99_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y99_SLICE_X96Y99_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y99_SLICE_X96Y99_DO5),
.O6(CLBLM_L_X64Y99_SLICE_X96Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ccccaaaaaaaa)
  ) CLBLM_L_X64Y99_SLICE_X96Y99_CLUT (
.I0(CLBLM_L_X62Y98_SLICE_X93Y98_CQ),
.I1(CLBLM_L_X64Y99_SLICE_X96Y99_CQ),
.I2(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I3(1'b1),
.I4(CLBLM_L_X64Y99_SLICE_X96Y99_BO5),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X64Y99_SLICE_X96Y99_CO5),
.O6(CLBLM_L_X64Y99_SLICE_X96Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h66ffcc0088880000)
  ) CLBLM_L_X64Y99_SLICE_X96Y99_BLUT (
.I0(CLBLM_R_X63Y99_SLICE_X94Y99_A5Q),
.I1(CLBLM_L_X64Y99_SLICE_X96Y99_BQ),
.I2(1'b1),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X64Y99_SLICE_X96Y99_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X64Y99_SLICE_X96Y99_BO5),
.O6(CLBLM_L_X64Y99_SLICE_X96Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0500050066aa66aa)
  ) CLBLM_L_X64Y99_SLICE_X96Y99_ALUT (
.I0(CLBLM_R_X63Y99_SLICE_X94Y99_A5Q),
.I1(CLBLM_L_X64Y99_SLICE_X96Y99_A5Q),
.I2(CLBLM_L_X64Y99_SLICE_X96Y99_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y99_SLICE_X96Y99_AO5),
.O6(CLBLM_L_X64Y99_SLICE_X96Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y99_SLICE_X97Y99_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y99_SLICE_X97Y99_AO5),
.Q(CLBLM_L_X64Y99_SLICE_X97Y99_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y99_SLICE_X97Y99_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y99_SLICE_X97Y99_BO5),
.Q(CLBLM_L_X64Y99_SLICE_X97Y99_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y99_SLICE_X97Y99_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y99_SLICE_X97Y99_AO6),
.Q(CLBLM_L_X64Y99_SLICE_X97Y99_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y99_SLICE_X97Y99_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y99_SLICE_X97Y99_BO6),
.Q(CLBLM_L_X64Y99_SLICE_X97Y99_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y99_SLICE_X97Y99_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y99_SLICE_X97Y99_DO5),
.O6(CLBLM_L_X64Y99_SLICE_X97Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y99_SLICE_X97Y99_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y99_SLICE_X97Y99_CO5),
.O6(CLBLM_L_X64Y99_SLICE_X97Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cf0ccf06accaacc)
  ) CLBLM_L_X64Y99_SLICE_X97Y99_BLUT (
.I0(CLBLM_L_X64Y99_SLICE_X97Y99_B5Q),
.I1(CLBLM_L_X64Y99_SLICE_X97Y99_BQ),
.I2(CLBLM_L_X64Y99_SLICE_X97Y99_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_R_X65Y99_SLICE_X99Y99_DQ),
.I5(1'b1),
.O5(CLBLM_L_X64Y99_SLICE_X97Y99_BO5),
.O6(CLBLM_L_X64Y99_SLICE_X97Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a6a6a6acc00cc00)
  ) CLBLM_L_X64Y99_SLICE_X97Y99_ALUT (
.I0(CLBLM_R_X65Y99_SLICE_X99Y99_DQ),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_L_X64Y99_SLICE_X97Y99_AQ),
.I3(CLBLM_L_X64Y99_SLICE_X96Y99_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y99_SLICE_X97Y99_AO5),
.O6(CLBLM_L_X64Y99_SLICE_X97Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y100_SLICE_X96Y100_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y100_SLICE_X96Y100_DO5),
.O6(CLBLM_L_X64Y100_SLICE_X96Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y100_SLICE_X96Y100_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y100_SLICE_X96Y100_CO5),
.O6(CLBLM_L_X64Y100_SLICE_X96Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y100_SLICE_X96Y100_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y100_SLICE_X96Y100_BO5),
.O6(CLBLM_L_X64Y100_SLICE_X96Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y100_SLICE_X96Y100_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y100_SLICE_X96Y100_AO5),
.O6(CLBLM_L_X64Y100_SLICE_X96Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y100_SLICE_X97Y100_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y100_SLICE_X97Y100_AO6),
.Q(CLBLM_L_X64Y100_SLICE_X97Y100_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y100_SLICE_X97Y100_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y100_SLICE_X97Y100_DO5),
.O6(CLBLM_L_X64Y100_SLICE_X97Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y100_SLICE_X97Y100_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y100_SLICE_X97Y100_CO5),
.O6(CLBLM_L_X64Y100_SLICE_X97Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y100_SLICE_X97Y100_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y100_SLICE_X97Y100_BO5),
.O6(CLBLM_L_X64Y100_SLICE_X97Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500ffaaf5a0)
  ) CLBLM_L_X64Y100_SLICE_X97Y100_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(1'b1),
.I2(CLBLM_L_X64Y100_SLICE_X97Y100_AQ),
.I3(CLBLM_L_X64Y99_SLICE_X96Y99_CQ),
.I4(CLBLM_R_X63Y98_SLICE_X95Y98_AO6),
.I5(CLBLM_L_X64Y103_SLICE_X97Y103_CO6),
.O5(CLBLM_L_X64Y100_SLICE_X97Y100_AO5),
.O6(CLBLM_L_X64Y100_SLICE_X97Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y101_SLICE_X96Y101_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y101_SLICE_X96Y101_AO5),
.Q(CLBLM_L_X64Y101_SLICE_X96Y101_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y101_SLICE_X96Y101_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y101_SLICE_X96Y101_BO5),
.Q(CLBLM_L_X64Y101_SLICE_X96Y101_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y101_SLICE_X96Y101_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y101_SLICE_X96Y101_CO5),
.Q(CLBLM_L_X64Y101_SLICE_X96Y101_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y101_SLICE_X96Y101_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y101_SLICE_X96Y101_AO6),
.Q(CLBLM_L_X64Y101_SLICE_X96Y101_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y101_SLICE_X96Y101_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y101_SLICE_X96Y101_BO6),
.Q(CLBLM_L_X64Y101_SLICE_X96Y101_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y101_SLICE_X96Y101_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y101_SLICE_X96Y101_CO6),
.Q(CLBLM_L_X64Y101_SLICE_X96Y101_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y101_SLICE_X96Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y101_SLICE_X96Y101_DO5),
.O6(CLBLM_L_X64Y101_SLICE_X96Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h050fff0044cccccc)
  ) CLBLM_L_X64Y101_SLICE_X96Y101_CLUT (
.I0(CLBLM_L_X62Y100_SLICE_X93Y100_AO6),
.I1(CLBLM_L_X64Y101_SLICE_X96Y101_CQ),
.I2(CLBLM_L_X64Y101_SLICE_X96Y101_C5Q),
.I3(CLBLM_L_X64Y101_SLICE_X96Y101_A5Q),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLM_L_X64Y101_SLICE_X96Y101_CO5),
.O6(CLBLM_L_X64Y101_SLICE_X96Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6aca6aca5faf50a0)
  ) CLBLM_L_X64Y101_SLICE_X96Y101_BLUT (
.I0(CLBLM_L_X64Y101_SLICE_X96Y101_B5Q),
.I1(CLBLM_L_X64Y101_SLICE_X96Y101_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X64Y103_SLICE_X97Y103_DO6),
.I4(CLBLM_L_X64Y101_SLICE_X96Y101_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X64Y101_SLICE_X96Y101_BO5),
.O6(CLBLM_L_X64Y101_SLICE_X96Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc00cc0faaf0aa)
  ) CLBLM_L_X64Y101_SLICE_X96Y101_ALUT (
.I0(CLBLM_R_X63Y101_SLICE_X94Y101_BQ),
.I1(CLBLM_L_X68Y101_SLICE_X102Y101_AQ),
.I2(CLBLM_L_X62Y100_SLICE_X93Y100_AO6),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X64Y101_SLICE_X96Y101_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X64Y101_SLICE_X96Y101_AO5),
.O6(CLBLM_L_X64Y101_SLICE_X96Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y101_SLICE_X97Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y101_SLICE_X97Y101_DO5),
.O6(CLBLM_L_X64Y101_SLICE_X97Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y101_SLICE_X97Y101_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y101_SLICE_X97Y101_CO5),
.O6(CLBLM_L_X64Y101_SLICE_X97Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y101_SLICE_X97Y101_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y101_SLICE_X97Y101_BO5),
.O6(CLBLM_L_X64Y101_SLICE_X97Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y101_SLICE_X97Y101_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y101_SLICE_X97Y101_AO5),
.O6(CLBLM_L_X64Y101_SLICE_X97Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y102_SLICE_X96Y102_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y102_SLICE_X96Y102_AO5),
.Q(CLBLM_L_X64Y102_SLICE_X96Y102_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y102_SLICE_X96Y102_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y102_SLICE_X96Y102_AO6),
.Q(CLBLM_L_X64Y102_SLICE_X96Y102_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y102_SLICE_X96Y102_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y102_SLICE_X96Y102_CO6),
.Q(CLBLM_L_X64Y102_SLICE_X96Y102_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffa599ffff0000)
  ) CLBLM_L_X64Y102_SLICE_X96Y102_DLUT (
.I0(CLBLM_L_X64Y101_SLICE_X96Y101_BQ),
.I1(CLBLM_L_X64Y101_SLICE_X96Y101_CQ),
.I2(CLBLM_L_X64Y101_SLICE_X96Y101_C5Q),
.I3(CLBLM_L_X64Y101_SLICE_X96Y101_B5Q),
.I4(CLBLM_L_X64Y102_SLICE_X97Y102_BQ),
.I5(CLBLM_L_X64Y103_SLICE_X97Y103_DO6),
.O5(CLBLM_L_X64Y102_SLICE_X96Y102_DO5),
.O6(CLBLM_L_X64Y102_SLICE_X96Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ddf0ccf088f0)
  ) CLBLM_L_X64Y102_SLICE_X96Y102_CLUT (
.I0(CLBLM_R_X63Y102_SLICE_X94Y102_DO5),
.I1(CLBLM_L_X64Y102_SLICE_X96Y102_CQ),
.I2(CLBLM_R_X63Y102_SLICE_X94Y102_BQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X64Y102_SLICE_X96Y102_BO5),
.I5(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.O5(CLBLM_L_X64Y102_SLICE_X96Y102_CO5),
.O6(CLBLM_L_X64Y102_SLICE_X96Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f5f5afafafaf)
  ) CLBLM_L_X64Y102_SLICE_X96Y102_BLUT (
.I0(CLBLM_L_X64Y105_SLICE_X96Y105_CQ),
.I1(1'b1),
.I2(CLBLM_L_X64Y105_SLICE_X96Y105_C5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y102_SLICE_X96Y102_BO5),
.O6(CLBLM_L_X64Y102_SLICE_X96Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aaa5aaa20f020f0)
  ) CLBLM_L_X64Y102_SLICE_X96Y102_ALUT (
.I0(CLBLM_R_X63Y102_SLICE_X95Y102_AQ),
.I1(CLBLM_L_X64Y102_SLICE_X96Y102_A5Q),
.I2(CLBLM_L_X64Y102_SLICE_X96Y102_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y102_SLICE_X96Y102_AO5),
.O6(CLBLM_L_X64Y102_SLICE_X96Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y102_SLICE_X97Y102_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y102_SLICE_X97Y102_AO6),
.Q(CLBLM_L_X64Y102_SLICE_X97Y102_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y102_SLICE_X97Y102_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y102_SLICE_X97Y102_BO6),
.Q(CLBLM_L_X64Y102_SLICE_X97Y102_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y102_SLICE_X97Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y102_SLICE_X97Y102_DO5),
.O6(CLBLM_L_X64Y102_SLICE_X97Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y102_SLICE_X97Y102_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y102_SLICE_X97Y102_CO5),
.O6(CLBLM_L_X64Y102_SLICE_X97Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h08aa000000aa0000)
  ) CLBLM_L_X64Y102_SLICE_X97Y102_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_R_X65Y104_SLICE_X98Y104_CQ),
.I2(CLBLM_R_X65Y104_SLICE_X98Y104_C5Q),
.I3(CLBLM_L_X64Y103_SLICE_X97Y103_DO6),
.I4(CLBLM_L_X64Y102_SLICE_X96Y102_DO6),
.I5(CLBLM_R_X65Y104_SLICE_X99Y104_DO6),
.O5(CLBLM_L_X64Y102_SLICE_X97Y102_BO5),
.O6(CLBLM_L_X64Y102_SLICE_X97Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h20000000f000f000)
  ) CLBLM_L_X64Y102_SLICE_X97Y102_ALUT (
.I0(CLBLM_R_X65Y104_SLICE_X99Y104_DO6),
.I1(CLBLM_R_X65Y104_SLICE_X98Y104_CQ),
.I2(CLBLM_R_X63Y99_SLICE_X95Y99_CO6),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_R_X65Y104_SLICE_X98Y104_C5Q),
.I5(CLBLM_L_X64Y103_SLICE_X97Y103_CO6),
.O5(CLBLM_L_X64Y102_SLICE_X97Y102_AO5),
.O6(CLBLM_L_X64Y102_SLICE_X97Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y103_SLICE_X96Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y103_SLICE_X96Y103_AO6),
.Q(CLBLM_L_X64Y103_SLICE_X96Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y103_SLICE_X96Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y103_SLICE_X96Y103_DO5),
.O6(CLBLM_L_X64Y103_SLICE_X96Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y103_SLICE_X96Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y103_SLICE_X96Y103_CO5),
.O6(CLBLM_L_X64Y103_SLICE_X96Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y103_SLICE_X96Y103_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y103_SLICE_X96Y103_BO5),
.O6(CLBLM_L_X64Y103_SLICE_X96Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaffaa30aa30aa)
  ) CLBLM_L_X64Y103_SLICE_X96Y103_ALUT (
.I0(CLBLM_R_X63Y102_SLICE_X95Y102_DQ),
.I1(CLBLM_L_X64Y103_SLICE_X97Y103_DO6),
.I2(CLBLM_L_X64Y103_SLICE_X96Y103_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(1'b1),
.I5(CLBLM_R_X63Y101_SLICE_X94Y101_DO6),
.O5(CLBLM_L_X64Y103_SLICE_X96Y103_AO5),
.O6(CLBLM_L_X64Y103_SLICE_X96Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y103_SLICE_X97Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y103_SLICE_X97Y103_AO6),
.Q(CLBLM_L_X64Y103_SLICE_X97Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y103_SLICE_X97Y103_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y103_SLICE_X97Y103_BO6),
.Q(CLBLM_L_X64Y103_SLICE_X97Y103_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f007f00ff00ff00)
  ) CLBLM_L_X64Y103_SLICE_X97Y103_DLUT (
.I0(CLBLM_R_X65Y104_SLICE_X98Y104_CQ),
.I1(CLBLM_R_X65Y104_SLICE_X98Y104_C5Q),
.I2(CLBLM_L_X64Y103_SLICE_X97Y103_BQ),
.I3(CLBLM_R_X65Y103_SLICE_X98Y103_A5Q),
.I4(1'b1),
.I5(CLBLM_R_X65Y103_SLICE_X99Y103_CO6),
.O5(CLBLM_L_X64Y103_SLICE_X97Y103_DO5),
.O6(CLBLM_L_X64Y103_SLICE_X97Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbff0000ffff0000)
  ) CLBLM_L_X64Y103_SLICE_X97Y103_CLUT (
.I0(CLBLM_R_X65Y104_SLICE_X98Y104_C5Q),
.I1(CLBLM_R_X65Y103_SLICE_X99Y103_CO6),
.I2(1'b1),
.I3(CLBLM_L_X64Y103_SLICE_X97Y103_AQ),
.I4(CLBLM_R_X65Y104_SLICE_X99Y104_B5Q),
.I5(CLBLM_R_X65Y104_SLICE_X98Y104_CQ),
.O5(CLBLM_L_X64Y103_SLICE_X97Y103_CO5),
.O6(CLBLM_L_X64Y103_SLICE_X97Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcf4fc3030b030)
  ) CLBLM_L_X64Y103_SLICE_X97Y103_BLUT (
.I0(CLBLM_R_X65Y104_SLICE_X99Y104_DO6),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_L_X64Y102_SLICE_X97Y102_BQ),
.I3(CLBLM_R_X65Y104_SLICE_X98Y104_CQ),
.I4(CLBLM_R_X65Y104_SLICE_X98Y104_C5Q),
.I5(CLBLM_L_X64Y103_SLICE_X97Y103_BQ),
.O5(CLBLM_L_X64Y103_SLICE_X97Y103_BO5),
.O6(CLBLM_L_X64Y103_SLICE_X97Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafefa020afafa0a0)
  ) CLBLM_L_X64Y103_SLICE_X97Y103_ALUT (
.I0(CLBLM_L_X64Y103_SLICE_X97Y103_AQ),
.I1(CLBLM_R_X65Y104_SLICE_X99Y104_DO6),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_R_X65Y104_SLICE_X98Y104_CQ),
.I4(CLBLM_L_X64Y102_SLICE_X97Y102_AQ),
.I5(CLBLM_R_X65Y104_SLICE_X98Y104_C5Q),
.O5(CLBLM_L_X64Y103_SLICE_X97Y103_AO5),
.O6(CLBLM_L_X64Y103_SLICE_X97Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y104_SLICE_X96Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y104_SLICE_X96Y104_AO6),
.Q(CLBLM_L_X64Y104_SLICE_X96Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y104_SLICE_X96Y104_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y104_SLICE_X96Y104_BO6),
.Q(CLBLM_L_X64Y104_SLICE_X96Y104_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y104_SLICE_X96Y104_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y104_SLICE_X96Y104_CO6),
.Q(CLBLM_L_X64Y104_SLICE_X96Y104_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y104_SLICE_X96Y104_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y104_SLICE_X96Y104_DO6),
.Q(CLBLM_L_X64Y104_SLICE_X96Y104_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h408cc00cc00cc00c)
  ) CLBLM_L_X64Y104_SLICE_X96Y104_DLUT (
.I0(CLBLM_L_X64Y105_SLICE_X96Y105_C5Q),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_L_X64Y104_SLICE_X96Y104_DQ),
.I3(CLBLL_R_X79Y99_SLICE_X122Y99_AO6),
.I4(CLBLM_L_X64Y105_SLICE_X96Y105_CQ),
.I5(CLBLM_L_X64Y102_SLICE_X96Y102_A5Q),
.O5(CLBLM_L_X64Y104_SLICE_X96Y104_DO5),
.O6(CLBLM_L_X64Y104_SLICE_X96Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5dfd5dfda808a808)
  ) CLBLM_L_X64Y104_SLICE_X96Y104_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X64Y104_SLICE_X96Y104_CQ),
.I2(CLBLM_R_X63Y101_SLICE_X94Y101_BO5),
.I3(CLBLM_L_X64Y104_SLICE_X96Y104_BQ),
.I4(1'b1),
.I5(CLBLM_L_X64Y104_SLICE_X96Y104_AQ),
.O5(CLBLM_L_X64Y104_SLICE_X96Y104_CO5),
.O6(CLBLM_L_X64Y104_SLICE_X96Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hecccffff4ccc0000)
  ) CLBLM_L_X64Y104_SLICE_X96Y104_BLUT (
.I0(CLBLM_L_X64Y105_SLICE_X96Y105_CQ),
.I1(CLBLM_L_X64Y104_SLICE_X96Y104_BQ),
.I2(CLBLM_L_X64Y105_SLICE_X96Y105_C5Q),
.I3(CLBLM_L_X64Y102_SLICE_X96Y102_A5Q),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X64Y104_SLICE_X96Y104_DQ),
.O5(CLBLM_L_X64Y104_SLICE_X96Y104_BO5),
.O6(CLBLM_L_X64Y104_SLICE_X96Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafcccc5050cccc)
  ) CLBLM_L_X64Y104_SLICE_X96Y104_ALUT (
.I0(CLBLM_R_X63Y101_SLICE_X94Y101_BO5),
.I1(CLBLM_L_X64Y104_SLICE_X96Y104_BQ),
.I2(CLBLM_L_X64Y104_SLICE_X96Y104_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_R_X63Y101_SLICE_X94Y101_DO6),
.O5(CLBLM_L_X64Y104_SLICE_X96Y104_AO5),
.O6(CLBLM_L_X64Y104_SLICE_X96Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y104_SLICE_X97Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y104_SLICE_X97Y104_AO6),
.Q(CLBLM_L_X64Y104_SLICE_X97Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y104_SLICE_X97Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y104_SLICE_X97Y104_DO5),
.O6(CLBLM_L_X64Y104_SLICE_X97Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y104_SLICE_X97Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y104_SLICE_X97Y104_CO5),
.O6(CLBLM_L_X64Y104_SLICE_X97Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y104_SLICE_X97Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y104_SLICE_X97Y104_BO5),
.O6(CLBLM_L_X64Y104_SLICE_X97Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcce4e4e4e4e4e4e4)
  ) CLBLM_L_X64Y104_SLICE_X97Y104_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_R_X65Y105_SLICE_X99Y105_C5Q),
.I2(CLBLM_L_X64Y104_SLICE_X97Y104_AQ),
.I3(CLBLM_L_X64Y105_SLICE_X96Y105_CQ),
.I4(CLBLM_L_X64Y105_SLICE_X96Y105_C5Q),
.I5(CLBLM_L_X64Y102_SLICE_X96Y102_A5Q),
.O5(CLBLM_L_X64Y104_SLICE_X97Y104_AO5),
.O6(CLBLM_L_X64Y104_SLICE_X97Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y105_SLICE_X96Y105_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y105_SLICE_X96Y105_CO5),
.Q(CLBLM_L_X64Y105_SLICE_X96Y105_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y105_SLICE_X96Y105_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y105_SLICE_X96Y105_CO6),
.Q(CLBLM_L_X64Y105_SLICE_X96Y105_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y105_SLICE_X96Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y105_SLICE_X96Y105_DO5),
.O6(CLBLM_L_X64Y105_SLICE_X96Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3fc03fc06cac6cac)
  ) CLBLM_L_X64Y105_SLICE_X96Y105_CLUT (
.I0(CLBLM_L_X64Y105_SLICE_X96Y105_C5Q),
.I1(CLBLM_L_X64Y105_SLICE_X96Y105_CQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X64Y102_SLICE_X96Y102_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y105_SLICE_X96Y105_CO5),
.O6(CLBLM_L_X64Y105_SLICE_X96Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5f5ffafafafa)
  ) CLBLM_L_X64Y105_SLICE_X96Y105_BLUT (
.I0(CLBLM_L_X64Y106_SLICE_X97Y106_B5Q),
.I1(1'b1),
.I2(CLBLM_L_X64Y106_SLICE_X97Y106_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y105_SLICE_X96Y105_BO5),
.O6(CLBLM_L_X64Y105_SLICE_X96Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f5f5afafafaf)
  ) CLBLM_L_X64Y105_SLICE_X96Y105_ALUT (
.I0(CLBLM_L_X64Y106_SLICE_X97Y106_B5Q),
.I1(1'b1),
.I2(CLBLM_L_X64Y106_SLICE_X97Y106_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y105_SLICE_X96Y105_AO5),
.O6(CLBLM_L_X64Y105_SLICE_X96Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y105_SLICE_X97Y105_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y105_SLICE_X97Y105_AO6),
.Q(CLBLM_L_X64Y105_SLICE_X97Y105_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y105_SLICE_X97Y105_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y105_SLICE_X97Y105_BO6),
.Q(CLBLM_L_X64Y105_SLICE_X97Y105_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y105_SLICE_X97Y105_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y105_SLICE_X97Y105_CO6),
.Q(CLBLM_L_X64Y105_SLICE_X97Y105_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaaaaa22aa)
  ) CLBLM_L_X64Y105_SLICE_X97Y105_DLUT (
.I0(CLBLM_R_X65Y105_SLICE_X98Y105_AQ),
.I1(CLBLM_R_X65Y103_SLICE_X99Y103_CO6),
.I2(1'b1),
.I3(CLBLM_L_X64Y105_SLICE_X97Y105_AQ),
.I4(CLBLM_R_X65Y104_SLICE_X98Y104_C5Q),
.I5(CLBLM_R_X65Y104_SLICE_X98Y104_CQ),
.O5(CLBLM_L_X64Y105_SLICE_X97Y105_DO5),
.O6(CLBLM_L_X64Y105_SLICE_X97Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7ddddddd28888888)
  ) CLBLM_L_X64Y105_SLICE_X97Y105_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X64Y105_SLICE_X97Y105_CQ),
.I2(CLBLM_L_X64Y105_SLICE_X96Y105_C5Q),
.I3(CLBLM_L_X64Y105_SLICE_X96Y105_CQ),
.I4(CLBLM_L_X64Y102_SLICE_X96Y102_A5Q),
.I5(CLBLM_L_X64Y104_SLICE_X96Y104_CQ),
.O5(CLBLM_L_X64Y105_SLICE_X97Y105_CO5),
.O6(CLBLM_L_X64Y105_SLICE_X97Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h80ff000000000000)
  ) CLBLM_L_X64Y105_SLICE_X97Y105_BLUT (
.I0(CLBLM_R_X65Y104_SLICE_X99Y104_DO6),
.I1(CLBLM_R_X65Y104_SLICE_X98Y104_CQ),
.I2(CLBLM_R_X65Y104_SLICE_X98Y104_C5Q),
.I3(CLBLM_L_X64Y105_SLICE_X97Y105_DO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_R_X63Y105_SLICE_X95Y105_DO6),
.O5(CLBLM_L_X64Y105_SLICE_X97Y105_BO5),
.O6(CLBLM_L_X64Y105_SLICE_X97Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcce4e4e4e4e4e4e4)
  ) CLBLM_L_X64Y105_SLICE_X97Y105_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X64Y105_SLICE_X97Y105_BQ),
.I2(CLBLM_L_X64Y105_SLICE_X97Y105_AQ),
.I3(CLBLM_R_X65Y104_SLICE_X98Y104_CQ),
.I4(CLBLM_R_X65Y104_SLICE_X98Y104_C5Q),
.I5(CLBLM_R_X65Y104_SLICE_X99Y104_DO6),
.O5(CLBLM_L_X64Y105_SLICE_X97Y105_AO5),
.O6(CLBLM_L_X64Y105_SLICE_X97Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y106_SLICE_X96Y106_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y106_SLICE_X92Y106_BQ),
.Q(CLBLM_L_X64Y106_SLICE_X96Y106_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y106_SLICE_X96Y106_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y106_SLICE_X96Y106_AO6),
.Q(CLBLM_L_X64Y106_SLICE_X96Y106_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y106_SLICE_X96Y106_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y106_SLICE_X96Y106_A5Q),
.Q(CLBLM_L_X64Y106_SLICE_X96Y106_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y106_SLICE_X96Y106_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y106_SLICE_X96Y106_CO6),
.Q(CLBLM_L_X64Y106_SLICE_X96Y106_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffccff33ff33ff)
  ) CLBLM_L_X64Y106_SLICE_X96Y106_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X64Y106_SLICE_X97Y106_BQ),
.I2(1'b1),
.I3(CLBLM_L_X64Y106_SLICE_X97Y106_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y106_SLICE_X96Y106_DO5),
.O6(CLBLM_L_X64Y106_SLICE_X96Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00d8ffd800)
  ) CLBLM_L_X64Y106_SLICE_X96Y106_CLUT (
.I0(CLBLM_L_X64Y105_SLICE_X96Y105_BO6),
.I1(CLBLM_L_X64Y106_SLICE_X96Y106_CQ),
.I2(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_R_X63Y106_SLICE_X95Y106_CQ),
.I5(CLBLM_L_X64Y106_SLICE_X96Y106_BO6),
.O5(CLBLM_L_X64Y106_SLICE_X96Y106_CO5),
.O6(CLBLM_L_X64Y106_SLICE_X96Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff0ffff00ff)
  ) CLBLM_L_X64Y106_SLICE_X96Y106_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X64Y106_SLICE_X97Y106_C5Q),
.I3(CLBLM_L_X64Y106_SLICE_X97Y106_BQ),
.I4(CLBLM_L_X64Y106_SLICE_X97Y106_CQ),
.I5(1'b1),
.O5(CLBLM_L_X64Y106_SLICE_X96Y106_BO5),
.O6(CLBLM_L_X64Y106_SLICE_X96Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0e2ffff0000)
  ) CLBLM_L_X64Y106_SLICE_X96Y106_ALUT (
.I0(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I1(CLBLM_L_X64Y106_SLICE_X97Y106_B5Q),
.I2(CLBLM_L_X64Y106_SLICE_X96Y106_AQ),
.I3(CLBLM_L_X64Y106_SLICE_X96Y106_BO6),
.I4(CLBLM_L_X64Y106_SLICE_X97Y106_AQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X64Y106_SLICE_X96Y106_AO5),
.O6(CLBLM_L_X64Y106_SLICE_X96Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y106_SLICE_X97Y106_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y106_SLICE_X97Y106_BO5),
.Q(CLBLM_L_X64Y106_SLICE_X97Y106_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y106_SLICE_X97Y106_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y106_SLICE_X97Y106_CO5),
.Q(CLBLM_L_X64Y106_SLICE_X97Y106_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y106_SLICE_X97Y106_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y106_SLICE_X97Y106_AO5),
.Q(CLBLM_L_X64Y106_SLICE_X97Y106_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y106_SLICE_X97Y106_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y106_SLICE_X97Y106_BO6),
.Q(CLBLM_L_X64Y106_SLICE_X97Y106_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y106_SLICE_X97Y106_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y106_SLICE_X97Y106_CO6),
.Q(CLBLM_L_X64Y106_SLICE_X97Y106_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y106_SLICE_X97Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y106_SLICE_X97Y106_DO5),
.O6(CLBLM_L_X64Y106_SLICE_X97Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cf03cf040cc40cc)
  ) CLBLM_L_X64Y106_SLICE_X97Y106_CLUT (
.I0(CLBLM_L_X64Y106_SLICE_X97Y106_C5Q),
.I1(CLBLM_L_X64Y106_SLICE_X97Y106_CQ),
.I2(CLBLM_L_X64Y106_SLICE_X97Y106_BQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y106_SLICE_X97Y106_CO5),
.O6(CLBLM_L_X64Y106_SLICE_X97Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000030305f5fa0a0)
  ) CLBLM_L_X64Y106_SLICE_X97Y106_BLUT (
.I0(CLBLM_L_X64Y106_SLICE_X97Y106_B5Q),
.I1(CLBLM_L_X64Y106_SLICE_X97Y106_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(1'b1),
.I4(CLBLM_L_X64Y106_SLICE_X97Y106_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X64Y106_SLICE_X97Y106_BO5),
.O6(CLBLM_L_X64Y106_SLICE_X97Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a000005aaaf0aa)
  ) CLBLM_L_X64Y106_SLICE_X97Y106_ALUT (
.I0(CLBLM_L_X64Y106_SLICE_X97Y106_B5Q),
.I1(1'b1),
.I2(CLBLM_L_X64Y106_SLICE_X97Y106_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X64Y106_SLICE_X97Y106_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X64Y106_SLICE_X97Y106_AO5),
.O6(CLBLM_L_X64Y106_SLICE_X97Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y122_SLICE_X96Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y121_SLICE_X102Y121_AQ),
.Q(CLBLM_L_X64Y122_SLICE_X96Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y122_SLICE_X96Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y122_SLICE_X96Y122_DO5),
.O6(CLBLM_L_X64Y122_SLICE_X96Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y122_SLICE_X96Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y122_SLICE_X96Y122_CO5),
.O6(CLBLM_L_X64Y122_SLICE_X96Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y122_SLICE_X96Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y122_SLICE_X96Y122_BO5),
.O6(CLBLM_L_X64Y122_SLICE_X96Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y122_SLICE_X96Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y122_SLICE_X96Y122_AO5),
.O6(CLBLM_L_X64Y122_SLICE_X96Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y122_SLICE_X97Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y122_SLICE_X97Y122_DO5),
.O6(CLBLM_L_X64Y122_SLICE_X97Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y122_SLICE_X97Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y122_SLICE_X97Y122_CO5),
.O6(CLBLM_L_X64Y122_SLICE_X97Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y122_SLICE_X97Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y122_SLICE_X97Y122_BO5),
.O6(CLBLM_L_X64Y122_SLICE_X97Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y122_SLICE_X97Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y122_SLICE_X97Y122_AO5),
.O6(CLBLM_L_X64Y122_SLICE_X97Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y95_SLICE_X102Y95_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y95_SLICE_X102Y95_AQ),
.Q(CLBLM_L_X68Y95_SLICE_X102Y95_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y95_SLICE_X102Y95_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y95_SLICE_X102Y95_AO6),
.Q(CLBLM_L_X68Y95_SLICE_X102Y95_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y95_SLICE_X102Y95_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y95_SLICE_X102Y95_DO5),
.O6(CLBLM_L_X68Y95_SLICE_X102Y95_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y95_SLICE_X102Y95_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y95_SLICE_X102Y95_CO5),
.O6(CLBLM_L_X68Y95_SLICE_X102Y95_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha000f00022003300)
  ) CLBLM_L_X68Y95_SLICE_X102Y95_BLUT (
.I0(CLBLM_L_X60Y94_SLICE_X90Y94_CQ),
.I1(CLBLM_L_X62Y95_SLICE_X92Y95_BQ),
.I2(CLBLM_L_X68Y95_SLICE_X102Y95_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X68Y99_SLICE_X102Y99_AQ),
.I5(CLBLM_L_X68Y95_SLICE_X102Y95_A5Q),
.O5(CLBLM_L_X68Y95_SLICE_X102Y95_BO5),
.O6(CLBLM_L_X68Y95_SLICE_X102Y95_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c005500cc005500)
  ) CLBLM_L_X68Y95_SLICE_X102Y95_ALUT (
.I0(CLBLM_L_X60Y94_SLICE_X90Y94_CQ),
.I1(CLBLM_L_X62Y95_SLICE_X92Y95_BQ),
.I2(CLBLM_L_X68Y95_SLICE_X102Y95_AQ),
.I3(CLBLM_L_X68Y95_SLICE_X102Y95_BO6),
.I4(CLBLM_L_X60Y94_SLICE_X90Y94_BQ),
.I5(CLBLM_L_X68Y95_SLICE_X102Y95_A5Q),
.O5(CLBLM_L_X68Y95_SLICE_X102Y95_AO5),
.O6(CLBLM_L_X68Y95_SLICE_X102Y95_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y95_SLICE_X103Y95_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y95_SLICE_X103Y95_DO5),
.O6(CLBLM_L_X68Y95_SLICE_X103Y95_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y95_SLICE_X103Y95_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y95_SLICE_X103Y95_CO5),
.O6(CLBLM_L_X68Y95_SLICE_X103Y95_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y95_SLICE_X103Y95_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y95_SLICE_X103Y95_BO5),
.O6(CLBLM_L_X68Y95_SLICE_X103Y95_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y95_SLICE_X103Y95_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y95_SLICE_X103Y95_AO5),
.O6(CLBLM_L_X68Y95_SLICE_X103Y95_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y96_SLICE_X102Y96_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y96_SLICE_X102Y96_AO6),
.Q(CLBLM_L_X68Y96_SLICE_X102Y96_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbbbbbb0000000)
  ) CLBLM_L_X68Y96_SLICE_X102Y96_DLUT (
.I0(CLBLM_L_X68Y96_SLICE_X102Y96_CO6),
.I1(CLBLM_L_X68Y96_SLICE_X103Y96_AO6),
.I2(CLBLM_L_X68Y96_SLICE_X102Y96_AQ),
.I3(CLBLM_L_X68Y99_SLICE_X102Y99_BO6),
.I4(CLBLM_L_X62Y95_SLICE_X92Y95_BQ),
.I5(CLBLM_L_X68Y96_SLICE_X102Y96_BO6),
.O5(CLBLM_L_X68Y96_SLICE_X102Y96_DO5),
.O6(CLBLM_L_X68Y96_SLICE_X102Y96_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000088880000f000)
  ) CLBLM_L_X68Y96_SLICE_X102Y96_CLUT (
.I0(CLBLM_L_X62Y95_SLICE_X92Y95_BQ),
.I1(CLBLM_R_X67Y97_SLICE_X100Y97_AQ),
.I2(CLBLM_R_X67Y98_SLICE_X101Y98_DQ),
.I3(CLBLM_L_X68Y95_SLICE_X102Y95_A5Q),
.I4(CLBLM_L_X68Y99_SLICE_X103Y99_CQ),
.I5(CLBLM_L_X68Y99_SLICE_X103Y99_C5Q),
.O5(CLBLM_L_X68Y96_SLICE_X102Y96_CO5),
.O6(CLBLM_L_X68Y96_SLICE_X102Y96_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h555d5555aaaeaaaa)
  ) CLBLM_L_X68Y96_SLICE_X102Y96_BLUT (
.I0(CLBLM_L_X68Y98_SLICE_X103Y98_A5Q),
.I1(CLBLM_L_X60Y94_SLICE_X90Y94_BQ),
.I2(CLBLM_L_X68Y99_SLICE_X103Y99_CQ),
.I3(CLBLM_L_X68Y99_SLICE_X103Y99_C5Q),
.I4(CLBLM_R_X67Y96_SLICE_X101Y96_CQ),
.I5(CLBLM_L_X68Y95_SLICE_X102Y95_AQ),
.O5(CLBLM_L_X68Y96_SLICE_X102Y96_BO5),
.O6(CLBLM_L_X68Y96_SLICE_X102Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3c0f3c0f3c0bb88)
  ) CLBLM_L_X68Y96_SLICE_X102Y96_ALUT (
.I0(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_L_X68Y96_SLICE_X102Y96_AQ),
.I3(CLBLM_L_X68Y98_SLICE_X102Y98_CQ),
.I4(CLBLM_R_X67Y98_SLICE_X101Y98_BO6),
.I5(CLBLM_R_X67Y98_SLICE_X100Y98_CO6),
.O5(CLBLM_L_X68Y96_SLICE_X102Y96_AO5),
.O6(CLBLM_L_X68Y96_SLICE_X102Y96_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y96_SLICE_X103Y96_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y96_SLICE_X103Y96_DO5),
.O6(CLBLM_L_X68Y96_SLICE_X103Y96_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y96_SLICE_X103Y96_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y96_SLICE_X103Y96_CO5),
.O6(CLBLM_L_X68Y96_SLICE_X103Y96_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800000088000000)
  ) CLBLM_L_X68Y96_SLICE_X103Y96_BLUT (
.I0(CLBLM_L_X68Y95_SLICE_X102Y95_A5Q),
.I1(CLBLM_L_X68Y95_SLICE_X102Y95_AQ),
.I2(1'b1),
.I3(CLBLM_L_X62Y95_SLICE_X92Y95_BQ),
.I4(CLBLM_L_X60Y94_SLICE_X90Y94_BQ),
.I5(1'b1),
.O5(CLBLM_L_X68Y96_SLICE_X103Y96_BO5),
.O6(CLBLM_L_X68Y96_SLICE_X103Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6666666606666666)
  ) CLBLM_L_X68Y96_SLICE_X103Y96_ALUT (
.I0(CLBLM_L_X68Y98_SLICE_X103Y98_A5Q),
.I1(CLBLM_L_X68Y95_SLICE_X102Y95_AQ),
.I2(CLBLM_L_X68Y98_SLICE_X102Y98_DQ),
.I3(CLBLM_L_X60Y94_SLICE_X90Y94_BQ),
.I4(CLBLM_L_X68Y99_SLICE_X103Y99_CQ),
.I5(CLBLM_L_X68Y99_SLICE_X103Y99_C5Q),
.O5(CLBLM_L_X68Y96_SLICE_X103Y96_AO5),
.O6(CLBLM_L_X68Y96_SLICE_X103Y96_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y97_SLICE_X102Y97_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y95_SLICE_X92Y95_CQ),
.Q(CLBLM_L_X68Y97_SLICE_X102Y97_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h153fff553f3fffff)
  ) CLBLM_L_X68Y97_SLICE_X102Y97_DLUT (
.I0(CLBLM_L_X68Y95_SLICE_X102Y95_A5Q),
.I1(CLBLM_L_X68Y98_SLICE_X103Y98_CQ),
.I2(CLBLM_L_X60Y97_SLICE_X90Y97_DQ),
.I3(CLBLM_L_X68Y95_SLICE_X102Y95_AQ),
.I4(CLBLM_L_X68Y98_SLICE_X103Y98_A5Q),
.I5(CLBLM_L_X68Y98_SLICE_X102Y98_CQ),
.O5(CLBLM_L_X68Y97_SLICE_X102Y97_DO5),
.O6(CLBLM_L_X68Y97_SLICE_X102Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaa2a2aaa2)
  ) CLBLM_L_X68Y97_SLICE_X102Y97_CLUT (
.I0(CLBLM_L_X70Y106_SLICE_X104Y106_CO6),
.I1(CLBLM_L_X68Y97_SLICE_X103Y97_CO6),
.I2(CLBLM_L_X68Y99_SLICE_X102Y99_CO6),
.I3(CLBLM_L_X68Y97_SLICE_X102Y97_AO5),
.I4(CLBLM_L_X68Y97_SLICE_X102Y97_DO6),
.I5(CLBLM_L_X68Y96_SLICE_X102Y96_DO6),
.O5(CLBLM_L_X68Y97_SLICE_X102Y97_CO5),
.O6(CLBLM_L_X68Y97_SLICE_X102Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h15ffffff3fffffff)
  ) CLBLM_L_X68Y97_SLICE_X102Y97_BLUT (
.I0(CLBLM_R_X67Y97_SLICE_X101Y97_CQ),
.I1(CLBLM_L_X68Y95_SLICE_X102Y95_AQ),
.I2(CLBLM_R_X67Y97_SLICE_X101Y97_BQ),
.I3(CLBLM_L_X68Y99_SLICE_X103Y99_C5Q),
.I4(CLBLM_L_X68Y99_SLICE_X103Y99_CQ),
.I5(CLBLM_L_X68Y97_SLICE_X103Y97_AQ),
.O5(CLBLM_L_X68Y97_SLICE_X102Y97_BO5),
.O6(CLBLM_L_X68Y97_SLICE_X102Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaeaa0f0f0000)
  ) CLBLM_L_X68Y97_SLICE_X102Y97_ALUT (
.I0(CLBLM_L_X68Y98_SLICE_X103Y98_A5Q),
.I1(CLBLM_L_X60Y97_SLICE_X90Y97_DQ),
.I2(CLBLM_L_X68Y99_SLICE_X103Y99_C5Q),
.I3(CLBLM_R_X67Y97_SLICE_X101Y97_DQ),
.I4(CLBLM_L_X68Y99_SLICE_X103Y99_CQ),
.I5(1'b1),
.O5(CLBLM_L_X68Y97_SLICE_X102Y97_AO5),
.O6(CLBLM_L_X68Y97_SLICE_X102Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y97_SLICE_X103Y97_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y99_SLICE_X102Y99_AQ),
.Q(CLBLM_L_X68Y97_SLICE_X103Y97_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8f0f8f0f0f0f0f0f)
  ) CLBLM_L_X68Y97_SLICE_X103Y97_DLUT (
.I0(CLBLM_L_X68Y99_SLICE_X103Y99_C5Q),
.I1(CLBLM_L_X62Y95_SLICE_X92Y95_CQ),
.I2(CLBLM_L_X68Y98_SLICE_X103Y98_A5Q),
.I3(CLBLM_L_X68Y99_SLICE_X103Y99_CQ),
.I4(1'b1),
.I5(CLBLM_L_X68Y99_SLICE_X103Y99_BQ),
.O5(CLBLM_L_X68Y97_SLICE_X103Y97_DO5),
.O6(CLBLM_L_X68Y97_SLICE_X103Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000cccc0050ccdc)
  ) CLBLM_L_X68Y97_SLICE_X103Y97_CLUT (
.I0(CLBLM_L_X68Y97_SLICE_X103Y97_AO6),
.I1(CLBLM_L_X68Y98_SLICE_X103Y98_DO6),
.I2(CLBLM_L_X68Y97_SLICE_X102Y97_BO6),
.I3(CLBLM_L_X68Y97_SLICE_X102Y97_AO6),
.I4(CLBLM_L_X68Y97_SLICE_X103Y97_DO6),
.I5(CLBLM_L_X68Y97_SLICE_X103Y97_BO6),
.O5(CLBLM_L_X68Y97_SLICE_X103Y97_CO5),
.O6(CLBLM_L_X68Y97_SLICE_X103Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a080a0008080000)
  ) CLBLM_L_X68Y97_SLICE_X103Y97_BLUT (
.I0(CLBLM_L_X68Y99_SLICE_X103Y99_CQ),
.I1(CLBLM_R_X67Y96_SLICE_X101Y96_BQ),
.I2(CLBLM_L_X68Y99_SLICE_X103Y99_C5Q),
.I3(CLBLM_L_X68Y99_SLICE_X102Y99_AQ),
.I4(CLBLM_L_X68Y97_SLICE_X102Y97_AQ),
.I5(CLBLM_R_X67Y97_SLICE_X101Y97_AQ),
.O5(CLBLM_L_X68Y97_SLICE_X103Y97_BO5),
.O6(CLBLM_L_X68Y97_SLICE_X103Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f00080008000800)
  ) CLBLM_L_X68Y97_SLICE_X103Y97_ALUT (
.I0(CLBLM_R_X67Y96_SLICE_X101Y96_DQ),
.I1(CLBLM_L_X62Y95_SLICE_X92Y95_CQ),
.I2(CLBLM_L_X68Y99_SLICE_X103Y99_CQ),
.I3(CLBLM_L_X68Y99_SLICE_X103Y99_C5Q),
.I4(CLBLM_R_X67Y96_SLICE_X101Y96_AQ),
.I5(CLBLM_L_X60Y94_SLICE_X90Y94_CQ),
.O5(CLBLM_L_X68Y97_SLICE_X103Y97_AO5),
.O6(CLBLM_L_X68Y97_SLICE_X103Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y98_SLICE_X102Y98_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y98_SLICE_X102Y98_AO6),
.Q(CLBLM_L_X68Y98_SLICE_X102Y98_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y98_SLICE_X102Y98_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y98_SLICE_X102Y98_BO6),
.Q(CLBLM_L_X68Y98_SLICE_X102Y98_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y98_SLICE_X102Y98_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y98_SLICE_X102Y98_CO6),
.Q(CLBLM_L_X68Y98_SLICE_X102Y98_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y98_SLICE_X102Y98_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y98_SLICE_X102Y98_DO6),
.Q(CLBLM_L_X68Y98_SLICE_X102Y98_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f3c0aaaaaaaa)
  ) CLBLM_L_X68Y98_SLICE_X102Y98_DLUT (
.I0(CLBLM_R_X67Y97_SLICE_X100Y97_AQ),
.I1(CLBLM_R_X67Y98_SLICE_X101Y98_CO5),
.I2(CLBLM_L_X68Y98_SLICE_X102Y98_DQ),
.I3(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I4(CLBLM_R_X67Y98_SLICE_X100Y98_CO5),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X68Y98_SLICE_X102Y98_DO5),
.O6(CLBLM_L_X68Y98_SLICE_X102Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccaaf0f0f0f0)
  ) CLBLM_L_X68Y98_SLICE_X102Y98_CLUT (
.I0(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I1(CLBLM_L_X68Y98_SLICE_X102Y98_CQ),
.I2(CLBLM_L_X68Y98_SLICE_X102Y98_BQ),
.I3(CLBLM_R_X67Y98_SLICE_X101Y98_BO6),
.I4(CLBLM_R_X67Y98_SLICE_X101Y98_AO5),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X68Y98_SLICE_X102Y98_CO5),
.O6(CLBLM_L_X68Y98_SLICE_X102Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccf0ccf0aaf0)
  ) CLBLM_L_X68Y98_SLICE_X102Y98_BLUT (
.I0(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I1(CLBLM_L_X68Y98_SLICE_X102Y98_BQ),
.I2(CLBLM_L_X68Y99_SLICE_X103Y99_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_R_X67Y98_SLICE_X101Y98_BO6),
.I5(CLBLM_R_X67Y98_SLICE_X101Y98_AO6),
.O5(CLBLM_L_X68Y98_SLICE_X102Y98_BO5),
.O6(CLBLM_L_X68Y98_SLICE_X102Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3c0f3c0f3c4f380)
  ) CLBLM_L_X68Y98_SLICE_X102Y98_ALUT (
.I0(CLBLM_R_X67Y98_SLICE_X100Y98_A5Q),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_L_X68Y98_SLICE_X102Y98_AQ),
.I3(CLBLM_L_X68Y101_SLICE_X102Y101_BQ),
.I4(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I5(CLBLM_R_X67Y98_SLICE_X101Y98_AO6),
.O5(CLBLM_L_X68Y98_SLICE_X102Y98_AO5),
.O6(CLBLM_L_X68Y98_SLICE_X102Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y98_SLICE_X103Y98_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y98_SLICE_X103Y98_AO5),
.Q(CLBLM_L_X68Y98_SLICE_X103Y98_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y98_SLICE_X103Y98_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y98_SLICE_X103Y98_AO6),
.Q(CLBLM_L_X68Y98_SLICE_X103Y98_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y98_SLICE_X103Y98_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y98_SLICE_X103Y98_BO6),
.Q(CLBLM_L_X68Y98_SLICE_X103Y98_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y98_SLICE_X103Y98_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y98_SLICE_X103Y98_CO6),
.Q(CLBLM_L_X68Y98_SLICE_X103Y98_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1fdf3fffdfdffff)
  ) CLBLM_L_X68Y98_SLICE_X103Y98_DLUT (
.I0(CLBLM_L_X68Y98_SLICE_X102Y98_AQ),
.I1(CLBLM_L_X68Y99_SLICE_X103Y99_C5Q),
.I2(CLBLM_L_X68Y99_SLICE_X103Y99_CQ),
.I3(CLBLM_L_X68Y98_SLICE_X103Y98_BQ),
.I4(CLBLM_L_X68Y99_SLICE_X102Y99_AQ),
.I5(CLBLM_L_X68Y97_SLICE_X103Y97_AQ),
.O5(CLBLM_L_X68Y98_SLICE_X103Y98_DO5),
.O6(CLBLM_L_X68Y98_SLICE_X103Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccddcc88f0f0f0f0)
  ) CLBLM_L_X68Y98_SLICE_X103Y98_CLUT (
.I0(CLBLM_R_X67Y98_SLICE_X100Y98_CO6),
.I1(CLBLM_L_X68Y98_SLICE_X103Y98_CQ),
.I2(CLBLM_L_X68Y98_SLICE_X103Y98_BQ),
.I3(CLBLM_R_X67Y98_SLICE_X101Y98_BO5),
.I4(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X68Y98_SLICE_X103Y98_CO5),
.O6(CLBLM_L_X68Y98_SLICE_X103Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00d8ffd800)
  ) CLBLM_L_X68Y98_SLICE_X103Y98_BLUT (
.I0(CLBLM_R_X67Y98_SLICE_X101Y98_AO5),
.I1(CLBLM_L_X68Y98_SLICE_X103Y98_BQ),
.I2(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X68Y98_SLICE_X102Y98_AQ),
.I5(CLBLM_R_X67Y98_SLICE_X101Y98_BO5),
.O5(CLBLM_L_X68Y98_SLICE_X103Y98_BO5),
.O6(CLBLM_L_X68Y98_SLICE_X103Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa0066f066f0)
  ) CLBLM_L_X68Y98_SLICE_X103Y98_ALUT (
.I0(CLBLM_L_X68Y98_SLICE_X103Y98_A5Q),
.I1(CLBLM_L_X68Y96_SLICE_X103Y96_BO6),
.I2(CLBLM_L_X68Y97_SLICE_X102Y97_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X72Y98_SLICE_X108Y98_BQ),
.I5(1'b1),
.O5(CLBLM_L_X68Y98_SLICE_X103Y98_AO5),
.O6(CLBLM_L_X68Y98_SLICE_X103Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y99_SLICE_X102Y99_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X60Y94_SLICE_X90Y94_CQ),
.Q(CLBLM_L_X68Y99_SLICE_X102Y99_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000800000000000)
  ) CLBLM_L_X68Y99_SLICE_X102Y99_DLUT (
.I0(CLBLM_L_X68Y98_SLICE_X103Y98_A5Q),
.I1(CLBLM_L_X68Y101_SLICE_X102Y101_CQ),
.I2(CLBLM_L_X68Y99_SLICE_X103Y99_C5Q),
.I3(CLBLM_L_X68Y99_SLICE_X103Y99_CQ),
.I4(1'b1),
.I5(CLBLM_L_X60Y94_SLICE_X90Y94_CQ),
.O5(CLBLM_L_X68Y99_SLICE_X102Y99_DO5),
.O6(CLBLM_L_X68Y99_SLICE_X102Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffff8000)
  ) CLBLM_L_X68Y99_SLICE_X102Y99_CLUT (
.I0(CLBLM_L_X68Y99_SLICE_X102Y99_AO6),
.I1(CLBLM_L_X68Y99_SLICE_X103Y99_AQ),
.I2(CLBLM_L_X68Y97_SLICE_X102Y97_AQ),
.I3(CLBLM_L_X68Y98_SLICE_X103Y98_A5Q),
.I4(CLBLM_L_X68Y99_SLICE_X102Y99_BO5),
.I5(CLBLM_L_X68Y99_SLICE_X102Y99_DO6),
.O5(CLBLM_L_X68Y99_SLICE_X102Y99_CO5),
.O6(CLBLM_L_X68Y99_SLICE_X102Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0000000008000)
  ) CLBLM_L_X68Y99_SLICE_X102Y99_BLUT (
.I0(CLBLM_L_X68Y95_SLICE_X102Y95_AQ),
.I1(CLBLM_L_X68Y98_SLICE_X103Y98_A5Q),
.I2(CLBLM_L_X68Y99_SLICE_X103Y99_C5Q),
.I3(CLBLM_L_X68Y98_SLICE_X102Y98_BQ),
.I4(CLBLM_L_X68Y99_SLICE_X103Y99_CQ),
.I5(1'b1),
.O5(CLBLM_L_X68Y99_SLICE_X102Y99_BO5),
.O6(CLBLM_L_X68Y99_SLICE_X102Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000f0f80000000)
  ) CLBLM_L_X68Y99_SLICE_X102Y99_ALUT (
.I0(CLBLM_L_X70Y106_SLICE_X104Y106_CO6),
.I1(CLBLM_L_X68Y98_SLICE_X103Y98_A5Q),
.I2(CLBLM_L_X68Y99_SLICE_X103Y99_C5Q),
.I3(CLBLM_L_X60Y94_SLICE_X90Y94_CQ),
.I4(CLBLM_L_X68Y99_SLICE_X103Y99_CQ),
.I5(1'b1),
.O5(CLBLM_L_X68Y99_SLICE_X102Y99_AO5),
.O6(CLBLM_L_X68Y99_SLICE_X102Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y99_SLICE_X103Y99_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y99_SLICE_X103Y99_CO5),
.Q(CLBLM_L_X68Y99_SLICE_X103Y99_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y99_SLICE_X103Y99_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y99_SLICE_X103Y99_DO5),
.Q(CLBLM_L_X68Y99_SLICE_X103Y99_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y99_SLICE_X103Y99_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y99_SLICE_X103Y99_AO6),
.Q(CLBLM_L_X68Y99_SLICE_X103Y99_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y99_SLICE_X103Y99_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y99_SLICE_X103Y99_BO6),
.Q(CLBLM_L_X68Y99_SLICE_X103Y99_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y99_SLICE_X103Y99_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y99_SLICE_X103Y99_CO6),
.Q(CLBLM_L_X68Y99_SLICE_X103Y99_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y99_SLICE_X103Y99_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y99_SLICE_X103Y99_DO6),
.Q(CLBLM_L_X68Y99_SLICE_X103Y99_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa77aa70f070f0)
  ) CLBLM_L_X68Y99_SLICE_X103Y99_DLUT (
.I0(CLBLM_L_X68Y98_SLICE_X103Y98_A5Q),
.I1(CLBLM_L_X68Y96_SLICE_X103Y96_BO6),
.I2(CLBLM_L_X68Y99_SLICE_X103Y99_DQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X68Y99_SLICE_X103Y99_D5Q),
.I5(1'b1),
.O5(CLBLM_L_X68Y99_SLICE_X103Y99_DO5),
.O6(CLBLM_L_X68Y99_SLICE_X103Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6caa6caa5aff5a00)
  ) CLBLM_L_X68Y99_SLICE_X103Y99_CLUT (
.I0(CLBLM_L_X68Y99_SLICE_X103Y99_C5Q),
.I1(CLBLM_L_X68Y99_SLICE_X103Y99_CQ),
.I2(CLBLM_L_X70Y106_SLICE_X104Y106_CO6),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X68Y99_SLICE_X103Y99_D5Q),
.I5(1'b1),
.O5(CLBLM_L_X68Y99_SLICE_X103Y99_CO5),
.O6(CLBLM_L_X68Y99_SLICE_X103Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccfc0aaaaaaaa)
  ) CLBLM_L_X68Y99_SLICE_X103Y99_BLUT (
.I0(CLBLM_L_X68Y98_SLICE_X103Y98_CQ),
.I1(CLBLM_L_X68Y99_SLICE_X103Y99_BQ),
.I2(CLBLM_R_X67Y98_SLICE_X100Y98_CO5),
.I3(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I4(CLBLM_R_X67Y98_SLICE_X101Y98_BO5),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X68Y99_SLICE_X103Y99_BO5),
.O6(CLBLM_L_X68Y99_SLICE_X103Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0faf050cccccccc)
  ) CLBLM_L_X68Y99_SLICE_X103Y99_ALUT (
.I0(CLBLM_R_X67Y98_SLICE_X100Y98_B5Q),
.I1(CLBLM_L_X68Y99_SLICE_X103Y99_BQ),
.I2(CLBLM_L_X68Y99_SLICE_X103Y99_AQ),
.I3(CLBLM_R_X67Y98_SLICE_X101Y98_BO5),
.I4(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X68Y99_SLICE_X103Y99_AO5),
.O6(CLBLM_L_X68Y99_SLICE_X103Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y100_SLICE_X102Y100_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y100_SLICE_X102Y100_DO5),
.O6(CLBLM_L_X68Y100_SLICE_X102Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y100_SLICE_X102Y100_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y100_SLICE_X102Y100_CO5),
.O6(CLBLM_L_X68Y100_SLICE_X102Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y100_SLICE_X102Y100_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y100_SLICE_X102Y100_BO5),
.O6(CLBLM_L_X68Y100_SLICE_X102Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y100_SLICE_X102Y100_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y100_SLICE_X102Y100_AO5),
.O6(CLBLM_L_X68Y100_SLICE_X102Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y100_SLICE_X103Y100_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y100_SLICE_X103Y100_DO5),
.O6(CLBLM_L_X68Y100_SLICE_X103Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y100_SLICE_X103Y100_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y100_SLICE_X103Y100_CO5),
.O6(CLBLM_L_X68Y100_SLICE_X103Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y100_SLICE_X103Y100_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y100_SLICE_X103Y100_BO5),
.O6(CLBLM_L_X68Y100_SLICE_X103Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heaeeeaaaaeaaaeee)
  ) CLBLM_L_X68Y100_SLICE_X103Y100_ALUT (
.I0(CLBLM_L_X68Y105_SLICE_X103Y105_BQ),
.I1(CLBLM_L_X70Y106_SLICE_X104Y106_CO6),
.I2(CLBLM_L_X68Y99_SLICE_X103Y99_D5Q),
.I3(CLBLM_L_X68Y99_SLICE_X103Y99_C5Q),
.I4(CLBLM_L_X68Y99_SLICE_X103Y99_DQ),
.I5(CLBLM_L_X68Y99_SLICE_X103Y99_CQ),
.O5(CLBLM_L_X68Y100_SLICE_X103Y100_AO5),
.O6(CLBLM_L_X68Y100_SLICE_X103Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y101_SLICE_X102Y101_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y105_SLICE_X102Y105_AQ),
.Q(CLBLM_L_X68Y101_SLICE_X102Y101_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y101_SLICE_X102Y101_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y101_SLICE_X102Y101_AO6),
.Q(CLBLM_L_X68Y101_SLICE_X102Y101_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y101_SLICE_X102Y101_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y101_SLICE_X102Y101_BO6),
.Q(CLBLM_L_X68Y101_SLICE_X102Y101_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y101_SLICE_X102Y101_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y101_SLICE_X102Y101_CO6),
.Q(CLBLM_L_X68Y101_SLICE_X102Y101_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y101_SLICE_X102Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y101_SLICE_X102Y101_DO5),
.O6(CLBLM_L_X68Y101_SLICE_X102Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fcfcff000c0c0)
  ) CLBLM_L_X68Y101_SLICE_X102Y101_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X68Y101_SLICE_X102Y101_CQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I4(CLBLM_L_X68Y101_SLICE_X102Y101_BO5),
.I5(CLBLM_L_X68Y98_SLICE_X102Y98_DQ),
.O5(CLBLM_L_X68Y101_SLICE_X102Y101_CO5),
.O6(CLBLM_L_X68Y101_SLICE_X102Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6fc06fc088008800)
  ) CLBLM_L_X68Y101_SLICE_X102Y101_BLUT (
.I0(CLBLM_R_X67Y98_SLICE_X100Y98_B5Q),
.I1(CLBLM_L_X68Y101_SLICE_X102Y101_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_R_X67Y98_SLICE_X100Y98_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y101_SLICE_X102Y101_BO5),
.O6(CLBLM_L_X68Y101_SLICE_X102Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00fff0ff0000fc00)
  ) CLBLM_L_X68Y101_SLICE_X102Y101_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X68Y105_SLICE_X102Y105_AQ),
.I2(CLBLM_L_X68Y101_SLICE_X102Y101_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X64Y101_SLICE_X96Y101_AQ),
.I5(CLBLM_L_X68Y101_SLICE_X102Y101_A5Q),
.O5(CLBLM_L_X68Y101_SLICE_X102Y101_AO5),
.O6(CLBLM_L_X68Y101_SLICE_X102Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y101_SLICE_X103Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y101_SLICE_X103Y101_DO5),
.O6(CLBLM_L_X68Y101_SLICE_X103Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y101_SLICE_X103Y101_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y101_SLICE_X103Y101_CO5),
.O6(CLBLM_L_X68Y101_SLICE_X103Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y101_SLICE_X103Y101_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y101_SLICE_X103Y101_BO5),
.O6(CLBLM_L_X68Y101_SLICE_X103Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y101_SLICE_X103Y101_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y101_SLICE_X103Y101_AO5),
.O6(CLBLM_L_X68Y101_SLICE_X103Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y102_SLICE_X102Y102_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y102_SLICE_X102Y102_AO6),
.Q(CLBLM_L_X68Y102_SLICE_X102Y102_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y102_SLICE_X102Y102_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y102_SLICE_X102Y102_BO6),
.Q(CLBLM_L_X68Y102_SLICE_X102Y102_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y102_SLICE_X102Y102_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y102_SLICE_X102Y102_CO6),
.Q(CLBLM_L_X68Y102_SLICE_X102Y102_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y102_SLICE_X102Y102_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y102_SLICE_X102Y102_DO6),
.Q(CLBLM_L_X68Y102_SLICE_X102Y102_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h708ff00f00000000)
  ) CLBLM_L_X68Y102_SLICE_X102Y102_DLUT (
.I0(CLBLM_L_X68Y101_SLICE_X102Y101_BQ),
.I1(CLBLM_R_X67Y98_SLICE_X100Y98_A5Q),
.I2(CLBLM_L_X68Y102_SLICE_X102Y102_DQ),
.I3(CLBLL_R_X79Y99_SLICE_X122Y99_AO6),
.I4(CLBLM_R_X67Y98_SLICE_X100Y98_B5Q),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X68Y102_SLICE_X102Y102_DO5),
.O6(CLBLM_L_X68Y102_SLICE_X102Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5acc5accf0f0f0f0)
  ) CLBLM_L_X68Y102_SLICE_X102Y102_CLUT (
.I0(CLBLM_L_X68Y102_SLICE_X102Y102_BQ),
.I1(CLBLM_L_X68Y102_SLICE_X102Y102_CQ),
.I2(CLBLM_L_X68Y102_SLICE_X102Y102_AQ),
.I3(CLBLM_L_X68Y99_SLICE_X102Y99_AO5),
.I4(1'b1),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X68Y102_SLICE_X102Y102_CO5),
.O6(CLBLM_L_X68Y102_SLICE_X102Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he4ccccccf0f0f0f0)
  ) CLBLM_L_X68Y102_SLICE_X102Y102_BLUT (
.I0(CLBLM_R_X67Y98_SLICE_X100Y98_B5Q),
.I1(CLBLM_L_X68Y102_SLICE_X102Y102_BQ),
.I2(CLBLM_L_X68Y102_SLICE_X102Y102_DQ),
.I3(CLBLM_R_X67Y98_SLICE_X100Y98_A5Q),
.I4(CLBLM_L_X68Y101_SLICE_X102Y101_BQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X68Y102_SLICE_X102Y102_BO5),
.O6(CLBLM_L_X68Y102_SLICE_X102Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc003cff3c00)
  ) CLBLM_L_X68Y102_SLICE_X102Y102_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X68Y97_SLICE_X102Y97_CO6),
.I2(CLBLM_L_X68Y102_SLICE_X102Y102_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X68Y102_SLICE_X102Y102_BQ),
.I5(CLBLM_L_X68Y99_SLICE_X102Y99_AO5),
.O5(CLBLM_L_X68Y102_SLICE_X102Y102_AO5),
.O6(CLBLM_L_X68Y102_SLICE_X102Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y102_SLICE_X103Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y102_SLICE_X103Y102_DO5),
.O6(CLBLM_L_X68Y102_SLICE_X103Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y102_SLICE_X103Y102_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y102_SLICE_X103Y102_CO5),
.O6(CLBLM_L_X68Y102_SLICE_X103Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y102_SLICE_X103Y102_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y102_SLICE_X103Y102_BO5),
.O6(CLBLM_L_X68Y102_SLICE_X103Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y102_SLICE_X103Y102_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y102_SLICE_X103Y102_AO5),
.O6(CLBLM_L_X68Y102_SLICE_X103Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y103_SLICE_X102Y103_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y103_SLICE_X102Y103_BO5),
.Q(CLBLM_L_X68Y103_SLICE_X102Y103_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y103_SLICE_X102Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y103_SLICE_X102Y103_AO6),
.Q(CLBLM_L_X68Y103_SLICE_X102Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y103_SLICE_X102Y103_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y103_SLICE_X102Y103_BO6),
.Q(CLBLM_L_X68Y103_SLICE_X102Y103_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y103_SLICE_X102Y103_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y103_SLICE_X102Y103_CO6),
.Q(CLBLM_L_X68Y103_SLICE_X102Y103_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y103_SLICE_X102Y103_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y103_SLICE_X102Y103_DO6),
.Q(CLBLM_L_X68Y103_SLICE_X102Y103_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacccacc3acc3acc)
  ) CLBLM_L_X68Y103_SLICE_X102Y103_DLUT (
.I0(CLBLM_L_X68Y103_SLICE_X102Y103_DQ),
.I1(CLBLM_L_X68Y103_SLICE_X102Y103_CQ),
.I2(CLBLM_L_X68Y101_SLICE_X102Y101_BO5),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(1'b1),
.I5(CLBLM_R_X67Y103_SLICE_X100Y103_B5Q),
.O5(CLBLM_L_X68Y103_SLICE_X102Y103_DO5),
.O6(CLBLM_L_X68Y103_SLICE_X102Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hec4cff00ccccff00)
  ) CLBLM_L_X68Y103_SLICE_X102Y103_CLUT (
.I0(CLBLM_L_X68Y101_SLICE_X102Y101_BQ),
.I1(CLBLM_L_X68Y103_SLICE_X102Y103_CQ),
.I2(CLBLM_R_X67Y98_SLICE_X100Y98_B5Q),
.I3(CLBLM_R_X67Y103_SLICE_X100Y103_B5Q),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_R_X67Y98_SLICE_X100Y98_A5Q),
.O5(CLBLM_L_X68Y103_SLICE_X102Y103_CO5),
.O6(CLBLM_L_X68Y103_SLICE_X102Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cff00ca3acccc)
  ) CLBLM_L_X68Y103_SLICE_X102Y103_BLUT (
.I0(CLBLM_L_X68Y103_SLICE_X102Y103_B5Q),
.I1(CLBLM_L_X68Y103_SLICE_X102Y103_BQ),
.I2(CLBLM_L_X68Y99_SLICE_X102Y99_AO5),
.I3(CLBLM_R_X67Y103_SLICE_X101Y103_AQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLM_L_X68Y103_SLICE_X102Y103_BO5),
.O6(CLBLM_L_X68Y103_SLICE_X102Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff33f3cccc00c0)
  ) CLBLM_L_X68Y103_SLICE_X102Y103_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_L_X68Y103_SLICE_X102Y103_AQ),
.I3(CLBLM_L_X70Y106_SLICE_X104Y106_CO6),
.I4(CLBLM_L_X68Y97_SLICE_X102Y97_CO6),
.I5(CLBLM_L_X68Y101_SLICE_X102Y101_CQ),
.O5(CLBLM_L_X68Y103_SLICE_X102Y103_AO5),
.O6(CLBLM_L_X68Y103_SLICE_X102Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y103_SLICE_X103Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y103_SLICE_X103Y103_DO5),
.O6(CLBLM_L_X68Y103_SLICE_X103Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y103_SLICE_X103Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y103_SLICE_X103Y103_CO5),
.O6(CLBLM_L_X68Y103_SLICE_X103Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y103_SLICE_X103Y103_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y103_SLICE_X103Y103_BO5),
.O6(CLBLM_L_X68Y103_SLICE_X103Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y103_SLICE_X103Y103_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y103_SLICE_X103Y103_AO5),
.O6(CLBLM_L_X68Y103_SLICE_X103Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y105_SLICE_X102Y105_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y106_SLICE_X102Y106_AO5),
.Q(CLBLM_L_X68Y105_SLICE_X102Y105_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y105_SLICE_X102Y105_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y105_SLICE_X102Y105_BO6),
.Q(CLBLM_L_X68Y105_SLICE_X102Y105_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y105_SLICE_X102Y105_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y105_SLICE_X102Y105_CO6),
.Q(CLBLM_L_X68Y105_SLICE_X102Y105_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffbbffb3)
  ) CLBLM_L_X68Y105_SLICE_X102Y105_DLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_R_X67Y105_SLICE_X101Y105_CO6),
.I2(CLBLM_R_X65Y105_SLICE_X98Y105_CQ),
.I3(CLBLM_L_X68Y105_SLICE_X102Y105_AO5),
.I4(CLBLM_R_X65Y106_SLICE_X99Y106_C5Q),
.I5(CLBLM_R_X65Y105_SLICE_X99Y105_BO5),
.O5(CLBLM_L_X68Y105_SLICE_X102Y105_DO5),
.O6(CLBLM_L_X68Y105_SLICE_X102Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff7f0080ff0000)
  ) CLBLM_L_X68Y105_SLICE_X102Y105_CLUT (
.I0(CLBLM_L_X68Y108_SLICE_X103Y108_AQ),
.I1(CLBLM_L_X68Y108_SLICE_X103Y108_A5Q),
.I2(CLBLM_L_X70Y106_SLICE_X104Y106_BQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X68Y105_SLICE_X102Y105_BQ),
.I5(CLBLM_L_X68Y105_SLICE_X102Y105_CQ),
.O5(CLBLM_L_X68Y105_SLICE_X102Y105_CO5),
.O6(CLBLM_L_X68Y105_SLICE_X102Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h46ccccccaaaaaaaa)
  ) CLBLM_L_X68Y105_SLICE_X102Y105_BLUT (
.I0(CLBLM_L_X68Y108_SLICE_X103Y108_A5Q),
.I1(CLBLM_L_X68Y105_SLICE_X102Y105_BQ),
.I2(CLBLM_L_X68Y105_SLICE_X102Y105_CQ),
.I3(CLBLM_L_X70Y106_SLICE_X104Y106_BQ),
.I4(CLBLM_L_X68Y108_SLICE_X103Y108_AQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X68Y105_SLICE_X102Y105_BO5),
.O6(CLBLM_L_X68Y105_SLICE_X102Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccc8ccc0ccc0)
  ) CLBLM_L_X68Y105_SLICE_X102Y105_ALUT (
.I0(CLBLM_R_X65Y105_SLICE_X98Y105_CQ),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_L_X70Y104_SLICE_X104Y104_BQ),
.I3(CLBLM_L_X70Y104_SLICE_X105Y104_D5Q),
.I4(CLBLM_R_X65Y106_SLICE_X99Y106_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X68Y105_SLICE_X102Y105_AO5),
.O6(CLBLM_L_X68Y105_SLICE_X102Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y105_SLICE_X103Y105_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y105_SLICE_X103Y105_AO6),
.Q(CLBLM_L_X68Y105_SLICE_X103Y105_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y105_SLICE_X103Y105_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y105_SLICE_X103Y105_BO6),
.Q(CLBLM_L_X68Y105_SLICE_X103Y105_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y105_SLICE_X103Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y105_SLICE_X103Y105_DO5),
.O6(CLBLM_L_X68Y105_SLICE_X103Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y105_SLICE_X103Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y105_SLICE_X103Y105_CO5),
.O6(CLBLM_L_X68Y105_SLICE_X103Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb000300030003000)
  ) CLBLM_L_X68Y105_SLICE_X103Y105_BLUT (
.I0(CLBLM_L_X68Y109_SLICE_X103Y109_BQ),
.I1(CLBLM_L_X70Y106_SLICE_X104Y106_CO6),
.I2(CLBLM_L_X68Y100_SLICE_X103Y100_AO6),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X68Y109_SLICE_X103Y109_B5Q),
.I5(CLBLM_L_X68Y108_SLICE_X103Y108_CO6),
.O5(CLBLM_L_X68Y105_SLICE_X103Y105_BO5),
.O6(CLBLM_L_X68Y105_SLICE_X103Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8ccf0ccf0ccf0cc)
  ) CLBLM_L_X68Y105_SLICE_X103Y105_ALUT (
.I0(CLBLM_L_X68Y109_SLICE_X103Y109_BQ),
.I1(CLBLM_L_X68Y105_SLICE_X103Y105_BQ),
.I2(CLBLM_L_X68Y105_SLICE_X103Y105_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X68Y109_SLICE_X103Y109_B5Q),
.I5(CLBLM_L_X68Y108_SLICE_X103Y108_CO6),
.O5(CLBLM_L_X68Y105_SLICE_X103Y105_AO5),
.O6(CLBLM_L_X68Y105_SLICE_X103Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffefffffffff)
  ) CLBLM_L_X68Y106_SLICE_X102Y106_DLUT (
.I0(CLBLM_L_X64Y104_SLICE_X96Y104_CQ),
.I1(CLBLM_R_X67Y109_SLICE_X100Y109_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X68Y102_SLICE_X102Y102_CQ),
.I4(CLBLM_L_X70Y104_SLICE_X105Y104_BQ),
.I5(CLBLM_R_X65Y100_SLICE_X98Y100_AQ),
.O5(CLBLM_L_X68Y106_SLICE_X102Y106_DO5),
.O6(CLBLM_L_X68Y106_SLICE_X102Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffef0f0f0f0)
  ) CLBLM_L_X68Y106_SLICE_X102Y106_CLUT (
.I0(CLBLM_R_X65Y100_SLICE_X98Y100_AQ),
.I1(CLBLL_R_X71Y108_SLICE_X106Y108_BQ),
.I2(CLBLM_L_X72Y105_SLICE_X108Y105_CQ),
.I3(CLBLM_R_X67Y109_SLICE_X100Y109_BQ),
.I4(CLBLM_L_X70Y104_SLICE_X105Y104_BQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X68Y106_SLICE_X102Y106_CO5),
.O6(CLBLM_L_X68Y106_SLICE_X102Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f5f5c4f531f5)
  ) CLBLM_L_X68Y106_SLICE_X102Y106_BLUT (
.I0(CLBLM_L_X68Y107_SLICE_X102Y107_AO5),
.I1(CLBLM_L_X64Y104_SLICE_X96Y104_CQ),
.I2(CLBLM_L_X68Y106_SLICE_X102Y106_DO6),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X68Y102_SLICE_X102Y102_CQ),
.I5(CLBLM_L_X68Y106_SLICE_X102Y106_CO6),
.O5(CLBLM_L_X68Y106_SLICE_X102Y106_BO5),
.O6(CLBLM_L_X68Y106_SLICE_X102Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaa8aaa8aaaa0000)
  ) CLBLM_L_X68Y106_SLICE_X102Y106_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X64Y104_SLICE_X96Y104_CQ),
.I2(CLBLM_L_X70Y104_SLICE_X105Y104_BQ),
.I3(CLBLM_R_X65Y100_SLICE_X98Y100_AQ),
.I4(CLBLM_L_X64Y105_SLICE_X96Y105_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X68Y106_SLICE_X102Y106_AO5),
.O6(CLBLM_L_X68Y106_SLICE_X102Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y106_SLICE_X103Y106_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y106_SLICE_X103Y106_BO5),
.Q(CLBLM_L_X68Y106_SLICE_X103Y106_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y106_SLICE_X103Y106_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y106_SLICE_X103Y106_BO6),
.Q(CLBLM_L_X68Y106_SLICE_X103Y106_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y106_SLICE_X103Y106_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y106_SLICE_X103Y106_CO6),
.Q(CLBLM_L_X68Y106_SLICE_X103Y106_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000200000000000)
  ) CLBLM_L_X68Y106_SLICE_X103Y106_DLUT (
.I0(CLBLM_L_X68Y108_SLICE_X103Y108_AQ),
.I1(CLBLM_L_X68Y106_SLICE_X103Y106_CQ),
.I2(CLBLM_L_X68Y106_SLICE_X103Y106_BQ),
.I3(CLBLM_L_X68Y108_SLICE_X103Y108_A5Q),
.I4(CLBLM_L_X68Y106_SLICE_X103Y106_B5Q),
.I5(CLBLM_L_X68Y105_SLICE_X102Y105_CQ),
.O5(CLBLM_L_X68Y106_SLICE_X103Y106_DO5),
.O6(CLBLM_L_X68Y106_SLICE_X103Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h70f08000f0f00000)
  ) CLBLM_L_X68Y106_SLICE_X103Y106_CLUT (
.I0(CLBLM_L_X68Y108_SLICE_X103Y108_AQ),
.I1(CLBLM_L_X70Y106_SLICE_X104Y106_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X68Y108_SLICE_X103Y108_A5Q),
.I4(CLBLM_L_X68Y106_SLICE_X103Y106_CQ),
.I5(CLBLM_L_X68Y105_SLICE_X102Y105_CQ),
.O5(CLBLM_L_X68Y106_SLICE_X103Y106_CO5),
.O6(CLBLM_L_X68Y106_SLICE_X103Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaa22aaaaf011f0)
  ) CLBLM_L_X68Y106_SLICE_X103Y106_BLUT (
.I0(CLBLM_L_X68Y106_SLICE_X103Y106_B5Q),
.I1(CLBLM_L_X68Y106_SLICE_X103Y106_BQ),
.I2(CLBLM_L_X68Y106_SLICE_X103Y106_CQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X68Y106_SLICE_X103Y106_AO5),
.I5(1'b1),
.O5(CLBLM_L_X68Y106_SLICE_X103Y106_BO5),
.O6(CLBLM_L_X68Y106_SLICE_X103Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h880088007fffffff)
  ) CLBLM_L_X68Y106_SLICE_X103Y106_ALUT (
.I0(CLBLM_L_X68Y108_SLICE_X103Y108_A5Q),
.I1(CLBLM_L_X70Y106_SLICE_X104Y106_BQ),
.I2(CLBLM_L_X68Y106_SLICE_X103Y106_CQ),
.I3(CLBLM_L_X68Y108_SLICE_X103Y108_AQ),
.I4(CLBLM_L_X68Y105_SLICE_X102Y105_CQ),
.I5(1'b1),
.O5(CLBLM_L_X68Y106_SLICE_X103Y106_AO5),
.O6(CLBLM_L_X68Y106_SLICE_X103Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0f0e0f0e0)
  ) CLBLM_L_X68Y107_SLICE_X102Y107_DLUT (
.I0(CLBLM_L_X68Y102_SLICE_X102Y102_CQ),
.I1(CLBLM_R_X67Y109_SLICE_X100Y109_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_R_X65Y106_SLICE_X98Y106_CQ),
.I4(1'b1),
.I5(CLBLL_R_X71Y108_SLICE_X106Y108_BQ),
.O5(CLBLM_L_X68Y107_SLICE_X102Y107_DO5),
.O6(CLBLM_L_X68Y107_SLICE_X102Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff01ff00ff54ff)
  ) CLBLM_L_X68Y107_SLICE_X102Y107_CLUT (
.I0(CLBLM_L_X68Y106_SLICE_X102Y106_AO6),
.I1(CLBLM_L_X72Y118_SLICE_X109Y118_BQ),
.I2(CLBLM_L_X74Y109_SLICE_X113Y109_A5Q),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X68Y107_SLICE_X102Y107_DO6),
.I5(CLBLM_L_X72Y105_SLICE_X108Y105_CQ),
.O5(CLBLM_L_X68Y107_SLICE_X102Y107_CO5),
.O6(CLBLM_L_X68Y107_SLICE_X102Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccfcfcccccfdf)
  ) CLBLM_L_X68Y107_SLICE_X102Y107_BLUT (
.I0(CLBLM_L_X72Y118_SLICE_X109Y118_BQ),
.I1(CLBLM_L_X68Y107_SLICE_X103Y107_BO6),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_R_X65Y106_SLICE_X98Y106_CQ),
.I4(CLBLM_L_X68Y106_SLICE_X102Y106_BO6),
.I5(CLBLM_L_X74Y109_SLICE_X113Y109_A5Q),
.O5(CLBLM_L_X68Y107_SLICE_X102Y107_BO5),
.O6(CLBLM_L_X68Y107_SLICE_X102Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f1f0f5f0f5f)
  ) CLBLM_L_X68Y107_SLICE_X102Y107_ALUT (
.I0(CLBLM_L_X72Y105_SLICE_X108Y105_CQ),
.I1(CLBLM_R_X67Y109_SLICE_X100Y109_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLL_R_X71Y108_SLICE_X106Y108_BQ),
.I4(CLBLM_L_X68Y102_SLICE_X102Y102_CQ),
.I5(1'b1),
.O5(CLBLM_L_X68Y107_SLICE_X102Y107_AO5),
.O6(CLBLM_L_X68Y107_SLICE_X102Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf4f4d8d8f4f4d8dd)
  ) CLBLM_L_X68Y107_SLICE_X103Y107_DLUT (
.I0(CLBLM_L_X68Y106_SLICE_X103Y106_CQ),
.I1(CLBLM_L_X70Y106_SLICE_X104Y106_BO6),
.I2(CLBLM_L_X68Y106_SLICE_X103Y106_B5Q),
.I3(CLBLM_L_X68Y109_SLICE_X103Y109_B5Q),
.I4(CLBLM_L_X68Y106_SLICE_X103Y106_BQ),
.I5(CLBLM_L_X68Y109_SLICE_X103Y109_BQ),
.O5(CLBLM_L_X68Y107_SLICE_X103Y107_DO5),
.O6(CLBLM_L_X68Y107_SLICE_X103Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X68Y107_SLICE_X103Y107_CLUT (
.I0(CLBLM_L_X68Y102_SLICE_X102Y102_CQ),
.I1(CLBLM_L_X72Y105_SLICE_X108Y105_CQ),
.I2(CLBLM_L_X64Y104_SLICE_X96Y104_CQ),
.I3(CLBLM_L_X74Y109_SLICE_X113Y109_A5Q),
.I4(CLBLM_R_X65Y100_SLICE_X98Y100_AQ),
.I5(CLBLM_L_X72Y118_SLICE_X109Y118_BQ),
.O5(CLBLM_L_X68Y107_SLICE_X103Y107_CO5),
.O6(CLBLM_L_X68Y107_SLICE_X103Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaabaaaaabbf)
  ) CLBLM_L_X68Y107_SLICE_X103Y107_BLUT (
.I0(CLBLM_L_X68Y107_SLICE_X102Y107_CO6),
.I1(CLBLL_R_X71Y108_SLICE_X106Y108_BQ),
.I2(CLBLM_L_X70Y104_SLICE_X105Y104_BQ),
.I3(CLBLM_R_X67Y109_SLICE_X100Y109_BQ),
.I4(CLBLM_L_X68Y107_SLICE_X103Y107_CO6),
.I5(CLBLM_R_X65Y106_SLICE_X98Y106_CQ),
.O5(CLBLM_L_X68Y107_SLICE_X103Y107_BO5),
.O6(CLBLM_L_X68Y107_SLICE_X103Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffbff33ff33ff)
  ) CLBLM_L_X68Y107_SLICE_X103Y107_ALUT (
.I0(CLBLM_L_X64Y104_SLICE_X96Y104_CQ),
.I1(CLBLM_L_X70Y108_SLICE_X105Y108_AO6),
.I2(CLBLM_L_X70Y104_SLICE_X105Y104_BQ),
.I3(CLBLM_L_X68Y107_SLICE_X102Y107_AO6),
.I4(CLBLM_R_X65Y100_SLICE_X98Y100_AQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X68Y107_SLICE_X103Y107_AO5),
.O6(CLBLM_L_X68Y107_SLICE_X103Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y108_SLICE_X102Y108_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y108_SLICE_X102Y108_AO5),
.Q(CLBLM_L_X68Y108_SLICE_X102Y108_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y108_SLICE_X102Y108_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y108_SLICE_X102Y108_BO5),
.Q(CLBLM_L_X68Y108_SLICE_X102Y108_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y108_SLICE_X102Y108_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y108_SLICE_X102Y108_AO6),
.Q(CLBLM_L_X68Y108_SLICE_X102Y108_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y108_SLICE_X102Y108_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y108_SLICE_X102Y108_BO6),
.Q(CLBLM_L_X68Y108_SLICE_X102Y108_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y108_SLICE_X102Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y108_SLICE_X102Y108_DO5),
.O6(CLBLM_L_X68Y108_SLICE_X102Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff88822282)
  ) CLBLM_L_X68Y108_SLICE_X102Y108_CLUT (
.I0(CLBLM_L_X70Y106_SLICE_X105Y106_DO6),
.I1(CLBLM_L_X68Y108_SLICE_X102Y108_AQ),
.I2(CLBLM_L_X68Y108_SLICE_X102Y108_BQ),
.I3(CLBLM_L_X68Y108_SLICE_X102Y108_A5Q),
.I4(CLBLM_L_X68Y108_SLICE_X102Y108_B5Q),
.I5(CLBLM_L_X68Y108_SLICE_X103Y108_BQ),
.O5(CLBLM_L_X68Y108_SLICE_X102Y108_CO5),
.O6(CLBLM_L_X68Y108_SLICE_X102Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f505f500ccccccc)
  ) CLBLM_L_X68Y108_SLICE_X102Y108_BLUT (
.I0(CLBLM_L_X68Y108_SLICE_X102Y108_B5Q),
.I1(CLBLM_L_X68Y108_SLICE_X102Y108_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X68Y109_SLICE_X102Y109_A5Q),
.I4(CLBLM_R_X67Y109_SLICE_X100Y109_DO5),
.I5(1'b1),
.O5(CLBLM_L_X68Y108_SLICE_X102Y108_BO5),
.O6(CLBLM_L_X68Y108_SLICE_X102Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cccf0cc33aaccaa)
  ) CLBLM_L_X68Y108_SLICE_X102Y108_ALUT (
.I0(CLBLM_L_X68Y108_SLICE_X102Y108_B5Q),
.I1(CLBLM_L_X68Y108_SLICE_X102Y108_A5Q),
.I2(CLBLM_L_X68Y108_SLICE_X102Y108_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X70Y106_SLICE_X105Y106_DO6),
.I5(1'b1),
.O5(CLBLM_L_X68Y108_SLICE_X102Y108_AO5),
.O6(CLBLM_L_X68Y108_SLICE_X102Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y108_SLICE_X103Y108_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y108_SLICE_X103Y108_AO5),
.Q(CLBLM_L_X68Y108_SLICE_X103Y108_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y108_SLICE_X103Y108_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y108_SLICE_X103Y108_AO6),
.Q(CLBLM_L_X68Y108_SLICE_X103Y108_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y108_SLICE_X103Y108_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y108_SLICE_X103Y108_BO6),
.Q(CLBLM_L_X68Y108_SLICE_X103Y108_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y108_SLICE_X103Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y108_SLICE_X103Y108_DO5),
.O6(CLBLM_L_X68Y108_SLICE_X103Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2222222200000000)
  ) CLBLM_L_X68Y108_SLICE_X103Y108_CLUT (
.I0(CLBLM_L_X68Y106_SLICE_X103Y106_BQ),
.I1(CLBLM_L_X68Y106_SLICE_X103Y106_B5Q),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X68Y106_SLICE_X103Y106_CQ),
.O5(CLBLM_L_X68Y108_SLICE_X103Y108_CO5),
.O6(CLBLM_L_X68Y108_SLICE_X103Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h20f0000000f00000)
  ) CLBLM_L_X68Y108_SLICE_X103Y108_BLUT (
.I0(CLBLM_L_X68Y109_SLICE_X103Y109_B5Q),
.I1(CLBLM_L_X68Y109_SLICE_X103Y109_BQ),
.I2(CLBLM_L_X68Y108_SLICE_X102Y108_CO6),
.I3(CLBLM_L_X70Y106_SLICE_X105Y106_DO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X68Y108_SLICE_X103Y108_CO6),
.O5(CLBLM_L_X68Y108_SLICE_X103Y108_BO5),
.O6(CLBLM_L_X68Y108_SLICE_X103Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff0ff003cccf0f0)
  ) CLBLM_L_X68Y108_SLICE_X103Y108_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X68Y108_SLICE_X103Y108_A5Q),
.I2(CLBLM_L_X68Y108_SLICE_X103Y108_AQ),
.I3(CLBLM_L_X70Y106_SLICE_X104Y106_BQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLM_L_X68Y108_SLICE_X103Y108_AO5),
.O6(CLBLM_L_X68Y108_SLICE_X103Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y109_SLICE_X102Y109_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y109_SLICE_X102Y109_AO5),
.Q(CLBLM_L_X68Y109_SLICE_X102Y109_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y109_SLICE_X102Y109_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y109_SLICE_X102Y109_AO6),
.Q(CLBLM_L_X68Y109_SLICE_X102Y109_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h88000000f8f0f0f0)
  ) CLBLM_L_X68Y109_SLICE_X102Y109_DLUT (
.I0(CLBLM_R_X67Y110_SLICE_X101Y110_AQ),
.I1(CLBLM_L_X68Y109_SLICE_X102Y109_BO6),
.I2(CLBLM_R_X67Y110_SLICE_X101Y110_DQ),
.I3(CLBLM_L_X68Y109_SLICE_X102Y109_A5Q),
.I4(CLBLM_R_X65Y111_SLICE_X98Y111_AQ),
.I5(CLBLM_R_X67Y108_SLICE_X101Y108_AO5),
.O5(CLBLM_L_X68Y109_SLICE_X102Y109_DO5),
.O6(CLBLM_L_X68Y109_SLICE_X102Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0e0f0f0f0f0)
  ) CLBLM_L_X68Y109_SLICE_X102Y109_CLUT (
.I0(CLBLM_R_X65Y108_SLICE_X99Y108_AO6),
.I1(CLBLM_L_X68Y109_SLICE_X102Y109_BO5),
.I2(CLBLM_L_X70Y106_SLICE_X105Y106_DO6),
.I3(CLBLM_R_X65Y110_SLICE_X99Y110_CO6),
.I4(CLBLM_L_X68Y109_SLICE_X102Y109_DO6),
.I5(CLBLM_R_X67Y109_SLICE_X101Y109_DO6),
.O5(CLBLM_L_X68Y109_SLICE_X102Y109_CO5),
.O6(CLBLM_L_X68Y109_SLICE_X102Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0c0c0c02000000)
  ) CLBLM_L_X68Y109_SLICE_X102Y109_BLUT (
.I0(CLBLM_R_X67Y109_SLICE_X101Y109_AQ),
.I1(CLBLM_L_X68Y108_SLICE_X102Y108_A5Q),
.I2(CLBLM_L_X68Y108_SLICE_X102Y108_AQ),
.I3(CLBLM_R_X65Y109_SLICE_X99Y109_A5Q),
.I4(CLBLM_L_X68Y109_SLICE_X102Y109_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X68Y109_SLICE_X102Y109_BO5),
.O6(CLBLM_L_X68Y109_SLICE_X102Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa55004e4ee4e4)
  ) CLBLM_L_X68Y109_SLICE_X102Y109_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_R_X65Y109_SLICE_X99Y109_A5Q),
.I2(CLBLM_R_X67Y109_SLICE_X100Y109_DO5),
.I3(CLBLM_L_X70Y114_SLICE_X104Y114_AQ),
.I4(CLBLM_L_X68Y109_SLICE_X102Y109_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X68Y109_SLICE_X102Y109_AO5),
.O6(CLBLM_L_X68Y109_SLICE_X102Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y109_SLICE_X103Y109_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y109_SLICE_X103Y109_BO5),
.Q(CLBLM_L_X68Y109_SLICE_X103Y109_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y109_SLICE_X103Y109_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y109_SLICE_X103Y109_AO6),
.Q(CLBLM_L_X68Y109_SLICE_X103Y109_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y109_SLICE_X103Y109_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y109_SLICE_X103Y109_BO6),
.Q(CLBLM_L_X68Y109_SLICE_X103Y109_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y109_SLICE_X103Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y109_SLICE_X103Y109_DO5),
.O6(CLBLM_L_X68Y109_SLICE_X103Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y109_SLICE_X103Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y109_SLICE_X103Y109_CO5),
.O6(CLBLM_L_X68Y109_SLICE_X103Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaa6caaaaf05af0)
  ) CLBLM_L_X68Y109_SLICE_X103Y109_BLUT (
.I0(CLBLM_L_X68Y109_SLICE_X103Y109_B5Q),
.I1(CLBLM_L_X68Y109_SLICE_X103Y109_BQ),
.I2(CLBLM_L_X68Y106_SLICE_X103Y106_BQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X68Y106_SLICE_X103Y106_AO5),
.I5(1'b1),
.O5(CLBLM_L_X68Y109_SLICE_X103Y109_BO5),
.O6(CLBLM_L_X68Y109_SLICE_X103Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3aaf3aaf0aaf0aa)
  ) CLBLM_L_X68Y109_SLICE_X103Y109_ALUT (
.I0(CLBLM_R_X67Y110_SLICE_X101Y110_DQ),
.I1(CLBLM_L_X70Y106_SLICE_X105Y106_DO6),
.I2(CLBLM_L_X68Y109_SLICE_X102Y109_CO6),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(1'b1),
.I5(CLBLM_L_X68Y109_SLICE_X103Y109_AQ),
.O5(CLBLM_L_X68Y109_SLICE_X103Y109_AO5),
.O6(CLBLM_L_X68Y109_SLICE_X103Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y112_SLICE_X102Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y112_SLICE_X102Y112_DO5),
.O6(CLBLM_L_X68Y112_SLICE_X102Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y112_SLICE_X102Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y112_SLICE_X102Y112_CO5),
.O6(CLBLM_L_X68Y112_SLICE_X102Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y112_SLICE_X102Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y112_SLICE_X102Y112_BO5),
.O6(CLBLM_L_X68Y112_SLICE_X102Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y112_SLICE_X102Y112_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y112_SLICE_X102Y112_AO5),
.O6(CLBLM_L_X68Y112_SLICE_X102Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y112_SLICE_X103Y112_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y112_SLICE_X106Y112_B5Q),
.Q(CLBLM_L_X68Y112_SLICE_X103Y112_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y112_SLICE_X103Y112_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X68Y112_SLICE_X103Y112_AQ),
.Q(CLBLM_L_X68Y112_SLICE_X103Y112_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y112_SLICE_X103Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y112_SLICE_X103Y112_DO5),
.O6(CLBLM_L_X68Y112_SLICE_X103Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y112_SLICE_X103Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y112_SLICE_X103Y112_CO5),
.O6(CLBLM_L_X68Y112_SLICE_X103Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y112_SLICE_X103Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y112_SLICE_X103Y112_BO5),
.O6(CLBLM_L_X68Y112_SLICE_X103Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y112_SLICE_X103Y112_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y112_SLICE_X103Y112_AO5),
.O6(CLBLM_L_X68Y112_SLICE_X103Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X68Y121_SLICE_X102Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y121_SLICE_X108Y121_AQ),
.Q(CLBLM_L_X68Y121_SLICE_X102Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y121_SLICE_X102Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y121_SLICE_X102Y121_DO5),
.O6(CLBLM_L_X68Y121_SLICE_X102Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y121_SLICE_X102Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y121_SLICE_X102Y121_CO5),
.O6(CLBLM_L_X68Y121_SLICE_X102Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y121_SLICE_X102Y121_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y121_SLICE_X102Y121_BO5),
.O6(CLBLM_L_X68Y121_SLICE_X102Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y121_SLICE_X102Y121_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y121_SLICE_X102Y121_AO5),
.O6(CLBLM_L_X68Y121_SLICE_X102Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y121_SLICE_X103Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y121_SLICE_X103Y121_DO5),
.O6(CLBLM_L_X68Y121_SLICE_X103Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y121_SLICE_X103Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y121_SLICE_X103Y121_CO5),
.O6(CLBLM_L_X68Y121_SLICE_X103Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y121_SLICE_X103Y121_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y121_SLICE_X103Y121_BO5),
.O6(CLBLM_L_X68Y121_SLICE_X103Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y121_SLICE_X103Y121_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y121_SLICE_X103Y121_AO5),
.O6(CLBLM_L_X68Y121_SLICE_X103Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y98_SLICE_X104Y98_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y99_SLICE_X104Y99_AQ),
.Q(CLBLM_L_X70Y98_SLICE_X104Y98_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y98_SLICE_X104Y98_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y98_SLICE_X104Y98_DO5),
.O6(CLBLM_L_X70Y98_SLICE_X104Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y98_SLICE_X104Y98_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y98_SLICE_X104Y98_CO5),
.O6(CLBLM_L_X70Y98_SLICE_X104Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y98_SLICE_X104Y98_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y98_SLICE_X104Y98_BO5),
.O6(CLBLM_L_X70Y98_SLICE_X104Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y98_SLICE_X104Y98_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y98_SLICE_X104Y98_AO5),
.O6(CLBLM_L_X70Y98_SLICE_X104Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y98_SLICE_X105Y98_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y98_SLICE_X105Y98_DO5),
.O6(CLBLM_L_X70Y98_SLICE_X105Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y98_SLICE_X105Y98_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y98_SLICE_X105Y98_CO5),
.O6(CLBLM_L_X70Y98_SLICE_X105Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y98_SLICE_X105Y98_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y98_SLICE_X105Y98_BO5),
.O6(CLBLM_L_X70Y98_SLICE_X105Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y98_SLICE_X105Y98_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y98_SLICE_X105Y98_AO5),
.O6(CLBLM_L_X70Y98_SLICE_X105Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y99_SLICE_X104Y99_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y101_SLICE_X105Y101_AQ),
.Q(CLBLM_L_X70Y99_SLICE_X104Y99_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5fffffff00000000)
  ) CLBLM_L_X70Y99_SLICE_X104Y99_DLUT (
.I0(CLBLM_L_X70Y100_SLICE_X105Y100_AQ),
.I1(1'b1),
.I2(CLBLM_L_X70Y99_SLICE_X104Y99_AQ),
.I3(CLBLM_L_X70Y100_SLICE_X105Y100_A5Q),
.I4(CLBLM_L_X70Y102_SLICE_X105Y102_CQ),
.I5(CLBLL_R_X71Y98_SLICE_X106Y98_A5Q),
.O5(CLBLM_L_X70Y99_SLICE_X104Y99_DO5),
.O6(CLBLM_L_X70Y99_SLICE_X104Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff000010ff1010)
  ) CLBLM_L_X70Y99_SLICE_X104Y99_CLUT (
.I0(CLBLM_L_X70Y99_SLICE_X104Y99_AO6),
.I1(CLBLM_L_X70Y99_SLICE_X105Y99_AO6),
.I2(CLBLM_L_X70Y100_SLICE_X104Y100_DO6),
.I3(CLBLL_R_X71Y101_SLICE_X106Y101_DO6),
.I4(CLBLM_L_X70Y99_SLICE_X104Y99_DO6),
.I5(CLBLM_L_X70Y99_SLICE_X104Y99_BO6),
.O5(CLBLM_L_X70Y99_SLICE_X104Y99_CO5),
.O6(CLBLM_L_X70Y99_SLICE_X104Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heca0000000000000)
  ) CLBLM_L_X70Y99_SLICE_X104Y99_BLUT (
.I0(CLBLM_L_X70Y100_SLICE_X104Y100_CQ),
.I1(CLBLM_L_X70Y101_SLICE_X104Y101_CQ),
.I2(CLBLM_L_X70Y101_SLICE_X104Y101_AQ),
.I3(CLBLL_R_X71Y100_SLICE_X106Y100_BQ),
.I4(CLBLM_L_X70Y100_SLICE_X105Y100_AQ),
.I5(CLBLM_L_X70Y100_SLICE_X105Y100_A5Q),
.O5(CLBLM_L_X70Y99_SLICE_X104Y99_BO5),
.O6(CLBLM_L_X70Y99_SLICE_X104Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000c8c000008800)
  ) CLBLM_L_X70Y99_SLICE_X104Y99_ALUT (
.I0(CLBLM_L_X70Y101_SLICE_X104Y101_BQ),
.I1(CLBLM_L_X70Y100_SLICE_X105Y100_A5Q),
.I2(CLBLM_L_X70Y99_SLICE_X104Y99_AQ),
.I3(CLBLM_L_X60Y97_SLICE_X90Y97_BQ),
.I4(CLBLM_L_X70Y100_SLICE_X105Y100_AQ),
.I5(CLBLM_L_X70Y99_SLICE_X105Y99_CQ),
.O5(CLBLM_L_X70Y99_SLICE_X104Y99_AO5),
.O6(CLBLM_L_X70Y99_SLICE_X104Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y99_SLICE_X105Y99_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y99_SLICE_X105Y99_BO6),
.Q(CLBLM_L_X70Y99_SLICE_X105Y99_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y99_SLICE_X105Y99_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y99_SLICE_X105Y99_CO6),
.Q(CLBLM_L_X70Y99_SLICE_X105Y99_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y99_SLICE_X105Y99_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y99_SLICE_X105Y99_DO5),
.O6(CLBLM_L_X70Y99_SLICE_X105Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccf0ddf088f0)
  ) CLBLM_L_X70Y99_SLICE_X105Y99_CLUT (
.I0(CLBLM_L_X70Y103_SLICE_X105Y103_CO6),
.I1(CLBLM_L_X70Y99_SLICE_X105Y99_CQ),
.I2(CLBLM_L_X70Y99_SLICE_X105Y99_BQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I5(CLBLM_L_X70Y103_SLICE_X105Y103_DO5),
.O5(CLBLM_L_X70Y99_SLICE_X105Y99_CO5),
.O6(CLBLM_L_X70Y99_SLICE_X105Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddddfd588888a80)
  ) CLBLM_L_X70Y99_SLICE_X105Y99_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X70Y99_SLICE_X105Y99_BQ),
.I2(CLBLM_L_X70Y103_SLICE_X105Y103_CO6),
.I3(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I4(CLBLM_L_X70Y103_SLICE_X105Y103_DO6),
.I5(CLBLM_L_X70Y100_SLICE_X104Y100_CQ),
.O5(CLBLM_L_X70Y99_SLICE_X105Y99_BO5),
.O6(CLBLM_L_X70Y99_SLICE_X105Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f4f055550000)
  ) CLBLM_L_X70Y99_SLICE_X105Y99_ALUT (
.I0(CLBLM_L_X70Y100_SLICE_X105Y100_A5Q),
.I1(CLBLM_L_X70Y99_SLICE_X105Y99_BQ),
.I2(CLBLL_R_X71Y98_SLICE_X106Y98_A5Q),
.I3(CLBLM_L_X70Y101_SLICE_X105Y101_AQ),
.I4(CLBLM_L_X70Y100_SLICE_X105Y100_AQ),
.I5(1'b1),
.O5(CLBLM_L_X70Y99_SLICE_X105Y99_AO5),
.O6(CLBLM_L_X70Y99_SLICE_X105Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y100_SLICE_X104Y100_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X60Y97_SLICE_X90Y97_BQ),
.Q(CLBLM_L_X70Y100_SLICE_X104Y100_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y100_SLICE_X104Y100_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y100_SLICE_X104Y100_AO6),
.Q(CLBLM_L_X70Y100_SLICE_X104Y100_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y100_SLICE_X104Y100_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y100_SLICE_X104Y100_BO6),
.Q(CLBLM_L_X70Y100_SLICE_X104Y100_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y100_SLICE_X104Y100_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y100_SLICE_X104Y100_CO6),
.Q(CLBLM_L_X70Y100_SLICE_X104Y100_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff135fffff)
  ) CLBLM_L_X70Y100_SLICE_X104Y100_DLUT (
.I0(CLBLM_L_X70Y100_SLICE_X104Y100_BQ),
.I1(CLBLM_L_X70Y100_SLICE_X104Y100_AQ),
.I2(CLBLM_L_X70Y98_SLICE_X104Y98_AQ),
.I3(CLBLM_L_X70Y100_SLICE_X104Y100_A5Q),
.I4(CLBLM_L_X70Y100_SLICE_X105Y100_AQ),
.I5(CLBLM_L_X70Y100_SLICE_X105Y100_A5Q),
.O5(CLBLM_L_X70Y100_SLICE_X104Y100_DO5),
.O6(CLBLM_L_X70Y100_SLICE_X104Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ddf0ccf088f0)
  ) CLBLM_L_X70Y100_SLICE_X104Y100_CLUT (
.I0(CLBLM_L_X70Y103_SLICE_X104Y103_DO5),
.I1(CLBLM_L_X70Y100_SLICE_X104Y100_CQ),
.I2(CLBLM_L_X70Y100_SLICE_X104Y100_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X70Y103_SLICE_X105Y103_CO6),
.I5(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.O5(CLBLM_L_X70Y100_SLICE_X104Y100_CO5),
.O6(CLBLM_L_X70Y100_SLICE_X104Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdc8cdc8cffff0000)
  ) CLBLM_L_X70Y100_SLICE_X104Y100_BLUT (
.I0(CLBLM_L_X70Y103_SLICE_X105Y103_CO6),
.I1(CLBLM_L_X70Y100_SLICE_X104Y100_BQ),
.I2(CLBLM_L_X70Y103_SLICE_X104Y103_C5Q),
.I3(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I4(CLBLM_L_X70Y99_SLICE_X105Y99_CQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X70Y100_SLICE_X104Y100_BO5),
.O6(CLBLM_L_X70Y100_SLICE_X104Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3c0c0f7b3c480)
  ) CLBLM_L_X70Y100_SLICE_X104Y100_ALUT (
.I0(CLBLM_L_X70Y103_SLICE_X105Y103_CO6),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_L_X70Y100_SLICE_X104Y100_AQ),
.I3(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I4(CLBLM_L_X70Y101_SLICE_X104Y101_BQ),
.I5(CLBLM_L_X70Y103_SLICE_X104Y103_DO6),
.O5(CLBLM_L_X70Y100_SLICE_X104Y100_AO5),
.O6(CLBLM_L_X70Y100_SLICE_X104Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y100_SLICE_X105Y100_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y100_SLICE_X105Y100_AO5),
.Q(CLBLM_L_X70Y100_SLICE_X105Y100_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y100_SLICE_X105Y100_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y100_SLICE_X105Y100_BO5),
.Q(CLBLM_L_X70Y100_SLICE_X105Y100_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y100_SLICE_X105Y100_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y100_SLICE_X105Y100_AO6),
.Q(CLBLM_L_X70Y100_SLICE_X105Y100_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y100_SLICE_X105Y100_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y100_SLICE_X105Y100_BO6),
.Q(CLBLM_L_X70Y100_SLICE_X105Y100_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y100_SLICE_X105Y100_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y108_SLICE_X118Y108_AQ),
.Q(CLBLM_L_X70Y100_SLICE_X105Y100_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff8ff080ff0ff000)
  ) CLBLM_L_X70Y100_SLICE_X105Y100_DLUT (
.I0(CLBLM_L_X70Y101_SLICE_X104Y101_AO6),
.I1(CLBLM_L_X70Y100_SLICE_X105Y100_CQ),
.I2(CLBLL_R_X71Y100_SLICE_X106Y100_AO6),
.I3(CLBLM_L_X70Y100_SLICE_X105Y100_CO6),
.I4(CLBLL_R_X71Y100_SLICE_X106Y100_CO6),
.I5(CLBLL_R_X71Y101_SLICE_X107Y101_AQ),
.O5(CLBLM_L_X70Y100_SLICE_X105Y100_DO5),
.O6(CLBLM_L_X70Y100_SLICE_X105Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa000000c000c0)
  ) CLBLM_L_X70Y100_SLICE_X105Y100_CLUT (
.I0(CLBLM_L_X60Y99_SLICE_X90Y99_AQ),
.I1(CLBLL_R_X77Y108_SLICE_X118Y108_AQ),
.I2(CLBLL_R_X71Y101_SLICE_X106Y101_AQ),
.I3(CLBLM_L_X70Y100_SLICE_X105Y100_A5Q),
.I4(CLBLM_L_X70Y101_SLICE_X105Y101_BQ),
.I5(CLBLM_L_X70Y100_SLICE_X105Y100_AQ),
.O5(CLBLM_L_X70Y100_SLICE_X105Y100_CO5),
.O6(CLBLM_L_X70Y100_SLICE_X105Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f5f50500ccccccc)
  ) CLBLM_L_X70Y100_SLICE_X105Y100_BLUT (
.I0(CLBLM_L_X70Y100_SLICE_X105Y100_B5Q),
.I1(CLBLM_L_X70Y100_SLICE_X105Y100_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLL_R_X71Y100_SLICE_X106Y100_AO5),
.I4(CLBLL_R_X71Y98_SLICE_X106Y98_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X70Y100_SLICE_X105Y100_BO5),
.O6(CLBLM_L_X70Y100_SLICE_X105Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cfff00033aaccaa)
  ) CLBLM_L_X70Y100_SLICE_X105Y100_ALUT (
.I0(CLBLM_L_X70Y100_SLICE_X105Y100_B5Q),
.I1(CLBLM_R_X65Y103_SLICE_X99Y103_DO6),
.I2(CLBLM_L_X70Y100_SLICE_X105Y100_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X70Y100_SLICE_X105Y100_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X70Y100_SLICE_X105Y100_AO5),
.O6(CLBLM_L_X70Y100_SLICE_X105Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y101_SLICE_X104Y101_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y100_SLICE_X104Y100_A5Q),
.Q(CLBLM_L_X70Y101_SLICE_X104Y101_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y101_SLICE_X104Y101_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y101_SLICE_X104Y101_BO6),
.Q(CLBLM_L_X70Y101_SLICE_X104Y101_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y101_SLICE_X104Y101_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y101_SLICE_X104Y101_CO6),
.Q(CLBLM_L_X70Y101_SLICE_X104Y101_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfef2f1fdf0f0f0f0)
  ) CLBLM_L_X70Y101_SLICE_X104Y101_DLUT (
.I0(CLBLM_L_X70Y100_SLICE_X105Y100_BQ),
.I1(CLBLM_L_X70Y100_SLICE_X105Y100_A5Q),
.I2(CLBLM_R_X65Y102_SLICE_X99Y102_AQ),
.I3(CLBLM_L_X70Y100_SLICE_X105Y100_B5Q),
.I4(CLBLM_L_X70Y100_SLICE_X105Y100_AQ),
.I5(CLBLM_R_X65Y103_SLICE_X99Y103_DO6),
.O5(CLBLM_L_X70Y101_SLICE_X104Y101_DO5),
.O6(CLBLM_L_X70Y101_SLICE_X104Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfdf8fc0c0d080)
  ) CLBLM_L_X70Y101_SLICE_X104Y101_CLUT (
.I0(CLBLM_L_X70Y103_SLICE_X105Y103_CO5),
.I1(CLBLM_L_X70Y101_SLICE_X104Y101_CQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I4(CLBLM_L_X70Y103_SLICE_X104Y103_DO6),
.I5(CLBLM_L_X70Y100_SLICE_X104Y100_BQ),
.O5(CLBLM_L_X70Y101_SLICE_X104Y101_CO5),
.O6(CLBLM_L_X70Y101_SLICE_X104Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddfd5d8888a808)
  ) CLBLM_L_X70Y101_SLICE_X104Y101_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X70Y101_SLICE_X104Y101_BQ),
.I2(CLBLM_L_X70Y103_SLICE_X104Y103_C5Q),
.I3(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I4(CLBLL_R_X71Y103_SLICE_X106Y103_BO6),
.I5(CLBLL_R_X71Y101_SLICE_X106Y101_CQ),
.O5(CLBLM_L_X70Y101_SLICE_X104Y101_BO5),
.O6(CLBLM_L_X70Y101_SLICE_X104Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aaaa80000000)
  ) CLBLM_L_X70Y101_SLICE_X104Y101_ALUT (
.I0(CLBLM_L_X70Y100_SLICE_X105Y100_A5Q),
.I1(CLBLM_R_X65Y103_SLICE_X99Y103_DO6),
.I2(CLBLL_R_X71Y98_SLICE_X106Y98_A5Q),
.I3(CLBLM_L_X60Y97_SLICE_X90Y97_BQ),
.I4(CLBLM_L_X70Y100_SLICE_X105Y100_AQ),
.I5(1'b1),
.O5(CLBLM_L_X70Y101_SLICE_X104Y101_AO5),
.O6(CLBLM_L_X70Y101_SLICE_X104Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y101_SLICE_X105Y101_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y101_SLICE_X104Y101_AQ),
.Q(CLBLM_L_X70Y101_SLICE_X105Y101_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y101_SLICE_X105Y101_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y101_SLICE_X105Y101_BO6),
.Q(CLBLM_L_X70Y101_SLICE_X105Y101_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff80ff00)
  ) CLBLM_L_X70Y101_SLICE_X105Y101_DLUT (
.I0(CLBLM_L_X70Y101_SLICE_X105Y101_AO6),
.I1(CLBLL_R_X71Y98_SLICE_X106Y98_A5Q),
.I2(CLBLM_L_X70Y98_SLICE_X104Y98_AQ),
.I3(CLBLM_L_X70Y101_SLICE_X105Y101_AO5),
.I4(CLBLM_L_X70Y102_SLICE_X105Y102_BQ),
.I5(CLBLM_L_X70Y102_SLICE_X104Y102_BO6),
.O5(CLBLM_L_X70Y101_SLICE_X105Y101_DO5),
.O6(CLBLM_L_X70Y101_SLICE_X105Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffbfbb00000000)
  ) CLBLM_L_X70Y101_SLICE_X105Y101_CLUT (
.I0(CLBLM_L_X70Y100_SLICE_X105Y100_DO6),
.I1(CLBLM_L_X70Y99_SLICE_X104Y99_CO6),
.I2(CLBLL_R_X71Y102_SLICE_X106Y102_DO6),
.I3(CLBLM_L_X70Y99_SLICE_X105Y99_AO5),
.I4(CLBLM_L_X70Y101_SLICE_X105Y101_DO6),
.I5(CLBLM_R_X65Y103_SLICE_X99Y103_DO6),
.O5(CLBLM_L_X70Y101_SLICE_X105Y101_CO5),
.O6(CLBLM_L_X70Y101_SLICE_X105Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccacccaffff0000)
  ) CLBLM_L_X70Y101_SLICE_X105Y101_BLUT (
.I0(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I1(CLBLM_L_X70Y101_SLICE_X105Y101_BQ),
.I2(CLBLM_L_X70Y103_SLICE_X105Y103_CO5),
.I3(CLBLM_L_X70Y103_SLICE_X105Y103_DO5),
.I4(CLBLL_R_X71Y101_SLICE_X107Y101_AQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X70Y101_SLICE_X105Y101_BO5),
.O6(CLBLM_L_X70Y101_SLICE_X105Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000555500008000)
  ) CLBLM_L_X70Y101_SLICE_X105Y101_ALUT (
.I0(CLBLM_L_X70Y100_SLICE_X105Y100_A5Q),
.I1(CLBLL_R_X71Y98_SLICE_X106Y98_A5Q),
.I2(CLBLM_L_X70Y102_SLICE_X105Y102_AQ),
.I3(CLBLL_R_X71Y100_SLICE_X106Y100_BQ),
.I4(CLBLM_L_X70Y100_SLICE_X105Y100_AQ),
.I5(1'b1),
.O5(CLBLM_L_X70Y101_SLICE_X105Y101_AO5),
.O6(CLBLM_L_X70Y101_SLICE_X105Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y102_SLICE_X104Y102_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y102_SLICE_X104Y102_AO6),
.Q(CLBLM_L_X70Y102_SLICE_X104Y102_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y102_SLICE_X104Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y102_SLICE_X104Y102_DO5),
.O6(CLBLM_L_X70Y102_SLICE_X104Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y102_SLICE_X104Y102_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y102_SLICE_X104Y102_CO5),
.O6(CLBLM_L_X70Y102_SLICE_X104Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc000000000000000)
  ) CLBLM_L_X70Y102_SLICE_X104Y102_BLUT (
.I0(1'b1),
.I1(CLBLL_R_X71Y98_SLICE_X106Y98_A5Q),
.I2(CLBLM_L_X70Y102_SLICE_X104Y102_AQ),
.I3(CLBLM_L_X60Y97_SLICE_X90Y97_BQ),
.I4(CLBLM_L_X70Y100_SLICE_X105Y100_AQ),
.I5(CLBLM_L_X70Y100_SLICE_X105Y100_A5Q),
.O5(CLBLM_L_X70Y102_SLICE_X104Y102_BO5),
.O6(CLBLM_L_X70Y102_SLICE_X104Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd75a820fd75a820)
  ) CLBLM_L_X70Y102_SLICE_X104Y102_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X70Y104_SLICE_X104Y104_CO5),
.I2(CLBLM_L_X70Y102_SLICE_X104Y102_AQ),
.I3(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I4(CLBLM_L_X70Y101_SLICE_X105Y101_BQ),
.I5(1'b1),
.O5(CLBLM_L_X70Y102_SLICE_X104Y102_AO5),
.O6(CLBLM_L_X70Y102_SLICE_X104Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y102_SLICE_X105Y102_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y102_SLICE_X105Y102_AO6),
.Q(CLBLM_L_X70Y102_SLICE_X105Y102_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y102_SLICE_X105Y102_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y102_SLICE_X105Y102_BO6),
.Q(CLBLM_L_X70Y102_SLICE_X105Y102_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y102_SLICE_X105Y102_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y102_SLICE_X105Y102_CO6),
.Q(CLBLM_L_X70Y102_SLICE_X105Y102_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff0000ffff0000)
  ) CLBLM_L_X70Y102_SLICE_X105Y102_DLUT (
.I0(CLBLM_L_X70Y100_SLICE_X105Y100_AQ),
.I1(CLBLM_L_X70Y100_SLICE_X105Y100_A5Q),
.I2(CLBLM_R_X65Y103_SLICE_X99Y103_DO6),
.I3(CLBLL_R_X71Y98_SLICE_X106Y98_A5Q),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X60Y97_SLICE_X90Y97_BQ),
.O5(CLBLM_L_X70Y102_SLICE_X105Y102_DO5),
.O6(CLBLM_L_X70Y102_SLICE_X105Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcaffcc00ca00)
  ) CLBLM_L_X70Y102_SLICE_X105Y102_CLUT (
.I0(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I1(CLBLM_L_X70Y102_SLICE_X105Y102_CQ),
.I2(CLBLL_R_X71Y103_SLICE_X106Y103_BO5),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X70Y103_SLICE_X105Y103_DO5),
.I5(CLBLL_R_X71Y102_SLICE_X106Y102_CQ),
.O5(CLBLM_L_X70Y102_SLICE_X105Y102_CO5),
.O6(CLBLM_L_X70Y102_SLICE_X105Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfccc0caaaaaaaa)
  ) CLBLM_L_X70Y102_SLICE_X105Y102_BLUT (
.I0(CLBLM_L_X70Y102_SLICE_X105Y102_CQ),
.I1(CLBLM_L_X70Y102_SLICE_X105Y102_BQ),
.I2(CLBLM_L_X70Y103_SLICE_X104Y103_C5Q),
.I3(CLBLL_R_X71Y103_SLICE_X106Y103_BO5),
.I4(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X70Y102_SLICE_X105Y102_BO5),
.O6(CLBLM_L_X70Y102_SLICE_X105Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f5a0cccccccc)
  ) CLBLM_L_X70Y102_SLICE_X105Y102_ALUT (
.I0(CLBLM_L_X70Y103_SLICE_X104Y103_DO6),
.I1(CLBLM_L_X70Y102_SLICE_X105Y102_BQ),
.I2(CLBLM_L_X70Y102_SLICE_X105Y102_AQ),
.I3(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I4(CLBLL_R_X71Y103_SLICE_X106Y103_BO6),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X70Y102_SLICE_X105Y102_AO5),
.O6(CLBLM_L_X70Y102_SLICE_X105Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y103_SLICE_X104Y103_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y103_SLICE_X104Y103_BO5),
.Q(CLBLM_L_X70Y103_SLICE_X104Y103_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y103_SLICE_X104Y103_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y103_SLICE_X104Y103_CO5),
.Q(CLBLM_L_X70Y103_SLICE_X104Y103_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y103_SLICE_X104Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y103_SLICE_X104Y103_AO6),
.Q(CLBLM_L_X70Y103_SLICE_X104Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y103_SLICE_X104Y103_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y103_SLICE_X104Y103_BO6),
.Q(CLBLM_L_X70Y103_SLICE_X104Y103_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y103_SLICE_X104Y103_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y103_SLICE_X104Y103_CO6),
.Q(CLBLM_L_X70Y103_SLICE_X104Y103_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefefefecfcfcfcf)
  ) CLBLM_L_X70Y103_SLICE_X104Y103_DLUT (
.I0(CLBLM_L_X70Y103_SLICE_X104Y103_C5Q),
.I1(CLBLM_L_X70Y103_SLICE_X104Y103_CQ),
.I2(CLBLM_L_X70Y103_SLICE_X104Y103_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y103_SLICE_X104Y103_DO5),
.O6(CLBLM_L_X70Y103_SLICE_X104Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ccff004400cccc)
  ) CLBLM_L_X70Y103_SLICE_X104Y103_CLUT (
.I0(CLBLM_L_X70Y103_SLICE_X104Y103_C5Q),
.I1(CLBLM_L_X70Y103_SLICE_X104Y103_CQ),
.I2(1'b1),
.I3(CLBLM_L_X70Y103_SLICE_X104Y103_BQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLM_L_X70Y103_SLICE_X104Y103_CO5),
.O6(CLBLM_L_X70Y103_SLICE_X104Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000030305f5fa0a0)
  ) CLBLM_L_X70Y103_SLICE_X104Y103_BLUT (
.I0(CLBLM_L_X70Y103_SLICE_X104Y103_B5Q),
.I1(CLBLM_L_X70Y103_SLICE_X104Y103_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(1'b1),
.I4(CLBLM_L_X70Y103_SLICE_X104Y103_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X70Y103_SLICE_X104Y103_BO5),
.O6(CLBLM_L_X70Y103_SLICE_X104Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffcccc3b3b0808)
  ) CLBLM_L_X70Y103_SLICE_X104Y103_ALUT (
.I0(CLBLM_L_X70Y103_SLICE_X104Y103_AQ),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_R_X65Y103_SLICE_X99Y103_DO6),
.I3(1'b1),
.I4(CLBLM_L_X70Y102_SLICE_X104Y102_AQ),
.I5(CLBLM_L_X70Y101_SLICE_X105Y101_CO6),
.O5(CLBLM_L_X70Y103_SLICE_X104Y103_AO5),
.O6(CLBLM_L_X70Y103_SLICE_X104Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y103_SLICE_X105Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y103_SLICE_X105Y103_AO6),
.Q(CLBLM_L_X70Y103_SLICE_X105Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y103_SLICE_X105Y103_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y103_SLICE_X105Y103_BO6),
.Q(CLBLM_L_X70Y103_SLICE_X105Y103_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffccff33ff33ff)
  ) CLBLM_L_X70Y103_SLICE_X105Y103_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X70Y103_SLICE_X104Y103_BQ),
.I2(1'b1),
.I3(CLBLM_L_X70Y103_SLICE_X104Y103_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y103_SLICE_X105Y103_DO5),
.O6(CLBLM_L_X70Y103_SLICE_X105Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f3f33f3f3f3f)
  ) CLBLM_L_X70Y103_SLICE_X105Y103_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X70Y104_SLICE_X104Y104_A5Q),
.I2(CLBLM_L_X70Y103_SLICE_X104Y103_B5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y103_SLICE_X105Y103_CO5),
.O6(CLBLM_L_X70Y103_SLICE_X105Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4cb30000cc330000)
  ) CLBLM_L_X70Y103_SLICE_X105Y103_BLUT (
.I0(CLBLM_L_X70Y103_SLICE_X104Y103_C5Q),
.I1(CLBLM_L_X70Y103_SLICE_X105Y103_BQ),
.I2(CLBLM_L_X70Y103_SLICE_X104Y103_B5Q),
.I3(CLBLL_R_X79Y99_SLICE_X122Y99_AO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X70Y104_SLICE_X104Y104_A5Q),
.O5(CLBLM_L_X70Y103_SLICE_X105Y103_BO5),
.O6(CLBLM_L_X70Y103_SLICE_X105Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdf80ccccff00cccc)
  ) CLBLM_L_X70Y103_SLICE_X105Y103_ALUT (
.I0(CLBLM_L_X70Y103_SLICE_X104Y103_C5Q),
.I1(CLBLM_L_X70Y103_SLICE_X105Y103_BQ),
.I2(CLBLM_L_X70Y103_SLICE_X104Y103_B5Q),
.I3(CLBLM_L_X70Y103_SLICE_X105Y103_AQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X70Y104_SLICE_X104Y104_A5Q),
.O5(CLBLM_L_X70Y103_SLICE_X105Y103_AO5),
.O6(CLBLM_L_X70Y103_SLICE_X105Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y104_SLICE_X104Y104_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y104_SLICE_X104Y104_CO6),
.Q(CLBLM_L_X70Y104_SLICE_X104Y104_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y104_SLICE_X104Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y104_SLICE_X104Y104_AO6),
.Q(CLBLM_L_X70Y104_SLICE_X104Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y104_SLICE_X104Y104_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y104_SLICE_X104Y104_BO6),
.Q(CLBLM_L_X70Y104_SLICE_X104Y104_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y104_SLICE_X104Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y104_SLICE_X104Y104_DO5),
.O6(CLBLM_L_X70Y104_SLICE_X104Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5fa0f5a0f0000000)
  ) CLBLM_L_X70Y104_SLICE_X104Y104_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(1'b1),
.I2(CLBLM_L_X70Y104_SLICE_X104Y104_A5Q),
.I3(CLBLM_L_X70Y103_SLICE_X104Y103_B5Q),
.I4(CLBLM_L_X70Y103_SLICE_X104Y103_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X70Y104_SLICE_X104Y104_CO5),
.O6(CLBLM_L_X70Y104_SLICE_X104Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a5ccccf0f0f0f0)
  ) CLBLM_L_X70Y104_SLICE_X104Y104_BLUT (
.I0(CLBLM_L_X70Y105_SLICE_X105Y105_A5Q),
.I1(CLBLM_L_X70Y104_SLICE_X104Y104_BQ),
.I2(CLBLM_L_X70Y104_SLICE_X104Y104_AQ),
.I3(1'b1),
.I4(CLBLM_L_X70Y104_SLICE_X104Y104_CO5),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X70Y104_SLICE_X104Y104_BO5),
.O6(CLBLM_L_X70Y104_SLICE_X104Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8f0aaaaf0f0aaaa)
  ) CLBLM_L_X70Y104_SLICE_X104Y104_ALUT (
.I0(CLBLM_L_X70Y105_SLICE_X105Y105_A5Q),
.I1(CLBLM_L_X70Y103_SLICE_X104Y103_C5Q),
.I2(CLBLM_L_X70Y104_SLICE_X104Y104_AQ),
.I3(CLBLM_L_X70Y103_SLICE_X104Y103_B5Q),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X70Y104_SLICE_X104Y104_A5Q),
.O5(CLBLM_L_X70Y104_SLICE_X104Y104_AO5),
.O6(CLBLM_L_X70Y104_SLICE_X104Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y104_SLICE_X105Y104_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y104_SLICE_X105Y104_DO5),
.Q(CLBLM_L_X70Y104_SLICE_X105Y104_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y104_SLICE_X105Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y104_SLICE_X105Y104_AO6),
.Q(CLBLM_L_X70Y104_SLICE_X105Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y104_SLICE_X105Y104_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y104_SLICE_X105Y104_BO6),
.Q(CLBLM_L_X70Y104_SLICE_X105Y104_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y104_SLICE_X105Y104_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y104_SLICE_X105Y104_CO6),
.Q(CLBLM_L_X70Y104_SLICE_X105Y104_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y104_SLICE_X105Y104_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y104_SLICE_X105Y104_DO6),
.Q(CLBLM_L_X70Y104_SLICE_X105Y104_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaaccf099f0aa)
  ) CLBLM_L_X70Y104_SLICE_X105Y104_DLUT (
.I0(CLBLM_L_X70Y104_SLICE_X105Y104_DQ),
.I1(CLBLM_L_X70Y104_SLICE_X105Y104_CQ),
.I2(CLBLM_L_X70Y104_SLICE_X105Y104_D5Q),
.I3(CLBLM_L_X70Y102_SLICE_X105Y102_DO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLM_L_X70Y104_SLICE_X105Y104_DO5),
.O6(CLBLM_L_X70Y104_SLICE_X105Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3caaccaaccaaccaa)
  ) CLBLM_L_X70Y104_SLICE_X105Y104_CLUT (
.I0(CLBLM_L_X70Y104_SLICE_X105Y104_BQ),
.I1(CLBLM_L_X70Y104_SLICE_X105Y104_CQ),
.I2(CLBLM_L_X70Y103_SLICE_X104Y103_B5Q),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X70Y104_SLICE_X104Y104_A5Q),
.I5(CLBLM_L_X70Y103_SLICE_X104Y103_C5Q),
.O5(CLBLM_L_X70Y104_SLICE_X105Y104_CO5),
.O6(CLBLM_L_X70Y104_SLICE_X105Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8d8dd8d8d8d8d8d8)
  ) CLBLM_L_X70Y104_SLICE_X105Y104_BLUT (
.I0(CLBLM_L_X70Y102_SLICE_X105Y102_DO6),
.I1(CLBLM_L_X70Y104_SLICE_X105Y104_BQ),
.I2(CLBLM_L_X70Y104_SLICE_X105Y104_AQ),
.I3(1'b1),
.I4(CLBLM_L_X70Y103_SLICE_X105Y103_AQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X70Y104_SLICE_X105Y104_BO5),
.O6(CLBLM_L_X70Y104_SLICE_X105Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55aa005ff50aa0)
  ) CLBLM_L_X70Y104_SLICE_X105Y104_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(1'b1),
.I2(CLBLM_L_X70Y104_SLICE_X105Y104_AQ),
.I3(CLBLM_L_X70Y101_SLICE_X105Y101_CO6),
.I4(CLBLM_L_X70Y103_SLICE_X105Y103_AQ),
.I5(CLBLM_L_X70Y101_SLICE_X104Y101_AO5),
.O5(CLBLM_L_X70Y104_SLICE_X105Y104_AO5),
.O6(CLBLM_L_X70Y104_SLICE_X105Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y105_SLICE_X104Y105_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y105_SLICE_X104Y105_AO6),
.Q(CLBLM_L_X70Y105_SLICE_X104Y105_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y105_SLICE_X104Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y105_SLICE_X104Y105_DO5),
.O6(CLBLM_L_X70Y105_SLICE_X104Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haf0faf0faa00aa00)
  ) CLBLM_L_X70Y105_SLICE_X104Y105_CLUT (
.I0(CLBLM_L_X68Y103_SLICE_X102Y103_AQ),
.I1(1'b1),
.I2(CLBLM_L_X72Y104_SLICE_X108Y104_DQ),
.I3(CLBLM_L_X70Y106_SLICE_X104Y106_AQ),
.I4(1'b1),
.I5(CLBLM_L_X70Y106_SLICE_X104Y106_BQ),
.O5(CLBLM_L_X70Y105_SLICE_X104Y105_CO5),
.O6(CLBLM_L_X70Y105_SLICE_X104Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f007f00ff00ff00)
  ) CLBLM_L_X70Y105_SLICE_X104Y105_BLUT (
.I0(CLBLM_L_X68Y106_SLICE_X103Y106_DO6),
.I1(CLBLM_L_X68Y109_SLICE_X103Y109_B5Q),
.I2(CLBLM_L_X70Y105_SLICE_X104Y105_AQ),
.I3(CLBLM_L_X70Y106_SLICE_X104Y106_BQ),
.I4(1'b1),
.I5(CLBLM_L_X68Y109_SLICE_X103Y109_BQ),
.O5(CLBLM_L_X70Y105_SLICE_X104Y105_BO5),
.O6(CLBLM_L_X70Y105_SLICE_X104Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf4b0ff00f0f0ff00)
  ) CLBLM_L_X70Y105_SLICE_X104Y105_ALUT (
.I0(CLBLM_L_X68Y109_SLICE_X103Y109_B5Q),
.I1(CLBLM_L_X68Y109_SLICE_X103Y109_BQ),
.I2(CLBLM_L_X70Y105_SLICE_X104Y105_AQ),
.I3(CLBLM_L_X70Y105_SLICE_X105Y105_BQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X68Y108_SLICE_X103Y108_CO6),
.O5(CLBLM_L_X70Y105_SLICE_X104Y105_AO5),
.O6(CLBLM_L_X70Y105_SLICE_X104Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y105_SLICE_X105Y105_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y105_SLICE_X105Y105_AO5),
.Q(CLBLM_L_X70Y105_SLICE_X105Y105_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y105_SLICE_X105Y105_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y105_SLICE_X105Y105_AO6),
.Q(CLBLM_L_X70Y105_SLICE_X105Y105_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y105_SLICE_X105Y105_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y105_SLICE_X105Y105_BO6),
.Q(CLBLM_L_X70Y105_SLICE_X105Y105_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y105_SLICE_X105Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y105_SLICE_X105Y105_DO5),
.O6(CLBLM_L_X70Y105_SLICE_X105Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y105_SLICE_X105Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y105_SLICE_X105Y105_CO5),
.O6(CLBLM_L_X70Y105_SLICE_X105Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2020a02020202020)
  ) CLBLM_L_X70Y105_SLICE_X105Y105_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X70Y105_SLICE_X104Y105_BO6),
.I2(CLBLM_L_X72Y104_SLICE_X109Y104_DO6),
.I3(CLBLM_L_X68Y108_SLICE_X103Y108_CO6),
.I4(CLBLM_L_X68Y109_SLICE_X103Y109_B5Q),
.I5(CLBLM_L_X68Y109_SLICE_X103Y109_BQ),
.O5(CLBLM_L_X70Y105_SLICE_X105Y105_BO5),
.O6(CLBLM_L_X70Y105_SLICE_X105Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h555500004ee44ee4)
  ) CLBLM_L_X70Y105_SLICE_X105Y105_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X70Y104_SLICE_X105Y104_D5Q),
.I2(CLBLM_L_X70Y105_SLICE_X105Y105_A5Q),
.I3(CLBLM_L_X70Y101_SLICE_X104Y101_AO5),
.I4(CLBLL_R_X75Y122_SLICE_X115Y122_AQ),
.I5(1'b1),
.O5(CLBLM_L_X70Y105_SLICE_X105Y105_AO5),
.O6(CLBLM_L_X70Y105_SLICE_X105Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y106_SLICE_X104Y106_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y106_SLICE_X104Y106_AQ),
.Q(CLBLM_L_X70Y106_SLICE_X104Y106_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y106_SLICE_X104Y106_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y106_SLICE_X104Y106_AO6),
.Q(CLBLM_L_X70Y106_SLICE_X104Y106_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y106_SLICE_X104Y106_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y106_SLICE_X105Y106_A5Q),
.Q(CLBLM_L_X70Y106_SLICE_X104Y106_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffff00)
  ) CLBLM_L_X70Y106_SLICE_X104Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X70Y106_SLICE_X104Y106_A5Q),
.I4(CLBLM_L_X70Y106_SLICE_X105Y106_A5Q),
.I5(CLBLM_L_X70Y106_SLICE_X104Y106_AQ),
.O5(CLBLM_L_X70Y106_SLICE_X104Y106_DO5),
.O6(CLBLM_L_X70Y106_SLICE_X104Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffdfffdf00000000)
  ) CLBLM_L_X70Y106_SLICE_X104Y106_CLUT (
.I0(CLBLM_L_X68Y105_SLICE_X103Y105_AQ),
.I1(CLBLM_L_X68Y109_SLICE_X103Y109_B5Q),
.I2(CLBLM_L_X68Y106_SLICE_X103Y106_DO6),
.I3(CLBLM_L_X68Y109_SLICE_X103Y109_BQ),
.I4(1'b1),
.I5(CLBLM_L_X70Y106_SLICE_X104Y106_AQ),
.O5(CLBLM_L_X70Y106_SLICE_X104Y106_CO5),
.O6(CLBLM_L_X70Y106_SLICE_X104Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f00ff55553333)
  ) CLBLM_L_X70Y106_SLICE_X104Y106_BLUT (
.I0(CLBLM_L_X70Y106_SLICE_X105Y106_AQ),
.I1(CLBLM_L_X68Y105_SLICE_X103Y105_AQ),
.I2(CLBLM_L_X70Y105_SLICE_X104Y105_AQ),
.I3(CLBLM_L_X70Y106_SLICE_X105Y106_BQ),
.I4(CLBLM_L_X68Y109_SLICE_X103Y109_B5Q),
.I5(CLBLM_L_X68Y109_SLICE_X103Y109_BQ),
.O5(CLBLM_L_X70Y106_SLICE_X104Y106_BO5),
.O6(CLBLM_L_X70Y106_SLICE_X104Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000040404)
  ) CLBLM_L_X70Y106_SLICE_X104Y106_ALUT (
.I0(CLBLM_L_X70Y106_SLICE_X105Y106_A5Q),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_L_X70Y106_SLICE_X104Y106_AQ),
.I3(CLBLM_L_X68Y105_SLICE_X102Y105_CQ),
.I4(CLBLM_L_X68Y106_SLICE_X103Y106_AO6),
.I5(CLBLM_L_X70Y106_SLICE_X104Y106_A5Q),
.O5(CLBLM_L_X70Y106_SLICE_X104Y106_AO5),
.O6(CLBLM_L_X70Y106_SLICE_X104Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y106_SLICE_X105Y106_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y106_SLICE_X104Y106_A5Q),
.Q(CLBLM_L_X70Y106_SLICE_X105Y106_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y106_SLICE_X105Y106_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y106_SLICE_X105Y106_AO6),
.Q(CLBLM_L_X70Y106_SLICE_X105Y106_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y106_SLICE_X105Y106_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y106_SLICE_X105Y106_BO6),
.Q(CLBLM_L_X70Y106_SLICE_X105Y106_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff3fffff00000000)
  ) CLBLM_L_X70Y106_SLICE_X105Y106_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X68Y109_SLICE_X103Y109_BQ),
.I2(CLBLM_L_X70Y106_SLICE_X105Y106_BQ),
.I3(CLBLM_L_X68Y109_SLICE_X103Y109_B5Q),
.I4(CLBLM_L_X68Y106_SLICE_X103Y106_DO6),
.I5(CLBLM_L_X70Y106_SLICE_X105Y106_A5Q),
.O5(CLBLM_L_X70Y106_SLICE_X105Y106_DO5),
.O6(CLBLM_L_X70Y106_SLICE_X105Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa2aaaaaaa2aaaaa)
  ) CLBLM_L_X70Y106_SLICE_X105Y106_CLUT (
.I0(CLBLM_L_X70Y106_SLICE_X104Y106_A5Q),
.I1(CLBLM_L_X68Y109_SLICE_X103Y109_B5Q),
.I2(CLBLM_L_X68Y106_SLICE_X103Y106_DO6),
.I3(CLBLM_L_X68Y109_SLICE_X103Y109_BQ),
.I4(CLBLM_L_X70Y106_SLICE_X105Y106_AQ),
.I5(1'b1),
.O5(CLBLM_L_X70Y106_SLICE_X105Y106_CO5),
.O6(CLBLM_L_X70Y106_SLICE_X105Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccff00ec4cff00)
  ) CLBLM_L_X70Y106_SLICE_X105Y106_BLUT (
.I0(CLBLM_L_X68Y108_SLICE_X103Y108_CO6),
.I1(CLBLM_L_X70Y106_SLICE_X105Y106_BQ),
.I2(CLBLM_L_X68Y109_SLICE_X103Y109_B5Q),
.I3(CLBLM_L_X68Y108_SLICE_X103Y108_BQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X68Y109_SLICE_X103Y109_BQ),
.O5(CLBLM_L_X70Y106_SLICE_X105Y106_BO5),
.O6(CLBLM_L_X70Y106_SLICE_X105Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaeffaa00a200)
  ) CLBLM_L_X70Y106_SLICE_X105Y106_ALUT (
.I0(CLBLM_L_X70Y106_SLICE_X105Y106_AQ),
.I1(CLBLM_L_X68Y108_SLICE_X103Y108_CO6),
.I2(CLBLM_L_X68Y109_SLICE_X103Y109_B5Q),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X68Y109_SLICE_X103Y109_BQ),
.I5(CLBLM_L_X70Y107_SLICE_X105Y107_BQ),
.O5(CLBLM_L_X70Y106_SLICE_X105Y106_AO5),
.O6(CLBLM_L_X70Y106_SLICE_X105Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y107_SLICE_X104Y107_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y107_SLICE_X104Y107_AO6),
.Q(CLBLM_L_X70Y107_SLICE_X104Y107_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y107_SLICE_X104Y107_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y107_SLICE_X104Y107_BO6),
.Q(CLBLM_L_X70Y107_SLICE_X104Y107_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y107_SLICE_X104Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y107_SLICE_X104Y107_DO5),
.O6(CLBLM_L_X70Y107_SLICE_X104Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff3f03300)
  ) CLBLM_L_X70Y107_SLICE_X104Y107_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X70Y107_SLICE_X105Y107_AQ),
.I2(CLBLM_L_X70Y106_SLICE_X105Y106_A5Q),
.I3(CLBLM_L_X70Y106_SLICE_X104Y106_A5Q),
.I4(CLBLM_L_X68Y109_SLICE_X103Y109_AQ),
.I5(CLBLM_L_X70Y105_SLICE_X104Y105_CO6),
.O5(CLBLM_L_X70Y107_SLICE_X104Y107_CO5),
.O6(CLBLM_L_X70Y107_SLICE_X104Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcfcfc30303074)
  ) CLBLM_L_X70Y107_SLICE_X104Y107_BLUT (
.I0(CLBLM_L_X68Y107_SLICE_X103Y107_DO6),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_L_X70Y107_SLICE_X104Y107_AQ),
.I3(CLBLM_L_X70Y106_SLICE_X104Y106_DO6),
.I4(CLBLM_L_X70Y106_SLICE_X104Y106_BQ),
.I5(CLBLM_L_X70Y107_SLICE_X104Y107_CO6),
.O5(CLBLM_L_X70Y107_SLICE_X104Y107_BO5),
.O6(CLBLM_L_X70Y107_SLICE_X104Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00000044)
  ) CLBLM_L_X70Y107_SLICE_X104Y107_ALUT (
.I0(CLBLM_L_X68Y107_SLICE_X103Y107_DO6),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(1'b1),
.I3(CLBLM_L_X70Y106_SLICE_X104Y106_DO6),
.I4(CLBLM_L_X70Y106_SLICE_X104Y106_BQ),
.I5(CLBLM_L_X70Y107_SLICE_X104Y107_CO6),
.O5(CLBLM_L_X70Y107_SLICE_X104Y107_AO5),
.O6(CLBLM_L_X70Y107_SLICE_X104Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y107_SLICE_X105Y107_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y107_SLICE_X105Y107_AO6),
.Q(CLBLM_L_X70Y107_SLICE_X105Y107_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y107_SLICE_X105Y107_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y107_SLICE_X105Y107_BO6),
.Q(CLBLM_L_X70Y107_SLICE_X105Y107_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y107_SLICE_X105Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y107_SLICE_X105Y107_DO5),
.O6(CLBLM_L_X70Y107_SLICE_X105Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y107_SLICE_X105Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y107_SLICE_X105Y107_CO5),
.O6(CLBLM_L_X70Y107_SLICE_X105Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000a0a02000a0a0)
  ) CLBLM_L_X70Y107_SLICE_X105Y107_BLUT (
.I0(CLBLL_R_X71Y107_SLICE_X106Y107_DO6),
.I1(CLBLM_L_X68Y109_SLICE_X103Y109_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X68Y108_SLICE_X103Y108_CO6),
.I4(CLBLM_L_X70Y106_SLICE_X105Y106_CO6),
.I5(CLBLM_L_X68Y109_SLICE_X103Y109_B5Q),
.O5(CLBLM_L_X70Y107_SLICE_X105Y107_BO5),
.O6(CLBLM_L_X70Y107_SLICE_X105Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbfbbbfb88c888c8)
  ) CLBLM_L_X70Y107_SLICE_X105Y107_ALUT (
.I0(CLBLM_L_X72Y106_SLICE_X108Y106_CO6),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_L_X70Y107_SLICE_X105Y107_AQ),
.I3(CLBLM_L_X70Y106_SLICE_X105Y106_CO6),
.I4(1'b1),
.I5(CLBLM_L_X72Y108_SLICE_X108Y108_DQ),
.O5(CLBLM_L_X70Y107_SLICE_X105Y107_AO5),
.O6(CLBLM_L_X70Y107_SLICE_X105Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y108_SLICE_X104Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y108_SLICE_X104Y108_DO5),
.O6(CLBLM_L_X70Y108_SLICE_X104Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y108_SLICE_X104Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y108_SLICE_X104Y108_CO5),
.O6(CLBLM_L_X70Y108_SLICE_X104Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y108_SLICE_X104Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y108_SLICE_X104Y108_BO5),
.O6(CLBLM_L_X70Y108_SLICE_X104Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y108_SLICE_X104Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y108_SLICE_X104Y108_AO5),
.O6(CLBLM_L_X70Y108_SLICE_X104Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y108_SLICE_X105Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y108_SLICE_X105Y108_DO5),
.O6(CLBLM_L_X70Y108_SLICE_X105Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y108_SLICE_X105Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y108_SLICE_X105Y108_CO5),
.O6(CLBLM_L_X70Y108_SLICE_X105Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y108_SLICE_X105Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y108_SLICE_X105Y108_BO5),
.O6(CLBLM_L_X70Y108_SLICE_X105Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f3facacacac)
  ) CLBLM_L_X70Y108_SLICE_X105Y108_ALUT (
.I0(CLBLL_R_X71Y108_SLICE_X107Y108_A5Q),
.I1(CLBLM_L_X72Y118_SLICE_X109Y118_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_R_X65Y106_SLICE_X98Y106_CQ),
.I4(CLBLM_L_X74Y109_SLICE_X113Y109_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X70Y108_SLICE_X105Y108_AO5),
.O6(CLBLM_L_X70Y108_SLICE_X105Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y109_SLICE_X104Y109_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y109_SLICE_X104Y109_AO5),
.Q(CLBLM_L_X70Y109_SLICE_X104Y109_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y109_SLICE_X104Y109_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y109_SLICE_X104Y109_BO5),
.Q(CLBLM_L_X70Y109_SLICE_X104Y109_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y109_SLICE_X104Y109_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y109_SLICE_X104Y109_AO6),
.Q(CLBLM_L_X70Y109_SLICE_X104Y109_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y109_SLICE_X104Y109_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y109_SLICE_X104Y109_BO6),
.Q(CLBLM_L_X70Y109_SLICE_X104Y109_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y109_SLICE_X104Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y109_SLICE_X104Y109_DO5),
.O6(CLBLM_L_X70Y109_SLICE_X104Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y109_SLICE_X104Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y109_SLICE_X104Y109_CO5),
.O6(CLBLM_L_X70Y109_SLICE_X104Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaf0faf0eecc44cc)
  ) CLBLM_L_X70Y109_SLICE_X104Y109_BLUT (
.I0(CLBLM_L_X70Y112_SLICE_X105Y112_B5Q),
.I1(CLBLM_L_X70Y109_SLICE_X104Y109_A5Q),
.I2(CLBLM_L_X70Y109_SLICE_X104Y109_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_R_X65Y106_SLICE_X99Y106_AQ),
.I5(1'b1),
.O5(CLBLM_L_X70Y109_SLICE_X104Y109_BO5),
.O6(CLBLM_L_X70Y109_SLICE_X104Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafaf0f0ee44cccc)
  ) CLBLM_L_X70Y109_SLICE_X104Y109_ALUT (
.I0(CLBLM_L_X70Y112_SLICE_X105Y112_B5Q),
.I1(CLBLM_L_X70Y109_SLICE_X104Y109_BQ),
.I2(CLBLM_L_X70Y113_SLICE_X104Y113_B5Q),
.I3(CLBLM_L_X70Y107_SLICE_X104Y107_BQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLM_L_X70Y109_SLICE_X104Y109_AO5),
.O6(CLBLM_L_X70Y109_SLICE_X104Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y109_SLICE_X105Y109_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y109_SLICE_X104Y109_B5Q),
.Q(CLBLM_L_X70Y109_SLICE_X105Y109_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y109_SLICE_X105Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y109_SLICE_X105Y109_DO5),
.O6(CLBLM_L_X70Y109_SLICE_X105Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y109_SLICE_X105Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y109_SLICE_X105Y109_CO5),
.O6(CLBLM_L_X70Y109_SLICE_X105Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y109_SLICE_X105Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y109_SLICE_X105Y109_BO5),
.O6(CLBLM_L_X70Y109_SLICE_X105Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y109_SLICE_X105Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y109_SLICE_X105Y109_AO5),
.O6(CLBLM_L_X70Y109_SLICE_X105Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y110_SLICE_X104Y110_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y110_SLICE_X104Y110_BO5),
.Q(CLBLM_L_X70Y110_SLICE_X104Y110_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y110_SLICE_X104Y110_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y110_SLICE_X104Y110_AO6),
.Q(CLBLM_L_X70Y110_SLICE_X104Y110_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y110_SLICE_X104Y110_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y110_SLICE_X104Y110_BO6),
.Q(CLBLM_L_X70Y110_SLICE_X104Y110_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y110_SLICE_X104Y110_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y110_SLICE_X104Y110_CO6),
.Q(CLBLM_L_X70Y110_SLICE_X104Y110_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y110_SLICE_X104Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y110_SLICE_X104Y110_DO5),
.O6(CLBLM_L_X70Y110_SLICE_X104Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5050505050505072)
  ) CLBLM_L_X70Y110_SLICE_X104Y110_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X70Y110_SLICE_X104Y110_AQ),
.I2(CLBLM_L_X70Y112_SLICE_X104Y112_A5Q),
.I3(CLBLM_L_X70Y110_SLICE_X104Y110_BQ),
.I4(CLBLM_L_X70Y110_SLICE_X104Y110_B5Q),
.I5(CLBLL_R_X71Y111_SLICE_X107Y111_BO6),
.O5(CLBLM_L_X70Y110_SLICE_X104Y110_CO5),
.O6(CLBLM_L_X70Y110_SLICE_X104Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc34f0f0aa62cccc)
  ) CLBLM_L_X70Y110_SLICE_X104Y110_BLUT (
.I0(CLBLM_L_X70Y110_SLICE_X104Y110_B5Q),
.I1(CLBLM_L_X70Y110_SLICE_X104Y110_BQ),
.I2(CLBLM_L_X70Y110_SLICE_X104Y110_AQ),
.I3(CLBLM_L_X70Y111_SLICE_X104Y111_CO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLM_L_X70Y110_SLICE_X104Y110_BO5),
.O6(CLBLM_L_X70Y110_SLICE_X104Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000070001000100)
  ) CLBLM_L_X70Y110_SLICE_X104Y110_ALUT (
.I0(CLBLM_L_X70Y110_SLICE_X104Y110_B5Q),
.I1(CLBLM_L_X70Y110_SLICE_X104Y110_BQ),
.I2(CLBLM_L_X70Y110_SLICE_X104Y110_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X70Y111_SLICE_X104Y111_CO6),
.I5(1'b1),
.O5(CLBLM_L_X70Y110_SLICE_X104Y110_AO5),
.O6(CLBLM_L_X70Y110_SLICE_X104Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y110_SLICE_X105Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y110_SLICE_X105Y110_DO5),
.O6(CLBLM_L_X70Y110_SLICE_X105Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y110_SLICE_X105Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y110_SLICE_X105Y110_CO5),
.O6(CLBLM_L_X70Y110_SLICE_X105Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y110_SLICE_X105Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y110_SLICE_X105Y110_BO5),
.O6(CLBLM_L_X70Y110_SLICE_X105Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y110_SLICE_X105Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y110_SLICE_X105Y110_AO5),
.O6(CLBLM_L_X70Y110_SLICE_X105Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y111_SLICE_X104Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y111_SLICE_X104Y111_BO6),
.Q(CLBLM_L_X70Y111_SLICE_X104Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y111_SLICE_X104Y111_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y111_SLICE_X104Y111_AO5),
.Q(CLBLM_L_X70Y111_SLICE_X104Y111_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000023213331)
  ) CLBLM_L_X70Y111_SLICE_X104Y111_DLUT (
.I0(CLBLM_L_X70Y110_SLICE_X104Y110_BQ),
.I1(CLBLL_R_X71Y111_SLICE_X107Y111_AQ),
.I2(CLBLM_L_X70Y110_SLICE_X104Y110_B5Q),
.I3(CLBLM_L_X72Y111_SLICE_X108Y111_BQ),
.I4(CLBLM_L_X70Y110_SLICE_X104Y110_AQ),
.I5(CLBLM_L_X70Y112_SLICE_X104Y112_AQ),
.O5(CLBLM_L_X70Y111_SLICE_X104Y111_DO5),
.O6(CLBLM_L_X70Y111_SLICE_X104Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfffffffffffffff)
  ) CLBLM_L_X70Y111_SLICE_X104Y111_CLUT (
.I0(CLBLM_L_X70Y111_SLICE_X104Y111_BQ),
.I1(CLBLL_R_X71Y111_SLICE_X107Y111_AQ),
.I2(CLBLM_L_X72Y111_SLICE_X109Y111_A5Q),
.I3(CLBLM_L_X70Y112_SLICE_X104Y112_A5Q),
.I4(CLBLM_L_X72Y111_SLICE_X109Y111_AQ),
.I5(CLBLM_L_X70Y112_SLICE_X104Y112_AQ),
.O5(CLBLM_L_X70Y111_SLICE_X104Y111_CO5),
.O6(CLBLM_L_X70Y111_SLICE_X104Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a07da00000c000)
  ) CLBLM_L_X70Y111_SLICE_X104Y111_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X70Y110_SLICE_X104Y110_BQ),
.I2(CLBLM_L_X70Y111_SLICE_X104Y111_AQ),
.I3(CLBLM_L_X70Y110_SLICE_X104Y110_B5Q),
.I4(CLBLM_L_X70Y111_SLICE_X104Y111_CO6),
.I5(1'b1),
.O5(CLBLM_L_X70Y111_SLICE_X104Y111_BO5),
.O6(CLBLM_L_X70Y111_SLICE_X104Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff7777000000f0)
  ) CLBLM_L_X70Y111_SLICE_X104Y111_ALUT (
.I0(CLBLM_L_X72Y111_SLICE_X109Y111_A5Q),
.I1(CLBLM_L_X72Y111_SLICE_X109Y111_AQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X72Y111_SLICE_X109Y111_CQ),
.I4(CLBLM_L_X70Y111_SLICE_X104Y111_BQ),
.I5(1'b1),
.O5(CLBLM_L_X70Y111_SLICE_X104Y111_AO5),
.O6(CLBLM_L_X70Y111_SLICE_X104Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y111_SLICE_X105Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y111_SLICE_X105Y111_AO6),
.Q(CLBLM_L_X70Y111_SLICE_X105Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y111_SLICE_X105Y111_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y111_SLICE_X105Y111_BO6),
.Q(CLBLM_L_X70Y111_SLICE_X105Y111_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaaaaaa8a8)
  ) CLBLM_L_X70Y111_SLICE_X105Y111_DLUT (
.I0(CLBLM_L_X70Y112_SLICE_X105Y112_AQ),
.I1(CLBLM_L_X70Y110_SLICE_X104Y110_B5Q),
.I2(CLBLL_R_X71Y112_SLICE_X106Y112_AQ),
.I3(1'b1),
.I4(CLBLM_L_X70Y110_SLICE_X104Y110_AQ),
.I5(CLBLM_L_X70Y110_SLICE_X104Y110_BQ),
.O5(CLBLM_L_X70Y111_SLICE_X105Y111_DO5),
.O6(CLBLM_L_X70Y111_SLICE_X105Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2000000000000000)
  ) CLBLM_L_X70Y111_SLICE_X105Y111_CLUT (
.I0(CLBLM_L_X70Y111_SLICE_X104Y111_AQ),
.I1(CLBLM_L_X70Y111_SLICE_X104Y111_CO6),
.I2(CLBLM_L_X70Y110_SLICE_X104Y110_BQ),
.I3(CLBLL_R_X71Y111_SLICE_X106Y111_BQ),
.I4(CLBLM_L_X70Y110_SLICE_X104Y110_B5Q),
.I5(CLBLL_R_X71Y111_SLICE_X106Y111_CQ),
.O5(CLBLM_L_X70Y111_SLICE_X105Y111_CO5),
.O6(CLBLM_L_X70Y111_SLICE_X105Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h30fcf0f000ccf0f0)
  ) CLBLM_L_X70Y111_SLICE_X105Y111_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X70Y111_SLICE_X105Y111_BQ),
.I2(CLBLM_L_X70Y111_SLICE_X105Y111_AQ),
.I3(CLBLM_L_X70Y111_SLICE_X104Y111_BO5),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X70Y111_SLICE_X105Y111_CO6),
.O5(CLBLM_L_X70Y111_SLICE_X105Y111_BO5),
.O6(CLBLM_L_X70Y111_SLICE_X105Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h12f0aaaa30f0aaaa)
  ) CLBLM_L_X70Y111_SLICE_X105Y111_ALUT (
.I0(CLBLL_R_X71Y111_SLICE_X106Y111_CQ),
.I1(CLBLM_L_X70Y111_SLICE_X105Y111_BQ),
.I2(CLBLM_L_X70Y111_SLICE_X105Y111_AQ),
.I3(CLBLM_L_X70Y111_SLICE_X104Y111_BO5),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X71Y111_SLICE_X106Y111_BQ),
.O5(CLBLM_L_X70Y111_SLICE_X105Y111_AO5),
.O6(CLBLM_L_X70Y111_SLICE_X105Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y112_SLICE_X104Y112_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y112_SLICE_X104Y112_BO6),
.Q(CLBLM_L_X70Y112_SLICE_X104Y112_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y112_SLICE_X104Y112_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y112_SLICE_X104Y112_CO5),
.Q(CLBLM_L_X70Y112_SLICE_X104Y112_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y112_SLICE_X104Y112_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y112_SLICE_X104Y112_AO6),
.Q(CLBLM_L_X70Y112_SLICE_X104Y112_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y112_SLICE_X104Y112_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y112_SLICE_X104Y112_CO6),
.Q(CLBLM_L_X70Y112_SLICE_X104Y112_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y112_SLICE_X104Y112_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y112_SLICE_X104Y112_DO6),
.Q(CLBLM_L_X70Y112_SLICE_X104Y112_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5500753055005500)
  ) CLBLM_L_X70Y112_SLICE_X104Y112_DLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X71Y111_SLICE_X107Y111_AQ),
.I2(CLBLM_L_X72Y111_SLICE_X109Y111_CQ),
.I3(CLBLM_L_X70Y110_SLICE_X104Y110_CQ),
.I4(CLBLM_L_X70Y112_SLICE_X104Y112_BO5),
.I5(CLBLM_L_X70Y110_SLICE_X104Y110_AO5),
.O5(CLBLM_L_X70Y112_SLICE_X104Y112_DO5),
.O6(CLBLM_L_X70Y112_SLICE_X104Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5fff0aaaeecceecc)
  ) CLBLM_L_X70Y112_SLICE_X104Y112_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X70Y112_SLICE_X105Y112_C5Q),
.I2(CLBLM_L_X70Y112_SLICE_X104Y112_DQ),
.I3(CLBLM_L_X70Y112_SLICE_X105Y112_B5Q),
.I4(CLBLM_L_X70Y113_SLICE_X104Y113_BQ),
.I5(1'b1),
.O5(CLBLM_L_X70Y112_SLICE_X104Y112_CO5),
.O6(CLBLM_L_X70Y112_SLICE_X104Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdff020f0fffff0f0)
  ) CLBLM_L_X70Y112_SLICE_X104Y112_BLUT (
.I0(CLBLL_R_X71Y111_SLICE_X107Y111_AQ),
.I1(CLBLM_L_X70Y111_SLICE_X104Y111_AO6),
.I2(CLBLM_L_X70Y112_SLICE_X104Y112_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X70Y112_SLICE_X104Y112_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X70Y112_SLICE_X104Y112_BO5),
.O6(CLBLM_L_X70Y112_SLICE_X104Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd2aaf0aaf0aaf0aa)
  ) CLBLM_L_X70Y112_SLICE_X104Y112_ALUT (
.I0(CLBLL_R_X71Y111_SLICE_X107Y111_AQ),
.I1(CLBLM_L_X70Y111_SLICE_X104Y111_BQ),
.I2(CLBLM_L_X70Y112_SLICE_X104Y112_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X72Y111_SLICE_X109Y111_AQ),
.I5(CLBLM_L_X72Y111_SLICE_X109Y111_A5Q),
.O5(CLBLM_L_X70Y112_SLICE_X104Y112_AO5),
.O6(CLBLM_L_X70Y112_SLICE_X104Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y112_SLICE_X105Y112_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y112_SLICE_X105Y112_AO5),
.Q(CLBLM_L_X70Y112_SLICE_X105Y112_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y112_SLICE_X105Y112_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y112_SLICE_X105Y112_BO5),
.Q(CLBLM_L_X70Y112_SLICE_X105Y112_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y112_SLICE_X105Y112_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y112_SLICE_X105Y112_CO5),
.Q(CLBLM_L_X70Y112_SLICE_X105Y112_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y112_SLICE_X105Y112_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y112_SLICE_X105Y112_DO5),
.Q(CLBLM_L_X70Y112_SLICE_X105Y112_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y112_SLICE_X105Y112_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y112_SLICE_X105Y112_AO6),
.Q(CLBLM_L_X70Y112_SLICE_X105Y112_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y112_SLICE_X105Y112_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y112_SLICE_X105Y112_BO6),
.Q(CLBLM_L_X70Y112_SLICE_X105Y112_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y112_SLICE_X105Y112_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y112_SLICE_X105Y112_CO6),
.Q(CLBLM_L_X70Y112_SLICE_X105Y112_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y112_SLICE_X105Y112_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y112_SLICE_X105Y112_DO6),
.Q(CLBLM_L_X70Y112_SLICE_X105Y112_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeeccccfafaf0f0)
  ) CLBLM_L_X70Y112_SLICE_X105Y112_DLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X70Y112_SLICE_X105Y112_CQ),
.I2(CLBLM_L_X70Y112_SLICE_X105Y112_DQ),
.I3(1'b1),
.I4(CLBLM_L_X70Y112_SLICE_X105Y112_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X70Y112_SLICE_X105Y112_DO5),
.O6(CLBLM_L_X70Y112_SLICE_X105Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaccaafff0ccf0)
  ) CLBLM_L_X70Y112_SLICE_X105Y112_CLUT (
.I0(CLBLM_L_X68Y112_SLICE_X103Y112_BQ),
.I1(CLBLL_R_X71Y111_SLICE_X106Y111_A5Q),
.I2(CLBLL_R_X71Y108_SLICE_X107Y108_A5Q),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X70Y112_SLICE_X105Y112_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X70Y112_SLICE_X105Y112_CO5),
.O6(CLBLM_L_X70Y112_SLICE_X105Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5050f0f01f1f1010)
  ) CLBLM_L_X70Y112_SLICE_X105Y112_BLUT (
.I0(CLBLL_R_X71Y112_SLICE_X106Y112_B5Q),
.I1(CLBLM_L_X70Y112_SLICE_X105Y112_A5Q),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(1'b1),
.I4(CLBLL_R_X71Y112_SLICE_X106Y112_BQ),
.I5(1'b1),
.O5(CLBLM_L_X70Y112_SLICE_X105Y112_BO5),
.O6(CLBLM_L_X70Y112_SLICE_X105Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee4444d8fad8d8)
  ) CLBLM_L_X70Y112_SLICE_X105Y112_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X70Y112_SLICE_X105Y112_BQ),
.I2(CLBLM_L_X70Y112_SLICE_X105Y112_AQ),
.I3(CLBLL_R_X71Y112_SLICE_X106Y112_BQ),
.I4(CLBLM_L_X70Y112_SLICE_X105Y112_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X70Y112_SLICE_X105Y112_AO5),
.O6(CLBLM_L_X70Y112_SLICE_X105Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y113_SLICE_X104Y113_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y113_SLICE_X104Y113_AO5),
.Q(CLBLM_L_X70Y113_SLICE_X104Y113_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y113_SLICE_X104Y113_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y113_SLICE_X104Y113_BO5),
.Q(CLBLM_L_X70Y113_SLICE_X104Y113_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y113_SLICE_X104Y113_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y113_SLICE_X104Y113_AO6),
.Q(CLBLM_L_X70Y113_SLICE_X104Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y113_SLICE_X104Y113_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y113_SLICE_X104Y113_BO6),
.Q(CLBLM_L_X70Y113_SLICE_X104Y113_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y113_SLICE_X104Y113_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y113_SLICE_X104Y113_CO6),
.Q(CLBLM_L_X70Y113_SLICE_X104Y113_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y113_SLICE_X104Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y113_SLICE_X104Y113_DO5),
.O6(CLBLM_L_X70Y113_SLICE_X104Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hddf5ddf588a088a0)
  ) CLBLM_L_X70Y113_SLICE_X104Y113_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_R_X65Y106_SLICE_X99Y106_DQ),
.I2(CLBLM_L_X70Y113_SLICE_X104Y113_BQ),
.I3(CLBLM_L_X70Y112_SLICE_X105Y112_B5Q),
.I4(1'b1),
.I5(CLBLM_L_X72Y111_SLICE_X108Y111_BQ),
.O5(CLBLM_L_X70Y113_SLICE_X104Y113_CO5),
.O6(CLBLM_L_X70Y113_SLICE_X104Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccccccfff0f0f0)
  ) CLBLM_L_X70Y113_SLICE_X104Y113_BLUT (
.I0(CLBLM_L_X70Y107_SLICE_X104Y107_AQ),
.I1(CLBLM_L_X70Y113_SLICE_X104Y113_A5Q),
.I2(CLBLM_L_X70Y112_SLICE_X104Y112_C5Q),
.I3(CLBLM_L_X70Y112_SLICE_X105Y112_B5Q),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLM_L_X70Y113_SLICE_X104Y113_BO5),
.O6(CLBLM_L_X70Y113_SLICE_X104Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccccccfff0f0f0)
  ) CLBLM_L_X70Y113_SLICE_X104Y113_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X70Y112_SLICE_X105Y112_D5Q),
.I2(CLBLM_L_X70Y113_SLICE_X104Y113_AQ),
.I3(CLBLM_L_X70Y112_SLICE_X105Y112_B5Q),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLM_L_X70Y113_SLICE_X104Y113_AO5),
.O6(CLBLM_L_X70Y113_SLICE_X104Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y113_SLICE_X105Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y113_SLICE_X105Y113_DO5),
.O6(CLBLM_L_X70Y113_SLICE_X105Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y113_SLICE_X105Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y113_SLICE_X105Y113_CO5),
.O6(CLBLM_L_X70Y113_SLICE_X105Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y113_SLICE_X105Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y113_SLICE_X105Y113_BO5),
.O6(CLBLM_L_X70Y113_SLICE_X105Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y113_SLICE_X105Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y113_SLICE_X105Y113_AO5),
.O6(CLBLM_L_X70Y113_SLICE_X105Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y114_SLICE_X104Y114_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y117_SLICE_X106Y117_B5Q),
.Q(CLBLM_L_X70Y114_SLICE_X104Y114_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y114_SLICE_X104Y114_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y114_SLICE_X104Y114_AO6),
.Q(CLBLM_L_X70Y114_SLICE_X104Y114_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y114_SLICE_X104Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y114_SLICE_X104Y114_DO5),
.O6(CLBLM_L_X70Y114_SLICE_X104Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y114_SLICE_X104Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y114_SLICE_X104Y114_CO5),
.O6(CLBLM_L_X70Y114_SLICE_X104Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y114_SLICE_X104Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y114_SLICE_X104Y114_BO5),
.O6(CLBLM_L_X70Y114_SLICE_X104Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f0ffff00fa0000)
  ) CLBLM_L_X70Y114_SLICE_X104Y114_ALUT (
.I0(CLBLL_R_X71Y117_SLICE_X106Y117_B5Q),
.I1(1'b1),
.I2(CLBLM_L_X70Y114_SLICE_X104Y114_AQ),
.I3(CLBLM_L_X68Y109_SLICE_X102Y109_AQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X70Y114_SLICE_X104Y114_A5Q),
.O5(CLBLM_L_X70Y114_SLICE_X104Y114_AO5),
.O6(CLBLM_L_X70Y114_SLICE_X104Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y114_SLICE_X105Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y114_SLICE_X105Y114_DO5),
.O6(CLBLM_L_X70Y114_SLICE_X105Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y114_SLICE_X105Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y114_SLICE_X105Y114_CO5),
.O6(CLBLM_L_X70Y114_SLICE_X105Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y114_SLICE_X105Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y114_SLICE_X105Y114_BO5),
.O6(CLBLM_L_X70Y114_SLICE_X105Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y114_SLICE_X105Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y114_SLICE_X105Y114_AO5),
.O6(CLBLM_L_X70Y114_SLICE_X105Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y119_SLICE_X104Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y119_SLICE_X104Y119_DO5),
.O6(CLBLM_L_X70Y119_SLICE_X104Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y119_SLICE_X104Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y119_SLICE_X104Y119_CO5),
.O6(CLBLM_L_X70Y119_SLICE_X104Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y119_SLICE_X104Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y119_SLICE_X104Y119_BO5),
.O6(CLBLM_L_X70Y119_SLICE_X104Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y119_SLICE_X104Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y119_SLICE_X104Y119_AO5),
.O6(CLBLM_L_X70Y119_SLICE_X104Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y119_SLICE_X105Y119_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y119_SLICE_X105Y119_AO5),
.Q(CLBLM_L_X70Y119_SLICE_X105Y119_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y119_SLICE_X105Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y119_SLICE_X105Y119_AO6),
.Q(CLBLM_L_X70Y119_SLICE_X105Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y119_SLICE_X105Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y119_SLICE_X105Y119_DO5),
.O6(CLBLM_L_X70Y119_SLICE_X105Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y119_SLICE_X105Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y119_SLICE_X105Y119_CO5),
.O6(CLBLM_L_X70Y119_SLICE_X105Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y119_SLICE_X105Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y119_SLICE_X105Y119_BO5),
.O6(CLBLM_L_X70Y119_SLICE_X105Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafafafac0c0c0c0)
  ) CLBLM_L_X70Y119_SLICE_X105Y119_ALUT (
.I0(CLBLM_L_X70Y123_SLICE_X104Y123_A5Q),
.I1(CLBLL_R_X71Y108_SLICE_X107Y108_A5Q),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y119_SLICE_X105Y119_AO5),
.O6(CLBLM_L_X70Y119_SLICE_X105Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y123_SLICE_X104Y123_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y123_SLICE_X104Y123_AO5),
.Q(CLBLM_L_X70Y123_SLICE_X104Y123_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y123_SLICE_X104Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y123_SLICE_X104Y123_AO6),
.Q(CLBLM_L_X70Y123_SLICE_X104Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y123_SLICE_X104Y123_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y123_SLICE_X104Y123_BO6),
.Q(CLBLM_L_X70Y123_SLICE_X104Y123_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y123_SLICE_X104Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y123_SLICE_X104Y123_DO5),
.O6(CLBLM_L_X70Y123_SLICE_X104Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdffffffffffffff)
  ) CLBLM_L_X70Y123_SLICE_X104Y123_CLUT (
.I0(CLBLM_L_X70Y119_SLICE_X105Y119_AQ),
.I1(CLBLM_L_X70Y123_SLICE_X104Y123_AQ),
.I2(CLBLL_R_X71Y126_SLICE_X107Y126_BQ),
.I3(CLBLM_L_X70Y123_SLICE_X104Y123_A5Q),
.I4(CLBLM_L_X70Y123_SLICE_X104Y123_BQ),
.I5(CLBLM_L_X70Y125_SLICE_X104Y125_AQ),
.O5(CLBLM_L_X70Y123_SLICE_X104Y123_CO5),
.O6(CLBLM_L_X70Y123_SLICE_X104Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafafafafafafafa)
  ) CLBLM_L_X70Y123_SLICE_X104Y123_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(1'b1),
.I2(CLBLM_L_X70Y123_SLICE_X104Y123_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y123_SLICE_X104Y123_BO5),
.O6(CLBLM_L_X70Y123_SLICE_X104Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaffaa50505050)
  ) CLBLM_L_X70Y123_SLICE_X104Y123_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(1'b1),
.I2(CLBLM_L_X70Y125_SLICE_X104Y125_AQ),
.I3(CLBLL_R_X71Y126_SLICE_X107Y126_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y123_SLICE_X104Y123_AO5),
.O6(CLBLM_L_X70Y123_SLICE_X104Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y123_SLICE_X105Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y123_SLICE_X105Y123_DO5),
.O6(CLBLM_L_X70Y123_SLICE_X105Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y123_SLICE_X105Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y123_SLICE_X105Y123_CO5),
.O6(CLBLM_L_X70Y123_SLICE_X105Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y123_SLICE_X105Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y123_SLICE_X105Y123_BO5),
.O6(CLBLM_L_X70Y123_SLICE_X105Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y123_SLICE_X105Y123_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y123_SLICE_X105Y123_AO5),
.O6(CLBLM_L_X70Y123_SLICE_X105Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y124_SLICE_X104Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y124_SLICE_X104Y124_AO6),
.Q(CLBLM_L_X70Y124_SLICE_X104Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y124_SLICE_X104Y124_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y124_SLICE_X104Y124_BO6),
.Q(CLBLM_L_X70Y124_SLICE_X104Y124_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y124_SLICE_X104Y124_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y124_SLICE_X104Y124_CO6),
.Q(CLBLM_L_X70Y124_SLICE_X104Y124_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7ffffffffffffff)
  ) CLBLM_L_X70Y124_SLICE_X104Y124_DLUT (
.I0(CLBLM_L_X70Y119_SLICE_X105Y119_AQ),
.I1(CLBLM_L_X70Y123_SLICE_X104Y123_A5Q),
.I2(CLBLM_L_X70Y123_SLICE_X104Y123_AQ),
.I3(CLBLM_L_X70Y125_SLICE_X104Y125_AQ),
.I4(CLBLM_L_X70Y123_SLICE_X104Y123_BQ),
.I5(CLBLL_R_X71Y126_SLICE_X107Y126_BQ),
.O5(CLBLM_L_X70Y124_SLICE_X104Y124_DO5),
.O6(CLBLM_L_X70Y124_SLICE_X104Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdcdc5050dcff5050)
  ) CLBLM_L_X70Y124_SLICE_X104Y124_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X70Y124_SLICE_X104Y124_CQ),
.I2(CLBLM_L_X70Y124_SLICE_X104Y124_AQ),
.I3(CLBLM_L_X72Y122_SLICE_X109Y122_BQ),
.I4(CLBLM_L_X70Y125_SLICE_X105Y125_AO5),
.I5(CLBLM_L_X70Y125_SLICE_X105Y125_BO6),
.O5(CLBLM_L_X70Y124_SLICE_X104Y124_CO5),
.O6(CLBLM_L_X70Y124_SLICE_X104Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8dff8dff8d008d00)
  ) CLBLM_L_X70Y124_SLICE_X104Y124_BLUT (
.I0(CLBLM_L_X70Y123_SLICE_X104Y123_CO6),
.I1(CLBLM_L_X70Y124_SLICE_X104Y124_BQ),
.I2(CLBLM_L_X70Y124_SLICE_X104Y124_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(1'b1),
.I5(CLBLM_L_X70Y126_SLICE_X104Y126_CQ),
.O5(CLBLM_L_X70Y124_SLICE_X104Y124_BO5),
.O6(CLBLM_L_X70Y124_SLICE_X104Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a2a2ffa0ffa2)
  ) CLBLM_L_X70Y124_SLICE_X104Y124_ALUT (
.I0(CLBLM_L_X70Y125_SLICE_X105Y125_AO5),
.I1(CLBLM_L_X70Y125_SLICE_X105Y125_BO6),
.I2(CLBLM_L_X70Y124_SLICE_X104Y124_AQ),
.I3(CLBLL_R_X71Y124_SLICE_X106Y124_AQ),
.I4(CLBLL_R_X73Y124_SLICE_X110Y124_AQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X70Y124_SLICE_X104Y124_AO5),
.O6(CLBLM_L_X70Y124_SLICE_X104Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_L_X70Y124_SLICE_X105Y124_DLUT (
.I0(CLBLM_L_X70Y119_SLICE_X105Y119_AQ),
.I1(CLBLM_L_X70Y125_SLICE_X104Y125_AQ),
.I2(CLBLM_L_X70Y123_SLICE_X104Y123_BQ),
.I3(CLBLM_L_X70Y123_SLICE_X104Y123_A5Q),
.I4(CLBLM_L_X70Y123_SLICE_X104Y123_AQ),
.I5(CLBLL_R_X71Y126_SLICE_X107Y126_BQ),
.O5(CLBLM_L_X70Y124_SLICE_X105Y124_DO5),
.O6(CLBLM_L_X70Y124_SLICE_X105Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff7fffffff)
  ) CLBLM_L_X70Y124_SLICE_X105Y124_CLUT (
.I0(CLBLM_L_X70Y119_SLICE_X105Y119_AQ),
.I1(CLBLM_L_X70Y125_SLICE_X104Y125_AQ),
.I2(CLBLM_L_X70Y123_SLICE_X104Y123_BQ),
.I3(CLBLM_L_X70Y123_SLICE_X104Y123_A5Q),
.I4(CLBLM_L_X70Y123_SLICE_X104Y123_AQ),
.I5(CLBLL_R_X71Y126_SLICE_X107Y126_BQ),
.O5(CLBLM_L_X70Y124_SLICE_X105Y124_CO5),
.O6(CLBLM_L_X70Y124_SLICE_X105Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0055005500550051)
  ) CLBLM_L_X70Y124_SLICE_X105Y124_BLUT (
.I0(CLBLM_L_X70Y123_SLICE_X104Y123_AQ),
.I1(CLBLM_L_X70Y123_SLICE_X104Y123_BQ),
.I2(CLBLM_L_X70Y119_SLICE_X105Y119_AQ),
.I3(CLBLL_R_X71Y126_SLICE_X107Y126_BQ),
.I4(CLBLM_L_X70Y125_SLICE_X104Y125_AQ),
.I5(CLBLM_L_X70Y123_SLICE_X104Y123_A5Q),
.O5(CLBLM_L_X70Y124_SLICE_X105Y124_BO5),
.O6(CLBLM_L_X70Y124_SLICE_X105Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000e0000000f)
  ) CLBLM_L_X70Y124_SLICE_X105Y124_ALUT (
.I0(CLBLM_L_X70Y123_SLICE_X104Y123_AQ),
.I1(CLBLL_R_X71Y126_SLICE_X107Y126_BQ),
.I2(CLBLL_R_X71Y126_SLICE_X107Y126_AQ),
.I3(CLBLM_L_X70Y124_SLICE_X105Y124_BO6),
.I4(CLBLM_L_X70Y125_SLICE_X105Y125_AQ),
.I5(CLBLM_L_X70Y125_SLICE_X104Y125_BQ),
.O5(CLBLM_L_X70Y124_SLICE_X105Y124_AO5),
.O6(CLBLM_L_X70Y124_SLICE_X105Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y125_SLICE_X104Y125_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y125_SLICE_X104Y125_AO5),
.Q(CLBLM_L_X70Y125_SLICE_X104Y125_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y125_SLICE_X104Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y125_SLICE_X104Y125_AO6),
.Q(CLBLM_L_X70Y125_SLICE_X104Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y125_SLICE_X104Y125_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y125_SLICE_X104Y125_BO6),
.Q(CLBLM_L_X70Y125_SLICE_X104Y125_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y125_SLICE_X104Y125_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y125_SLICE_X104Y125_CO6),
.Q(CLBLM_L_X70Y125_SLICE_X104Y125_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0207a2a75257f2f7)
  ) CLBLM_L_X70Y125_SLICE_X104Y125_DLUT (
.I0(CLBLL_R_X71Y126_SLICE_X107Y126_BQ),
.I1(CLBLM_L_X70Y125_SLICE_X104Y125_CQ),
.I2(CLBLM_L_X70Y123_SLICE_X104Y123_AQ),
.I3(CLBLM_L_X70Y125_SLICE_X104Y125_BQ),
.I4(CLBLL_R_X71Y125_SLICE_X107Y125_AQ),
.I5(CLBLL_R_X71Y125_SLICE_X106Y125_AQ),
.O5(CLBLM_L_X70Y125_SLICE_X104Y125_DO5),
.O6(CLBLM_L_X70Y125_SLICE_X104Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0cfffffc0cf0000)
  ) CLBLM_L_X70Y125_SLICE_X104Y125_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X70Y125_SLICE_X104Y125_CQ),
.I2(CLBLM_L_X70Y124_SLICE_X104Y124_DO6),
.I3(CLBLM_L_X70Y126_SLICE_X104Y126_BQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X71Y125_SLICE_X106Y125_AQ),
.O5(CLBLM_L_X70Y125_SLICE_X104Y125_CO5),
.O6(CLBLM_L_X70Y125_SLICE_X104Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22eeee222222ee)
  ) CLBLM_L_X70Y125_SLICE_X104Y125_BLUT (
.I0(CLBLM_L_X70Y125_SLICE_X104Y125_CQ),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(1'b1),
.I3(CLBLM_L_X70Y123_SLICE_X104Y123_CO6),
.I4(CLBLM_L_X70Y126_SLICE_X104Y126_AQ),
.I5(CLBLM_L_X70Y125_SLICE_X104Y125_BQ),
.O5(CLBLM_L_X70Y125_SLICE_X104Y125_BO5),
.O6(CLBLM_L_X70Y125_SLICE_X104Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33330000ffccffcc)
  ) CLBLM_L_X70Y125_SLICE_X104Y125_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(1'b1),
.I3(CLBLM_L_X70Y125_SLICE_X105Y125_BQ),
.I4(CLBLM_L_X70Y123_SLICE_X104Y123_BQ),
.I5(1'b1),
.O5(CLBLM_L_X70Y125_SLICE_X104Y125_AO5),
.O6(CLBLM_L_X70Y125_SLICE_X104Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y125_SLICE_X105Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(RIOB33_X105Y51_IOB_X1Y51_I),
.Q(CLBLM_L_X70Y125_SLICE_X105Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y125_SLICE_X105Y125_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y125_SLICE_X105Y125_AO6),
.Q(CLBLM_L_X70Y125_SLICE_X105Y125_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd5d5ddddd5d55555)
  ) CLBLM_L_X70Y125_SLICE_X105Y125_DLUT (
.I0(CLBLM_L_X70Y124_SLICE_X105Y124_DO6),
.I1(CLBLL_R_X71Y126_SLICE_X107Y126_AQ),
.I2(CLBLL_R_X71Y125_SLICE_X107Y125_AQ),
.I3(1'b1),
.I4(CLBLM_L_X70Y125_SLICE_X105Y125_AQ),
.I5(CLBLL_R_X71Y125_SLICE_X106Y125_AQ),
.O5(CLBLM_L_X70Y125_SLICE_X105Y125_DO5),
.O6(CLBLM_L_X70Y125_SLICE_X105Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fcfef0f0fdff)
  ) CLBLM_L_X70Y125_SLICE_X105Y125_CLUT (
.I0(CLBLM_L_X70Y125_SLICE_X105Y125_AQ),
.I1(CLBLL_R_X71Y126_SLICE_X107Y126_AQ),
.I2(CLBLM_L_X70Y126_SLICE_X105Y126_DO6),
.I3(CLBLM_L_X70Y125_SLICE_X104Y125_CQ),
.I4(CLBLM_L_X70Y125_SLICE_X105Y125_DO6),
.I5(CLBLM_L_X70Y125_SLICE_X104Y125_BQ),
.O5(CLBLM_L_X70Y125_SLICE_X105Y125_CO5),
.O6(CLBLM_L_X70Y125_SLICE_X105Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc00f000f3fffffff)
  ) CLBLM_L_X70Y125_SLICE_X105Y125_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X70Y123_SLICE_X104Y123_BQ),
.I2(CLBLM_L_X70Y119_SLICE_X105Y119_AQ),
.I3(CLBLM_L_X70Y123_SLICE_X104Y123_A5Q),
.I4(CLBLM_L_X70Y125_SLICE_X104Y125_AQ),
.I5(1'b1),
.O5(CLBLM_L_X70Y125_SLICE_X105Y125_BO5),
.O6(CLBLM_L_X70Y125_SLICE_X105Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0fff0fc00ff00)
  ) CLBLM_L_X70Y125_SLICE_X105Y125_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X70Y123_SLICE_X104Y123_A5Q),
.I2(CLBLM_L_X70Y119_SLICE_X105Y119_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X70Y125_SLICE_X104Y125_AQ),
.I5(1'b1),
.O5(CLBLM_L_X70Y125_SLICE_X105Y125_AO5),
.O6(CLBLM_L_X70Y125_SLICE_X105Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y126_SLICE_X104Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y126_SLICE_X104Y126_AO6),
.Q(CLBLM_L_X70Y126_SLICE_X104Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y126_SLICE_X104Y126_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y126_SLICE_X104Y126_BO6),
.Q(CLBLM_L_X70Y126_SLICE_X104Y126_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y126_SLICE_X104Y126_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y126_SLICE_X104Y126_CO6),
.Q(CLBLM_L_X70Y126_SLICE_X104Y126_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0033ff33550f550f)
  ) CLBLM_L_X70Y126_SLICE_X104Y126_DLUT (
.I0(CLBLM_L_X70Y126_SLICE_X105Y126_AQ),
.I1(CLBLM_L_X70Y126_SLICE_X104Y126_CQ),
.I2(CLBLM_L_X70Y124_SLICE_X104Y124_BQ),
.I3(CLBLM_L_X70Y123_SLICE_X104Y123_AQ),
.I4(CLBLL_R_X71Y126_SLICE_X106Y126_AQ),
.I5(CLBLL_R_X71Y126_SLICE_X107Y126_BQ),
.O5(CLBLM_L_X70Y126_SLICE_X104Y126_DO5),
.O6(CLBLM_L_X70Y126_SLICE_X104Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcaca0afacaca0afa)
  ) CLBLM_L_X70Y126_SLICE_X104Y126_CLUT (
.I0(CLBLM_L_X70Y126_SLICE_X105Y126_AQ),
.I1(CLBLM_L_X70Y126_SLICE_X104Y126_CQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X70Y124_SLICE_X104Y124_CQ),
.I4(CLBLM_L_X70Y124_SLICE_X104Y124_DO6),
.I5(1'b1),
.O5(CLBLM_L_X70Y126_SLICE_X104Y126_CO5),
.O6(CLBLM_L_X70Y126_SLICE_X104Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd5c0d5c0d5c0f5f0)
  ) CLBLM_L_X70Y126_SLICE_X104Y126_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X70Y126_SLICE_X104Y126_BQ),
.I2(CLBLM_L_X70Y125_SLICE_X105Y125_AO5),
.I3(CLBLM_L_X70Y126_SLICE_X104Y126_AQ),
.I4(CLBLM_L_X70Y125_SLICE_X105Y125_BO6),
.I5(CLBLM_L_X70Y129_SLICE_X104Y129_BQ),
.O5(CLBLM_L_X70Y126_SLICE_X104Y126_BO5),
.O6(CLBLM_L_X70Y126_SLICE_X104Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd5d5d5ddc0c0c0cc)
  ) CLBLM_L_X70Y126_SLICE_X104Y126_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X70Y125_SLICE_X105Y125_AO5),
.I2(CLBLM_L_X70Y126_SLICE_X104Y126_AQ),
.I3(CLBLM_L_X70Y133_SLICE_X104Y133_BQ),
.I4(CLBLM_L_X70Y125_SLICE_X105Y125_BO6),
.I5(CLBLM_L_X70Y125_SLICE_X104Y125_A5Q),
.O5(CLBLM_L_X70Y126_SLICE_X104Y126_AO5),
.O6(CLBLM_L_X70Y126_SLICE_X104Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y126_SLICE_X105Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y126_SLICE_X105Y126_AO6),
.Q(CLBLM_L_X70Y126_SLICE_X105Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y126_SLICE_X105Y126_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y126_SLICE_X105Y126_BO6),
.Q(CLBLM_L_X70Y126_SLICE_X105Y126_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000ef000000ea)
  ) CLBLM_L_X70Y126_SLICE_X105Y126_DLUT (
.I0(CLBLL_R_X71Y126_SLICE_X107Y126_AQ),
.I1(CLBLM_L_X70Y128_SLICE_X104Y128_CQ),
.I2(CLBLM_L_X70Y125_SLICE_X105Y125_AQ),
.I3(CLBLL_R_X71Y126_SLICE_X107Y126_AO5),
.I4(CLBLM_L_X70Y124_SLICE_X105Y124_DO6),
.I5(CLBLM_L_X70Y133_SLICE_X105Y133_BQ),
.O5(CLBLM_L_X70Y126_SLICE_X105Y126_DO5),
.O6(CLBLM_L_X70Y126_SLICE_X105Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000f0d0000)
  ) CLBLM_L_X70Y126_SLICE_X105Y126_CLUT (
.I0(CLBLM_L_X70Y125_SLICE_X104Y125_CQ),
.I1(CLBLM_L_X70Y123_SLICE_X104Y123_AQ),
.I2(CLBLL_R_X71Y126_SLICE_X107Y126_AQ),
.I3(CLBLL_R_X71Y126_SLICE_X107Y126_BQ),
.I4(CLBLM_L_X70Y125_SLICE_X105Y125_AQ),
.I5(CLBLM_L_X70Y124_SLICE_X105Y124_BO6),
.O5(CLBLM_L_X70Y126_SLICE_X105Y126_CO5),
.O6(CLBLM_L_X70Y126_SLICE_X105Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddf5555cccf0000)
  ) CLBLM_L_X70Y126_SLICE_X105Y126_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X70Y126_SLICE_X105Y126_BQ),
.I2(CLBLM_L_X70Y125_SLICE_X105Y125_BO6),
.I3(CLBLL_R_X73Y126_SLICE_X110Y126_BQ),
.I4(CLBLM_L_X70Y125_SLICE_X105Y125_AO5),
.I5(CLBLM_L_X70Y124_SLICE_X104Y124_CQ),
.O5(CLBLM_L_X70Y126_SLICE_X105Y126_BO5),
.O6(CLBLM_L_X70Y126_SLICE_X105Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a077227722)
  ) CLBLM_L_X70Y126_SLICE_X105Y126_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X70Y126_SLICE_X105Y126_BQ),
.I2(CLBLM_L_X70Y126_SLICE_X105Y126_AQ),
.I3(CLBLL_R_X71Y126_SLICE_X106Y126_AQ),
.I4(1'b1),
.I5(CLBLM_L_X70Y124_SLICE_X105Y124_CO6),
.O5(CLBLM_L_X70Y126_SLICE_X105Y126_AO5),
.O6(CLBLM_L_X70Y126_SLICE_X105Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y128_SLICE_X104Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y128_SLICE_X104Y128_BO6),
.Q(CLBLM_L_X70Y128_SLICE_X104Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y128_SLICE_X104Y128_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y128_SLICE_X104Y128_AO5),
.Q(CLBLM_L_X70Y128_SLICE_X104Y128_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y128_SLICE_X104Y128_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y128_SLICE_X104Y128_CO6),
.Q(CLBLM_L_X70Y128_SLICE_X104Y128_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y128_SLICE_X104Y128_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y128_SLICE_X104Y128_DO6),
.Q(CLBLM_L_X70Y128_SLICE_X104Y128_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c3cccccf0f0cccc)
  ) CLBLM_L_X70Y128_SLICE_X104Y128_DLUT (
.I0(CLBLM_L_X70Y129_SLICE_X104Y129_AQ),
.I1(CLBLM_L_X70Y128_SLICE_X104Y128_CQ),
.I2(CLBLM_L_X70Y128_SLICE_X104Y128_DQ),
.I3(CLBLM_L_X70Y128_SLICE_X104Y128_AQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X70Y126_SLICE_X105Y126_CO6),
.O5(CLBLM_L_X70Y128_SLICE_X104Y128_DO5),
.O6(CLBLM_L_X70Y128_SLICE_X104Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaccaaccaa)
  ) CLBLM_L_X70Y128_SLICE_X104Y128_CLUT (
.I0(CLBLM_L_X70Y128_SLICE_X104Y128_BQ),
.I1(CLBLM_L_X70Y128_SLICE_X104Y128_CQ),
.I2(CLBLM_L_X70Y128_SLICE_X105Y128_AO6),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(1'b1),
.I5(CLBLM_L_X70Y126_SLICE_X105Y126_CO6),
.O5(CLBLM_L_X70Y128_SLICE_X104Y128_CO5),
.O6(CLBLM_L_X70Y128_SLICE_X104Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff500a0ffff0fff)
  ) CLBLM_L_X70Y128_SLICE_X104Y128_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(1'b1),
.I2(CLBLM_L_X70Y128_SLICE_X104Y128_AQ),
.I3(CLBLM_L_X70Y126_SLICE_X105Y126_CO6),
.I4(CLBLM_L_X70Y129_SLICE_X104Y129_AQ),
.I5(1'b1),
.O5(CLBLM_L_X70Y128_SLICE_X104Y128_BO5),
.O6(CLBLM_L_X70Y128_SLICE_X104Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfcfcff5dda088)
  ) CLBLM_L_X70Y128_SLICE_X104Y128_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X70Y128_SLICE_X104Y128_BQ),
.I2(CLBLM_L_X70Y128_SLICE_X104Y128_AQ),
.I3(CLBLM_L_X70Y126_SLICE_X105Y126_CO6),
.I4(CLBLM_L_X70Y128_SLICE_X105Y128_AQ),
.I5(1'b1),
.O5(CLBLM_L_X70Y128_SLICE_X104Y128_AO5),
.O6(CLBLM_L_X70Y128_SLICE_X104Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y128_SLICE_X105Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y128_SLICE_X104Y128_AQ),
.Q(CLBLM_L_X70Y128_SLICE_X105Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y128_SLICE_X105Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y128_SLICE_X105Y128_DO5),
.O6(CLBLM_L_X70Y128_SLICE_X105Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff050fffff55ff)
  ) CLBLM_L_X70Y128_SLICE_X105Y128_CLUT (
.I0(CLBLM_L_X70Y129_SLICE_X104Y129_AQ),
.I1(1'b1),
.I2(CLBLM_L_X70Y130_SLICE_X105Y130_CQ),
.I3(CLBLM_L_X70Y129_SLICE_X105Y129_BQ),
.I4(CLBLM_L_X70Y128_SLICE_X104Y128_AQ),
.I5(CLBLM_L_X70Y128_SLICE_X104Y128_BQ),
.O5(CLBLM_L_X70Y128_SLICE_X105Y128_CO5),
.O6(CLBLM_L_X70Y128_SLICE_X105Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0cff00000c0c0000)
  ) CLBLM_L_X70Y128_SLICE_X105Y128_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X70Y130_SLICE_X105Y130_BQ),
.I2(CLBLM_L_X70Y129_SLICE_X104Y129_AQ),
.I3(CLBLM_L_X70Y128_SLICE_X104Y128_BQ),
.I4(CLBLM_L_X70Y128_SLICE_X104Y128_AQ),
.I5(CLBLM_L_X70Y129_SLICE_X105Y129_CQ),
.O5(CLBLM_L_X70Y128_SLICE_X105Y128_BO5),
.O6(CLBLM_L_X70Y128_SLICE_X105Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heaafeaaaffffffff)
  ) CLBLM_L_X70Y128_SLICE_X105Y128_ALUT (
.I0(CLBLM_L_X70Y128_SLICE_X105Y128_BO6),
.I1(CLBLM_L_X70Y130_SLICE_X104Y130_BQ),
.I2(CLBLM_L_X70Y129_SLICE_X104Y129_AQ),
.I3(CLBLM_L_X70Y128_SLICE_X104Y128_BQ),
.I4(CLBLM_L_X70Y129_SLICE_X105Y129_AQ),
.I5(CLBLM_L_X70Y128_SLICE_X105Y128_CO6),
.O5(CLBLM_L_X70Y128_SLICE_X105Y128_AO5),
.O6(CLBLM_L_X70Y128_SLICE_X105Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y129_SLICE_X104Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y129_SLICE_X104Y129_AO6),
.Q(CLBLM_L_X70Y129_SLICE_X104Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y129_SLICE_X104Y129_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y129_SLICE_X104Y129_BO6),
.Q(CLBLM_L_X70Y129_SLICE_X104Y129_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y129_SLICE_X104Y129_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y129_SLICE_X104Y129_CO6),
.Q(CLBLM_L_X70Y129_SLICE_X104Y129_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y129_SLICE_X104Y129_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y129_SLICE_X104Y129_DO6),
.Q(CLBLM_L_X70Y129_SLICE_X104Y129_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4ee4e4e4e4e4e4e4)
  ) CLBLM_L_X70Y129_SLICE_X104Y129_DLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X70Y129_SLICE_X104Y129_CQ),
.I2(CLBLM_L_X70Y129_SLICE_X104Y129_DQ),
.I3(CLBLM_L_X70Y126_SLICE_X105Y126_CO6),
.I4(CLBLM_L_X70Y129_SLICE_X104Y129_AQ),
.I5(CLBLM_L_X70Y128_SLICE_X104Y128_BQ),
.O5(CLBLM_L_X70Y129_SLICE_X104Y129_DO5),
.O6(CLBLM_L_X70Y129_SLICE_X104Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd8855aadd88ff00)
  ) CLBLM_L_X70Y129_SLICE_X104Y129_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X70Y129_SLICE_X104Y129_CQ),
.I2(1'b1),
.I3(CLBLM_L_X70Y128_SLICE_X104Y128_DQ),
.I4(CLBLM_L_X70Y128_SLICE_X104Y128_BO5),
.I5(CLBLM_L_X70Y131_SLICE_X104Y131_BQ),
.O5(CLBLM_L_X70Y129_SLICE_X104Y129_CO5),
.O6(CLBLM_L_X70Y129_SLICE_X104Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc5ffc500ccffcc00)
  ) CLBLM_L_X70Y129_SLICE_X104Y129_BLUT (
.I0(CLBLL_R_X71Y130_SLICE_X106Y130_AO6),
.I1(CLBLM_L_X70Y129_SLICE_X104Y129_BQ),
.I2(CLBLM_L_X70Y128_SLICE_X104Y128_AO6),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X70Y129_SLICE_X105Y129_AQ),
.I5(CLBLM_L_X70Y126_SLICE_X105Y126_CO6),
.O5(CLBLM_L_X70Y129_SLICE_X104Y129_BO5),
.O6(CLBLM_L_X70Y129_SLICE_X104Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5055ccccf0f0cccc)
  ) CLBLM_L_X70Y129_SLICE_X104Y129_ALUT (
.I0(CLBLM_L_X70Y128_SLICE_X104Y128_BQ),
.I1(CLBLM_L_X70Y129_SLICE_X104Y129_BQ),
.I2(CLBLM_L_X70Y129_SLICE_X104Y129_AQ),
.I3(CLBLM_L_X70Y128_SLICE_X104Y128_AQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X70Y126_SLICE_X105Y126_CO6),
.O5(CLBLM_L_X70Y129_SLICE_X104Y129_AO5),
.O6(CLBLM_L_X70Y129_SLICE_X104Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y129_SLICE_X105Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y129_SLICE_X105Y129_AO6),
.Q(CLBLM_L_X70Y129_SLICE_X105Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y129_SLICE_X105Y129_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y129_SLICE_X105Y129_BO6),
.Q(CLBLM_L_X70Y129_SLICE_X105Y129_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y129_SLICE_X105Y129_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y129_SLICE_X105Y129_CO6),
.Q(CLBLM_L_X70Y129_SLICE_X105Y129_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y129_SLICE_X105Y129_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y129_SLICE_X105Y129_DO6),
.Q(CLBLM_L_X70Y129_SLICE_X105Y129_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000e1ffe100)
  ) CLBLM_L_X70Y129_SLICE_X105Y129_DLUT (
.I0(CLBLM_L_X70Y130_SLICE_X105Y130_A5Q),
.I1(CLBLM_L_X70Y130_SLICE_X105Y130_AQ),
.I2(CLBLM_L_X70Y129_SLICE_X105Y129_DQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X70Y130_SLICE_X104Y130_DQ),
.I5(CLBLM_L_X72Y132_SLICE_X109Y132_AO6),
.O5(CLBLM_L_X70Y129_SLICE_X105Y129_DO5),
.O6(CLBLM_L_X70Y129_SLICE_X105Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8d8d8d8d8fa50)
  ) CLBLM_L_X70Y129_SLICE_X105Y129_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X70Y129_SLICE_X105Y129_CQ),
.I2(CLBLM_L_X70Y130_SLICE_X105Y130_CQ),
.I3(CLBLM_L_X72Y133_SLICE_X109Y133_AO6),
.I4(CLBLM_L_X72Y132_SLICE_X109Y132_AO6),
.I5(CLBLM_L_X70Y130_SLICE_X105Y130_DO5),
.O5(CLBLM_L_X70Y129_SLICE_X105Y129_CO5),
.O6(CLBLM_L_X70Y129_SLICE_X105Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcafacacaca0acaca)
  ) CLBLM_L_X70Y129_SLICE_X105Y129_BLUT (
.I0(CLBLM_L_X70Y129_SLICE_X105Y129_CQ),
.I1(CLBLM_L_X70Y129_SLICE_X105Y129_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X72Y132_SLICE_X109Y132_AO6),
.I4(CLBLL_R_X71Y130_SLICE_X106Y130_AO6),
.I5(CLBLM_L_X72Y133_SLICE_X109Y133_AO6),
.O5(CLBLM_L_X70Y129_SLICE_X105Y129_BO5),
.O6(CLBLM_L_X70Y129_SLICE_X105Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f0cccca0f0cccc)
  ) CLBLM_L_X70Y129_SLICE_X105Y129_ALUT (
.I0(CLBLM_L_X70Y130_SLICE_X104Y130_AO6),
.I1(CLBLM_L_X70Y129_SLICE_X105Y129_BQ),
.I2(CLBLM_L_X70Y129_SLICE_X105Y129_AQ),
.I3(CLBLM_L_X70Y130_SLICE_X105Y130_A5Q),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X72Y133_SLICE_X109Y133_AO6),
.O5(CLBLM_L_X70Y129_SLICE_X105Y129_AO5),
.O6(CLBLM_L_X70Y129_SLICE_X105Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y130_SLICE_X104Y130_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y130_SLICE_X104Y130_BO6),
.Q(CLBLM_L_X70Y130_SLICE_X104Y130_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y130_SLICE_X104Y130_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y130_SLICE_X104Y130_CO6),
.Q(CLBLM_L_X70Y130_SLICE_X104Y130_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y130_SLICE_X104Y130_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y130_SLICE_X104Y130_DO6),
.Q(CLBLM_L_X70Y130_SLICE_X104Y130_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcce4cce466e466e4)
  ) CLBLM_L_X70Y130_SLICE_X104Y130_DLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X70Y130_SLICE_X104Y130_CQ),
.I2(CLBLM_L_X70Y130_SLICE_X104Y130_DQ),
.I3(CLBLM_L_X70Y130_SLICE_X104Y130_AO5),
.I4(1'b1),
.I5(CLBLM_L_X70Y129_SLICE_X104Y129_DQ),
.O5(CLBLM_L_X70Y130_SLICE_X104Y130_DO5),
.O6(CLBLM_L_X70Y130_SLICE_X104Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcdffcc00c800)
  ) CLBLM_L_X70Y130_SLICE_X104Y130_CLUT (
.I0(CLBLM_L_X70Y130_SLICE_X105Y130_AQ),
.I1(CLBLM_L_X70Y130_SLICE_X104Y130_CQ),
.I2(CLBLM_L_X72Y132_SLICE_X109Y132_AO6),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X70Y130_SLICE_X105Y130_A5Q),
.I5(CLBLM_L_X70Y129_SLICE_X104Y129_DQ),
.O5(CLBLM_L_X70Y130_SLICE_X104Y130_CO5),
.O6(CLBLM_L_X70Y130_SLICE_X104Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500dd88dd88)
  ) CLBLM_L_X70Y130_SLICE_X104Y130_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X70Y130_SLICE_X104Y130_BQ),
.I2(1'b1),
.I3(CLBLM_L_X70Y131_SLICE_X104Y131_BQ),
.I4(CLBLM_L_X72Y133_SLICE_X109Y133_AO6),
.I5(CLBLM_L_X70Y130_SLICE_X104Y130_AO5),
.O5(CLBLM_L_X70Y130_SLICE_X104Y130_BO5),
.O6(CLBLM_L_X70Y130_SLICE_X104Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccffff00001111)
  ) CLBLM_L_X70Y130_SLICE_X104Y130_ALUT (
.I0(CLBLM_L_X70Y130_SLICE_X105Y130_A5Q),
.I1(CLBLM_L_X72Y132_SLICE_X109Y132_AO6),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X70Y130_SLICE_X105Y130_AQ),
.I5(1'b1),
.O5(CLBLM_L_X70Y130_SLICE_X104Y130_AO5),
.O6(CLBLM_L_X70Y130_SLICE_X104Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y130_SLICE_X105Y130_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y130_SLICE_X105Y130_AO5),
.Q(CLBLM_L_X70Y130_SLICE_X105Y130_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y130_SLICE_X105Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y130_SLICE_X105Y130_AO6),
.Q(CLBLM_L_X70Y130_SLICE_X105Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y130_SLICE_X105Y130_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y130_SLICE_X105Y130_BO6),
.Q(CLBLM_L_X70Y130_SLICE_X105Y130_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y130_SLICE_X105Y130_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y130_SLICE_X105Y130_CO6),
.Q(CLBLM_L_X70Y130_SLICE_X105Y130_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccffccf0fff0ff)
  ) CLBLM_L_X70Y130_SLICE_X105Y130_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X72Y132_SLICE_X109Y132_AO6),
.I2(CLBLL_R_X71Y130_SLICE_X106Y130_AQ),
.I3(CLBLM_L_X70Y130_SLICE_X105Y130_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y130_SLICE_X105Y130_DO5),
.O6(CLBLM_L_X70Y130_SLICE_X105Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfc0caaaaaaaa)
  ) CLBLM_L_X70Y130_SLICE_X105Y130_CLUT (
.I0(CLBLM_L_X70Y130_SLICE_X105Y130_BQ),
.I1(CLBLM_L_X70Y130_SLICE_X105Y130_CQ),
.I2(CLBLL_R_X71Y130_SLICE_X106Y130_AQ),
.I3(CLBLM_L_X72Y133_SLICE_X109Y133_AO6),
.I4(CLBLM_L_X70Y130_SLICE_X105Y130_DO6),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X70Y130_SLICE_X105Y130_CO5),
.O6(CLBLM_L_X70Y130_SLICE_X105Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccacaff00ff00)
  ) CLBLM_L_X70Y130_SLICE_X105Y130_BLUT (
.I0(CLBLM_L_X72Y133_SLICE_X109Y133_AO6),
.I1(CLBLM_L_X70Y130_SLICE_X105Y130_BQ),
.I2(CLBLM_L_X70Y130_SLICE_X104Y130_AO6),
.I3(CLBLM_L_X70Y130_SLICE_X104Y130_BQ),
.I4(CLBLL_R_X71Y130_SLICE_X106Y130_AQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X70Y130_SLICE_X105Y130_BO5),
.O6(CLBLM_L_X70Y130_SLICE_X105Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb000b100ddff8800)
  ) CLBLM_L_X70Y130_SLICE_X105Y130_ALUT (
.I0(CLBLM_L_X72Y132_SLICE_X109Y132_AO6),
.I1(CLBLM_L_X70Y130_SLICE_X105Y130_A5Q),
.I2(CLBLM_L_X70Y130_SLICE_X105Y130_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLL_R_X71Y130_SLICE_X106Y130_AQ),
.I5(1'b1),
.O5(CLBLM_L_X70Y130_SLICE_X105Y130_AO5),
.O6(CLBLM_L_X70Y130_SLICE_X105Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y131_SLICE_X104Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y131_SLICE_X104Y131_AO6),
.Q(CLBLM_L_X70Y131_SLICE_X104Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y131_SLICE_X104Y131_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y131_SLICE_X104Y131_BO6),
.Q(CLBLM_L_X70Y131_SLICE_X104Y131_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y131_SLICE_X104Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y131_SLICE_X104Y131_DO5),
.O6(CLBLM_L_X70Y131_SLICE_X104Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y131_SLICE_X104Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y131_SLICE_X104Y131_CO5),
.O6(CLBLM_L_X70Y131_SLICE_X104Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8d8d8d8d8d8f0)
  ) CLBLM_L_X70Y131_SLICE_X104Y131_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X70Y131_SLICE_X104Y131_BQ),
.I2(CLBLM_L_X70Y131_SLICE_X104Y131_AQ),
.I3(CLBLM_L_X72Y132_SLICE_X109Y132_AO6),
.I4(CLBLM_L_X70Y130_SLICE_X105Y130_AQ),
.I5(CLBLM_L_X70Y130_SLICE_X105Y130_A5Q),
.O5(CLBLM_L_X70Y131_SLICE_X104Y131_BO5),
.O6(CLBLM_L_X70Y131_SLICE_X104Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd2ffd2ffd200e200)
  ) CLBLM_L_X70Y131_SLICE_X104Y131_ALUT (
.I0(CLBLM_L_X72Y133_SLICE_X109Y133_AO5),
.I1(CLBLM_L_X72Y132_SLICE_X109Y132_AO6),
.I2(CLBLM_L_X70Y131_SLICE_X104Y131_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X70Y130_SLICE_X105Y130_AQ),
.I5(CLBLM_L_X70Y130_SLICE_X105Y130_A5Q),
.O5(CLBLM_L_X70Y131_SLICE_X104Y131_AO5),
.O6(CLBLM_L_X70Y131_SLICE_X104Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y131_SLICE_X105Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y131_SLICE_X105Y131_DO5),
.O6(CLBLM_L_X70Y131_SLICE_X105Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y131_SLICE_X105Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y131_SLICE_X105Y131_CO5),
.O6(CLBLM_L_X70Y131_SLICE_X105Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y131_SLICE_X105Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y131_SLICE_X105Y131_BO5),
.O6(CLBLM_L_X70Y131_SLICE_X105Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y131_SLICE_X105Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y131_SLICE_X105Y131_AO5),
.O6(CLBLM_L_X70Y131_SLICE_X105Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y132_SLICE_X104Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y132_SLICE_X104Y132_DO5),
.O6(CLBLM_L_X70Y132_SLICE_X104Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y132_SLICE_X104Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y132_SLICE_X104Y132_CO5),
.O6(CLBLM_L_X70Y132_SLICE_X104Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y132_SLICE_X104Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y132_SLICE_X104Y132_BO5),
.O6(CLBLM_L_X70Y132_SLICE_X104Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y132_SLICE_X104Y132_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y132_SLICE_X104Y132_AO5),
.O6(CLBLM_L_X70Y132_SLICE_X104Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y132_SLICE_X105Y132_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y135_SLICE_X105Y135_AQ),
.Q(CLBLM_L_X70Y132_SLICE_X105Y132_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y132_SLICE_X105Y132_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y133_SLICE_X104Y133_A5Q),
.Q(CLBLM_L_X70Y132_SLICE_X105Y132_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y132_SLICE_X105Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y132_SLICE_X105Y132_DO5),
.O6(CLBLM_L_X70Y132_SLICE_X105Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y132_SLICE_X105Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y132_SLICE_X105Y132_CO5),
.O6(CLBLM_L_X70Y132_SLICE_X105Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y132_SLICE_X105Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y132_SLICE_X105Y132_BO5),
.O6(CLBLM_L_X70Y132_SLICE_X105Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y132_SLICE_X105Y132_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y132_SLICE_X105Y132_AO5),
.O6(CLBLM_L_X70Y132_SLICE_X105Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y133_SLICE_X104Y133_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y133_SLICE_X104Y133_CO6),
.Q(CLBLM_L_X70Y133_SLICE_X104Y133_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y133_SLICE_X104Y133_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y133_SLICE_X104Y133_AO6),
.Q(CLBLM_L_X70Y133_SLICE_X104Y133_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y133_SLICE_X104Y133_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y133_SLICE_X104Y133_BO6),
.Q(CLBLM_L_X70Y133_SLICE_X104Y133_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff9fff8fff1fff0)
  ) CLBLM_L_X70Y133_SLICE_X104Y133_DLUT (
.I0(CLBLM_L_X70Y133_SLICE_X105Y133_AQ),
.I1(CLBLM_L_X70Y133_SLICE_X104Y133_AQ),
.I2(CLBLM_L_X70Y134_SLICE_X104Y134_DO6),
.I3(CLBLM_L_X70Y134_SLICE_X104Y134_CO6),
.I4(CLBLM_L_X70Y134_SLICE_X104Y134_AQ),
.I5(CLBLM_L_X70Y134_SLICE_X105Y134_BQ),
.O5(CLBLM_L_X70Y133_SLICE_X104Y133_DO5),
.O6(CLBLM_L_X70Y133_SLICE_X104Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8ccd8ccdfdfdfdf)
  ) CLBLM_L_X70Y133_SLICE_X104Y133_CLUT (
.I0(CLBLM_L_X70Y124_SLICE_X105Y124_AO6),
.I1(CLBLM_L_X70Y133_SLICE_X104Y133_AQ),
.I2(CLBLM_L_X70Y133_SLICE_X104Y133_A5Q),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y133_SLICE_X104Y133_CO5),
.O6(CLBLM_L_X70Y133_SLICE_X104Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5ccc5cccffff0000)
  ) CLBLM_L_X70Y133_SLICE_X104Y133_BLUT (
.I0(CLBLL_R_X71Y133_SLICE_X106Y133_AO6),
.I1(CLBLM_L_X70Y133_SLICE_X104Y133_BQ),
.I2(CLBLM_L_X70Y124_SLICE_X105Y124_AO6),
.I3(CLBLM_L_X70Y134_SLICE_X104Y134_CO5),
.I4(CLBLM_L_X70Y134_SLICE_X104Y134_AQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X70Y133_SLICE_X104Y133_BO5),
.O6(CLBLM_L_X70Y133_SLICE_X104Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0accaacc0accfacc)
  ) CLBLM_L_X70Y133_SLICE_X104Y133_ALUT (
.I0(CLBLM_L_X70Y133_SLICE_X104Y133_AQ),
.I1(CLBLM_L_X70Y133_SLICE_X104Y133_BQ),
.I2(CLBLM_L_X70Y124_SLICE_X105Y124_AO6),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X70Y133_SLICE_X105Y133_AQ),
.I5(CLBLM_L_X70Y133_SLICE_X104Y133_A5Q),
.O5(CLBLM_L_X70Y133_SLICE_X104Y133_AO5),
.O6(CLBLM_L_X70Y133_SLICE_X104Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y133_SLICE_X105Y133_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y133_SLICE_X105Y133_AO6),
.Q(CLBLM_L_X70Y133_SLICE_X105Y133_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y133_SLICE_X105Y133_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y133_SLICE_X105Y133_BO6),
.Q(CLBLM_L_X70Y133_SLICE_X105Y133_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y133_SLICE_X105Y133_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y133_SLICE_X105Y133_CO6),
.Q(CLBLM_L_X70Y133_SLICE_X105Y133_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y133_SLICE_X105Y133_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y133_SLICE_X105Y133_DO6),
.Q(CLBLM_L_X70Y133_SLICE_X105Y133_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he466e466e4cce4cc)
  ) CLBLM_L_X70Y133_SLICE_X105Y133_DLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X70Y133_SLICE_X105Y133_CQ),
.I2(CLBLM_L_X70Y133_SLICE_X105Y133_DQ),
.I3(CLBLM_L_X70Y133_SLICE_X104Y133_CO5),
.I4(1'b1),
.I5(CLBLM_L_X70Y134_SLICE_X105Y134_CQ),
.O5(CLBLM_L_X70Y133_SLICE_X105Y133_DO5),
.O6(CLBLM_L_X70Y133_SLICE_X105Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6ce46c6cf0f0f0f0)
  ) CLBLM_L_X70Y133_SLICE_X105Y133_CLUT (
.I0(CLBLM_L_X70Y124_SLICE_X105Y124_AO6),
.I1(CLBLM_L_X70Y133_SLICE_X105Y133_CQ),
.I2(CLBLM_L_X70Y133_SLICE_X105Y133_BQ),
.I3(CLBLM_L_X70Y133_SLICE_X104Y133_AQ),
.I4(CLBLM_L_X70Y133_SLICE_X104Y133_A5Q),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X70Y133_SLICE_X105Y133_CO5),
.O6(CLBLM_L_X70Y133_SLICE_X105Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc30fcfcfc303030)
  ) CLBLM_L_X70Y133_SLICE_X105Y133_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_L_X70Y133_SLICE_X105Y133_AQ),
.I3(CLBLM_L_X70Y133_SLICE_X104Y133_DO6),
.I4(CLBLM_L_X70Y124_SLICE_X105Y124_AO6),
.I5(CLBLM_L_X70Y133_SLICE_X105Y133_BQ),
.O5(CLBLM_L_X70Y133_SLICE_X105Y133_BO5),
.O6(CLBLM_L_X70Y133_SLICE_X105Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88f3c0bb88f3c0)
  ) CLBLM_L_X70Y133_SLICE_X105Y133_ALUT (
.I0(CLBLM_L_X70Y133_SLICE_X104Y133_A5Q),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_L_X70Y133_SLICE_X105Y133_AQ),
.I3(CLBLM_L_X70Y132_SLICE_X105Y132_BQ),
.I4(CLBLM_L_X70Y124_SLICE_X105Y124_AO6),
.I5(1'b1),
.O5(CLBLM_L_X70Y133_SLICE_X105Y133_AO5),
.O6(CLBLM_L_X70Y133_SLICE_X105Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y134_SLICE_X104Y134_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y134_SLICE_X104Y134_AO6),
.Q(CLBLM_L_X70Y134_SLICE_X104Y134_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y134_SLICE_X104Y134_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y134_SLICE_X104Y134_BO6),
.Q(CLBLM_L_X70Y134_SLICE_X104Y134_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5450545044004400)
  ) CLBLM_L_X70Y134_SLICE_X104Y134_DLUT (
.I0(CLBLM_L_X70Y133_SLICE_X104Y133_A5Q),
.I1(CLBLM_L_X70Y133_SLICE_X105Y133_AQ),
.I2(CLBLM_L_X70Y134_SLICE_X104Y134_BQ),
.I3(CLBLM_L_X70Y135_SLICE_X104Y135_AQ),
.I4(1'b1),
.I5(CLBLM_L_X70Y133_SLICE_X104Y133_AQ),
.O5(CLBLM_L_X70Y134_SLICE_X104Y134_DO5),
.O6(CLBLM_L_X70Y134_SLICE_X104Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c8c00880c0c0c0c)
  ) CLBLM_L_X70Y134_SLICE_X104Y134_CLUT (
.I0(CLBLM_L_X70Y134_SLICE_X105Y134_AQ),
.I1(CLBLM_L_X70Y133_SLICE_X104Y133_A5Q),
.I2(CLBLM_L_X70Y133_SLICE_X105Y133_AQ),
.I3(CLBLM_L_X70Y133_SLICE_X104Y133_AQ),
.I4(CLBLM_L_X70Y135_SLICE_X104Y135_BQ),
.I5(1'b1),
.O5(CLBLM_L_X70Y134_SLICE_X104Y134_CO5),
.O6(CLBLM_L_X70Y134_SLICE_X104Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88f5a0dd88)
  ) CLBLM_L_X70Y134_SLICE_X104Y134_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X70Y134_SLICE_X104Y134_BQ),
.I2(CLBLM_L_X72Y134_SLICE_X109Y134_AO6),
.I3(CLBLM_L_X70Y135_SLICE_X104Y135_BQ),
.I4(CLBLL_R_X71Y133_SLICE_X106Y133_AO6),
.I5(CLBLM_L_X72Y133_SLICE_X109Y133_CO6),
.O5(CLBLM_L_X70Y134_SLICE_X104Y134_BO5),
.O6(CLBLM_L_X70Y134_SLICE_X104Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3aac0aaf0aaf0aa)
  ) CLBLM_L_X70Y134_SLICE_X104Y134_ALUT (
.I0(CLBLM_L_X70Y134_SLICE_X104Y134_BQ),
.I1(CLBLM_L_X70Y134_SLICE_X105Y134_DO5),
.I2(CLBLM_L_X70Y134_SLICE_X104Y134_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X72Y134_SLICE_X109Y134_AO6),
.I5(CLBLM_L_X70Y135_SLICE_X105Y135_A5Q),
.O5(CLBLM_L_X70Y134_SLICE_X104Y134_AO5),
.O6(CLBLM_L_X70Y134_SLICE_X104Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y134_SLICE_X105Y134_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y134_SLICE_X105Y134_AO6),
.Q(CLBLM_L_X70Y134_SLICE_X105Y134_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y134_SLICE_X105Y134_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y134_SLICE_X105Y134_BO6),
.Q(CLBLM_L_X70Y134_SLICE_X105Y134_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y134_SLICE_X105Y134_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y134_SLICE_X105Y134_CO6),
.Q(CLBLM_L_X70Y134_SLICE_X105Y134_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00001111ffff5555)
  ) CLBLM_L_X70Y134_SLICE_X105Y134_DLUT (
.I0(CLBLM_L_X70Y135_SLICE_X105Y135_AQ),
.I1(CLBLM_L_X70Y135_SLICE_X105Y135_A5Q),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X72Y133_SLICE_X109Y133_CO6),
.I5(1'b1),
.O5(CLBLM_L_X70Y134_SLICE_X105Y134_DO5),
.O6(CLBLM_L_X70Y134_SLICE_X105Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0ffe00f001f00)
  ) CLBLM_L_X70Y134_SLICE_X105Y134_CLUT (
.I0(CLBLM_L_X70Y135_SLICE_X105Y135_AQ),
.I1(CLBLM_L_X70Y135_SLICE_X105Y135_A5Q),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLL_R_X71Y134_SLICE_X106Y134_BQ),
.I4(CLBLM_L_X72Y133_SLICE_X109Y133_CO6),
.I5(CLBLM_L_X70Y134_SLICE_X105Y134_CQ),
.O5(CLBLM_L_X70Y134_SLICE_X105Y134_CO5),
.O6(CLBLM_L_X70Y134_SLICE_X105Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44f0f0ee44f0f0)
  ) CLBLM_L_X70Y134_SLICE_X105Y134_BLUT (
.I0(CLBLM_L_X70Y134_SLICE_X105Y134_DO6),
.I1(CLBLM_L_X70Y134_SLICE_X105Y134_BQ),
.I2(CLBLM_L_X70Y134_SLICE_X105Y134_CQ),
.I3(CLBLM_L_X72Y134_SLICE_X109Y134_AO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLM_L_X70Y134_SLICE_X105Y134_BO5),
.O6(CLBLM_L_X70Y134_SLICE_X105Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f5f0a0cccccccc)
  ) CLBLM_L_X70Y134_SLICE_X105Y134_ALUT (
.I0(CLBLL_R_X71Y133_SLICE_X106Y133_AQ),
.I1(CLBLM_L_X70Y134_SLICE_X105Y134_BQ),
.I2(CLBLM_L_X70Y134_SLICE_X105Y134_AQ),
.I3(CLBLM_L_X70Y134_SLICE_X105Y134_DO5),
.I4(CLBLM_L_X72Y134_SLICE_X109Y134_AO6),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X70Y134_SLICE_X105Y134_AO5),
.O6(CLBLM_L_X70Y134_SLICE_X105Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y135_SLICE_X104Y135_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y135_SLICE_X104Y135_AO6),
.Q(CLBLM_L_X70Y135_SLICE_X104Y135_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y135_SLICE_X104Y135_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y135_SLICE_X104Y135_BO6),
.Q(CLBLM_L_X70Y135_SLICE_X104Y135_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y135_SLICE_X104Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y135_SLICE_X104Y135_DO5),
.O6(CLBLM_L_X70Y135_SLICE_X104Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h44444444fcfcfcfc)
  ) CLBLM_L_X70Y135_SLICE_X104Y135_CLUT (
.I0(CLBLL_R_X71Y133_SLICE_X106Y133_AQ),
.I1(CLBLM_L_X70Y135_SLICE_X105Y135_A5Q),
.I2(CLBLM_L_X72Y133_SLICE_X109Y133_CO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y135_SLICE_X104Y135_CO5),
.O6(CLBLM_L_X70Y135_SLICE_X104Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8fa50d8d8d8d8)
  ) CLBLM_L_X70Y135_SLICE_X104Y135_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X70Y135_SLICE_X104Y135_BQ),
.I2(CLBLM_L_X70Y135_SLICE_X104Y135_AQ),
.I3(CLBLM_L_X72Y134_SLICE_X109Y134_AO6),
.I4(CLBLM_L_X72Y133_SLICE_X109Y133_CO6),
.I5(CLBLM_L_X70Y135_SLICE_X104Y135_CO6),
.O5(CLBLM_L_X70Y135_SLICE_X104Y135_BO5),
.O6(CLBLM_L_X70Y135_SLICE_X104Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2eee2e2e222e2)
  ) CLBLM_L_X70Y135_SLICE_X104Y135_ALUT (
.I0(CLBLM_L_X70Y134_SLICE_X105Y134_AQ),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_L_X70Y135_SLICE_X104Y135_AQ),
.I3(CLBLL_R_X71Y133_SLICE_X106Y133_AQ),
.I4(CLBLM_L_X70Y135_SLICE_X104Y135_CO5),
.I5(CLBLM_L_X72Y134_SLICE_X109Y134_AO6),
.O5(CLBLM_L_X70Y135_SLICE_X104Y135_AO5),
.O6(CLBLM_L_X70Y135_SLICE_X104Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y135_SLICE_X105Y135_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y135_SLICE_X105Y135_AO5),
.Q(CLBLM_L_X70Y135_SLICE_X105Y135_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y135_SLICE_X105Y135_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y135_SLICE_X105Y135_AO6),
.Q(CLBLM_L_X70Y135_SLICE_X105Y135_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y135_SLICE_X105Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y135_SLICE_X105Y135_DO5),
.O6(CLBLM_L_X70Y135_SLICE_X105Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y135_SLICE_X105Y135_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y135_SLICE_X105Y135_CO5),
.O6(CLBLM_L_X70Y135_SLICE_X105Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y135_SLICE_X105Y135_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y135_SLICE_X105Y135_BO5),
.O6(CLBLM_L_X70Y135_SLICE_X105Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8080c0c4ff887700)
  ) CLBLM_L_X70Y135_SLICE_X105Y135_ALUT (
.I0(CLBLM_L_X72Y133_SLICE_X109Y133_CO6),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_L_X70Y135_SLICE_X105Y135_AQ),
.I3(CLBLL_R_X71Y133_SLICE_X106Y133_AQ),
.I4(CLBLM_L_X70Y135_SLICE_X105Y135_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X70Y135_SLICE_X105Y135_AO5),
.O6(CLBLM_L_X70Y135_SLICE_X105Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y136_SLICE_X104Y136_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y136_SLICE_X104Y136_AO6),
.Q(CLBLM_L_X70Y136_SLICE_X104Y136_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y136_SLICE_X104Y136_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y136_SLICE_X104Y136_BO6),
.Q(CLBLM_L_X70Y136_SLICE_X104Y136_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y136_SLICE_X104Y136_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y136_SLICE_X104Y136_DO5),
.O6(CLBLM_L_X70Y136_SLICE_X104Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y136_SLICE_X104Y136_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y136_SLICE_X104Y136_CO5),
.O6(CLBLM_L_X70Y136_SLICE_X104Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h46aaccaaccaaccaa)
  ) CLBLM_L_X70Y136_SLICE_X104Y136_BLUT (
.I0(CLBLM_L_X70Y136_SLICE_X105Y136_BQ),
.I1(CLBLM_L_X70Y136_SLICE_X104Y136_BQ),
.I2(CLBLM_L_X70Y136_SLICE_X104Y136_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X70Y136_SLICE_X105Y136_AQ),
.I5(CLBLL_R_X73Y133_SLICE_X111Y133_A5Q),
.O5(CLBLM_L_X70Y136_SLICE_X104Y136_BO5),
.O6(CLBLM_L_X70Y136_SLICE_X104Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h58ccf0ccf0ccf0cc)
  ) CLBLM_L_X70Y136_SLICE_X104Y136_ALUT (
.I0(CLBLM_L_X70Y136_SLICE_X105Y136_BQ),
.I1(CLBLM_L_X70Y136_SLICE_X104Y136_BQ),
.I2(CLBLM_L_X70Y136_SLICE_X104Y136_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X70Y136_SLICE_X105Y136_AQ),
.I5(CLBLL_R_X73Y133_SLICE_X111Y133_A5Q),
.O5(CLBLM_L_X70Y136_SLICE_X104Y136_AO5),
.O6(CLBLM_L_X70Y136_SLICE_X104Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y136_SLICE_X105Y136_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y136_SLICE_X105Y136_AO5),
.Q(CLBLM_L_X70Y136_SLICE_X105Y136_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y136_SLICE_X105Y136_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y136_SLICE_X105Y136_AO6),
.Q(CLBLM_L_X70Y136_SLICE_X105Y136_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y136_SLICE_X105Y136_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y136_SLICE_X105Y136_BO6),
.Q(CLBLM_L_X70Y136_SLICE_X105Y136_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y136_SLICE_X105Y136_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y136_SLICE_X105Y136_DO5),
.O6(CLBLM_L_X70Y136_SLICE_X105Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000040004)
  ) CLBLM_L_X70Y136_SLICE_X105Y136_CLUT (
.I0(CLBLM_L_X70Y136_SLICE_X104Y136_AQ),
.I1(CLBLL_R_X75Y133_SLICE_X115Y133_BQ),
.I2(CLBLM_L_X70Y136_SLICE_X105Y136_BQ),
.I3(CLBLM_L_X70Y136_SLICE_X105Y136_AQ),
.I4(1'b1),
.I5(CLBLM_L_X70Y136_SLICE_X104Y136_BQ),
.O5(CLBLM_L_X70Y136_SLICE_X105Y136_CO5),
.O6(CLBLM_L_X70Y136_SLICE_X105Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6aca6aca88000000)
  ) CLBLM_L_X70Y136_SLICE_X105Y136_BLUT (
.I0(CLBLM_L_X70Y136_SLICE_X105Y136_AQ),
.I1(CLBLM_L_X70Y136_SLICE_X105Y136_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLL_R_X73Y133_SLICE_X111Y133_A5Q),
.I4(CLBLM_L_X70Y136_SLICE_X104Y136_AQ),
.I5(1'b1),
.O5(CLBLM_L_X70Y136_SLICE_X105Y136_BO5),
.O6(CLBLM_L_X70Y136_SLICE_X105Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3ccc3cccaaffaa00)
  ) CLBLM_L_X70Y136_SLICE_X105Y136_ALUT (
.I0(CLBLM_L_X76Y125_SLICE_X116Y125_AQ),
.I1(CLBLL_R_X73Y133_SLICE_X111Y133_A5Q),
.I2(CLBLM_L_X70Y136_SLICE_X105Y136_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X70Y136_SLICE_X104Y136_AQ),
.I5(1'b1),
.O5(CLBLM_L_X70Y136_SLICE_X105Y136_AO5),
.O6(CLBLM_L_X70Y136_SLICE_X105Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y98_SLICE_X108Y98_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y118_SLICE_X108Y118_D5Q),
.Q(CLBLM_L_X72Y98_SLICE_X108Y98_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y98_SLICE_X108Y98_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y119_SLICE_X108Y119_C5Q),
.Q(CLBLM_L_X72Y98_SLICE_X108Y98_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y98_SLICE_X108Y98_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y98_SLICE_X108Y98_AO6),
.Q(CLBLM_L_X72Y98_SLICE_X108Y98_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y98_SLICE_X108Y98_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y98_SLICE_X108Y98_BO6),
.Q(CLBLM_L_X72Y98_SLICE_X108Y98_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y98_SLICE_X108Y98_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y98_SLICE_X108Y98_DO5),
.O6(CLBLM_L_X72Y98_SLICE_X108Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y98_SLICE_X108Y98_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y98_SLICE_X108Y98_CO5),
.O6(CLBLM_L_X72Y98_SLICE_X108Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0d0c0d0caaaaaaaa)
  ) CLBLM_L_X72Y98_SLICE_X108Y98_BLUT (
.I0(CLBLM_L_X72Y98_SLICE_X108Y98_B5Q),
.I1(CLBLM_L_X72Y98_SLICE_X108Y98_BQ),
.I2(CLBLM_L_X68Y98_SLICE_X103Y98_AQ),
.I3(CLBLM_L_X72Y119_SLICE_X108Y119_C5Q),
.I4(1'b1),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X72Y98_SLICE_X108Y98_BO5),
.O6(CLBLM_L_X72Y98_SLICE_X108Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55f555f500aa00a0)
  ) CLBLM_L_X72Y98_SLICE_X108Y98_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(1'b1),
.I2(CLBLM_L_X72Y98_SLICE_X108Y98_AQ),
.I3(CLBLL_R_X71Y98_SLICE_X106Y98_AQ),
.I4(CLBLM_L_X72Y118_SLICE_X108Y118_D5Q),
.I5(CLBLM_L_X72Y98_SLICE_X108Y98_A5Q),
.O5(CLBLM_L_X72Y98_SLICE_X108Y98_AO5),
.O6(CLBLM_L_X72Y98_SLICE_X108Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y98_SLICE_X109Y98_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y98_SLICE_X109Y98_DO5),
.O6(CLBLM_L_X72Y98_SLICE_X109Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y98_SLICE_X109Y98_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y98_SLICE_X109Y98_CO5),
.O6(CLBLM_L_X72Y98_SLICE_X109Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y98_SLICE_X109Y98_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y98_SLICE_X109Y98_BO5),
.O6(CLBLM_L_X72Y98_SLICE_X109Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y98_SLICE_X109Y98_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y98_SLICE_X109Y98_AO5),
.O6(CLBLM_L_X72Y98_SLICE_X109Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y103_SLICE_X108Y103_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y103_SLICE_X108Y103_AO5),
.Q(CLBLM_L_X72Y103_SLICE_X108Y103_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y103_SLICE_X108Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y103_SLICE_X108Y103_AO6),
.Q(CLBLM_L_X72Y103_SLICE_X108Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbbbbb77777777)
  ) CLBLM_L_X72Y103_SLICE_X108Y103_DLUT (
.I0(CLBLM_L_X72Y104_SLICE_X109Y104_AQ),
.I1(CLBLM_L_X72Y103_SLICE_X108Y103_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y103_SLICE_X108Y103_DO5),
.O6(CLBLM_L_X72Y103_SLICE_X108Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f3f3fcfcfcfc)
  ) CLBLM_L_X72Y103_SLICE_X108Y103_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X72Y104_SLICE_X109Y104_A5Q),
.I2(CLBLL_R_X73Y104_SLICE_X110Y104_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y103_SLICE_X108Y103_CO5),
.O6(CLBLM_L_X72Y103_SLICE_X108Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffccff00ffff)
  ) CLBLM_L_X72Y103_SLICE_X108Y103_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X72Y103_SLICE_X108Y103_A5Q),
.I2(1'b1),
.I3(CLBLM_L_X72Y103_SLICE_X108Y103_AQ),
.I4(CLBLM_L_X72Y104_SLICE_X109Y104_AQ),
.I5(1'b1),
.O5(CLBLM_L_X72Y103_SLICE_X108Y103_BO5),
.O6(CLBLM_L_X72Y103_SLICE_X108Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ffff0003f000f00)
  ) CLBLM_L_X72Y103_SLICE_X108Y103_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X72Y103_SLICE_X108Y103_A5Q),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X72Y103_SLICE_X108Y103_AQ),
.I4(CLBLM_L_X72Y104_SLICE_X109Y104_AQ),
.I5(1'b1),
.O5(CLBLM_L_X72Y103_SLICE_X108Y103_AO5),
.O6(CLBLM_L_X72Y103_SLICE_X108Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y103_SLICE_X109Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y103_SLICE_X110Y103_A5Q),
.Q(CLBLM_L_X72Y103_SLICE_X109Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y103_SLICE_X109Y103_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y103_SLICE_X109Y103_BO6),
.Q(CLBLM_L_X72Y103_SLICE_X109Y103_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000aca00c00)
  ) CLBLM_L_X72Y103_SLICE_X109Y103_DLUT (
.I0(CLBLM_L_X72Y103_SLICE_X109Y103_BQ),
.I1(CLBLL_R_X73Y104_SLICE_X110Y104_CQ),
.I2(CLBLM_L_X72Y104_SLICE_X109Y104_B5Q),
.I3(CLBLL_R_X73Y103_SLICE_X110Y103_A5Q),
.I4(CLBLM_L_X72Y103_SLICE_X109Y103_AQ),
.I5(CLBLM_L_X72Y104_SLICE_X109Y104_BQ),
.O5(CLBLM_L_X72Y103_SLICE_X109Y103_DO5),
.O6(CLBLM_L_X72Y103_SLICE_X109Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h70f0f0f0f0f0f0f0)
  ) CLBLM_L_X72Y103_SLICE_X109Y103_CLUT (
.I0(CLBLM_L_X70Y105_SLICE_X104Y105_BO6),
.I1(CLBLL_R_X73Y104_SLICE_X110Y104_A5Q),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X60Y101_SLICE_X90Y101_AQ),
.I4(CLBLM_L_X72Y104_SLICE_X109Y104_B5Q),
.I5(CLBLM_L_X72Y104_SLICE_X109Y104_BQ),
.O5(CLBLM_L_X72Y103_SLICE_X109Y103_CO5),
.O6(CLBLM_L_X72Y103_SLICE_X109Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccfaaaaccc0aaaa)
  ) CLBLM_L_X72Y103_SLICE_X109Y103_BLUT (
.I0(CLBLL_R_X73Y104_SLICE_X110Y104_CQ),
.I1(CLBLM_L_X72Y103_SLICE_X109Y103_BQ),
.I2(CLBLM_L_X72Y103_SLICE_X108Y103_CO5),
.I3(CLBLM_L_X72Y103_SLICE_X108Y103_BO5),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.O5(CLBLM_L_X72Y103_SLICE_X109Y103_BO5),
.O6(CLBLM_L_X72Y103_SLICE_X109Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000550055)
  ) CLBLM_L_X72Y103_SLICE_X109Y103_ALUT (
.I0(CLBLM_L_X72Y104_SLICE_X109Y104_B5Q),
.I1(CLBLL_R_X73Y104_SLICE_X110Y104_A5Q),
.I2(CLBLM_L_X60Y101_SLICE_X90Y101_AQ),
.I3(CLBLM_L_X72Y104_SLICE_X109Y104_BQ),
.I4(CLBLM_L_X70Y105_SLICE_X104Y105_BO6),
.I5(1'b1),
.O5(CLBLM_L_X72Y103_SLICE_X109Y103_AO5),
.O6(CLBLM_L_X72Y103_SLICE_X109Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y104_SLICE_X108Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y104_SLICE_X108Y104_AO6),
.Q(CLBLM_L_X72Y104_SLICE_X108Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y104_SLICE_X108Y104_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y104_SLICE_X108Y104_BO6),
.Q(CLBLM_L_X72Y104_SLICE_X108Y104_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y104_SLICE_X108Y104_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y104_SLICE_X108Y104_CO6),
.Q(CLBLM_L_X72Y104_SLICE_X108Y104_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y104_SLICE_X108Y104_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y104_SLICE_X108Y104_DO6),
.Q(CLBLM_L_X72Y104_SLICE_X108Y104_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff30aaaaff30aaaa)
  ) CLBLM_L_X72Y104_SLICE_X108Y104_DLUT (
.I0(CLBLL_R_X73Y104_SLICE_X111Y104_BQ),
.I1(CLBLM_L_X70Y105_SLICE_X104Y105_BO6),
.I2(CLBLM_L_X72Y104_SLICE_X108Y104_DQ),
.I3(CLBLL_R_X73Y103_SLICE_X111Y103_BO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLM_L_X72Y104_SLICE_X108Y104_DO5),
.O6(CLBLM_L_X72Y104_SLICE_X108Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa5a5acacacaca)
  ) CLBLM_L_X72Y104_SLICE_X108Y104_CLUT (
.I0(CLBLM_L_X72Y104_SLICE_X108Y104_BQ),
.I1(CLBLM_L_X72Y104_SLICE_X108Y104_CQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(1'b1),
.I4(CLBLM_L_X72Y105_SLICE_X108Y105_A5Q),
.I5(CLBLL_R_X73Y104_SLICE_X110Y104_BO5),
.O5(CLBLM_L_X72Y104_SLICE_X108Y104_CO5),
.O6(CLBLM_L_X72Y104_SLICE_X108Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hacccccccaaaaaaaa)
  ) CLBLM_L_X72Y104_SLICE_X108Y104_BLUT (
.I0(CLBLM_L_X72Y105_SLICE_X108Y105_A5Q),
.I1(CLBLM_L_X72Y104_SLICE_X108Y104_BQ),
.I2(CLBLM_L_X72Y104_SLICE_X109Y104_A5Q),
.I3(CLBLL_R_X73Y104_SLICE_X110Y104_BQ),
.I4(CLBLM_L_X72Y103_SLICE_X108Y103_A5Q),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X72Y104_SLICE_X108Y104_BO5),
.O6(CLBLM_L_X72Y104_SLICE_X108Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd887d28dd887d28)
  ) CLBLM_L_X72Y104_SLICE_X108Y104_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X73Y103_SLICE_X111Y103_BO6),
.I2(CLBLM_L_X72Y104_SLICE_X108Y104_AQ),
.I3(CLBLM_L_X72Y105_SLICE_X108Y105_BQ),
.I4(CLBLM_L_X72Y103_SLICE_X109Y103_AO6),
.I5(1'b1),
.O5(CLBLM_L_X72Y104_SLICE_X108Y104_AO5),
.O6(CLBLM_L_X72Y104_SLICE_X108Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y104_SLICE_X109Y104_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y104_SLICE_X109Y104_AO5),
.Q(CLBLM_L_X72Y104_SLICE_X109Y104_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y104_SLICE_X109Y104_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y104_SLICE_X109Y104_BO5),
.Q(CLBLM_L_X72Y104_SLICE_X109Y104_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y104_SLICE_X109Y104_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y104_SLICE_X109Y104_CO5),
.Q(CLBLM_L_X72Y104_SLICE_X109Y104_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y104_SLICE_X109Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y104_SLICE_X109Y104_AO6),
.Q(CLBLM_L_X72Y104_SLICE_X109Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y104_SLICE_X109Y104_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y104_SLICE_X109Y104_BO6),
.Q(CLBLM_L_X72Y104_SLICE_X109Y104_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y104_SLICE_X109Y104_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y104_SLICE_X109Y104_CO6),
.Q(CLBLM_L_X72Y104_SLICE_X109Y104_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa5ffc3ff00ff00)
  ) CLBLM_L_X72Y104_SLICE_X109Y104_DLUT (
.I0(CLBLM_L_X72Y104_SLICE_X109Y104_C5Q),
.I1(CLBLM_L_X72Y104_SLICE_X109Y104_CQ),
.I2(CLBLM_L_X72Y104_SLICE_X109Y104_BQ),
.I3(CLBLM_L_X70Y105_SLICE_X105Y105_BQ),
.I4(CLBLM_L_X72Y104_SLICE_X109Y104_B5Q),
.I5(CLBLM_L_X70Y105_SLICE_X104Y105_BO6),
.O5(CLBLM_L_X72Y104_SLICE_X109Y104_DO5),
.O6(CLBLM_L_X72Y104_SLICE_X109Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0555f0f00ccccccc)
  ) CLBLM_L_X72Y104_SLICE_X109Y104_CLUT (
.I0(CLBLM_L_X72Y104_SLICE_X109Y104_C5Q),
.I1(CLBLM_L_X72Y104_SLICE_X109Y104_CQ),
.I2(CLBLL_R_X73Y104_SLICE_X110Y104_A5Q),
.I3(CLBLL_R_X73Y104_SLICE_X111Y104_DO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLM_L_X72Y104_SLICE_X109Y104_CO5),
.O6(CLBLM_L_X72Y104_SLICE_X109Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6fc06fc05faf50a0)
  ) CLBLM_L_X72Y104_SLICE_X109Y104_BLUT (
.I0(CLBLM_L_X70Y105_SLICE_X104Y105_BO6),
.I1(CLBLM_L_X72Y104_SLICE_X109Y104_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X72Y104_SLICE_X109Y104_B5Q),
.I4(CLBLM_L_X72Y104_SLICE_X109Y104_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X72Y104_SLICE_X109Y104_BO5),
.O6(CLBLM_L_X72Y104_SLICE_X109Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0500050066aa66aa)
  ) CLBLM_L_X72Y104_SLICE_X109Y104_ALUT (
.I0(CLBLM_L_X72Y103_SLICE_X108Y103_A5Q),
.I1(CLBLM_L_X72Y104_SLICE_X109Y104_A5Q),
.I2(CLBLM_L_X72Y104_SLICE_X109Y104_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y104_SLICE_X109Y104_AO5),
.O6(CLBLM_L_X72Y104_SLICE_X109Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y105_SLICE_X108Y105_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y105_SLICE_X108Y105_AO5),
.Q(CLBLM_L_X72Y105_SLICE_X108Y105_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y105_SLICE_X108Y105_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y105_SLICE_X108Y105_AO6),
.Q(CLBLM_L_X72Y105_SLICE_X108Y105_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y105_SLICE_X108Y105_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y105_SLICE_X108Y105_BO6),
.Q(CLBLM_L_X72Y105_SLICE_X108Y105_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y105_SLICE_X108Y105_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y105_SLICE_X108Y105_CO6),
.Q(CLBLM_L_X72Y105_SLICE_X108Y105_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y105_SLICE_X108Y105_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y105_SLICE_X108Y105_DO6),
.Q(CLBLM_L_X72Y105_SLICE_X108Y105_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h20a08a0aa0a00a0a)
  ) CLBLM_L_X72Y105_SLICE_X108Y105_DLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X73Y104_SLICE_X110Y104_BQ),
.I2(CLBLM_L_X72Y105_SLICE_X108Y105_DQ),
.I3(CLBLM_L_X72Y104_SLICE_X109Y104_A5Q),
.I4(CLBLL_R_X79Y99_SLICE_X122Y99_AO6),
.I5(CLBLM_L_X72Y103_SLICE_X108Y103_A5Q),
.O5(CLBLM_L_X72Y105_SLICE_X108Y105_DO5),
.O6(CLBLM_L_X72Y105_SLICE_X108Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc5a5aaaaa)
  ) CLBLM_L_X72Y105_SLICE_X108Y105_CLUT (
.I0(CLBLM_L_X72Y104_SLICE_X108Y104_AQ),
.I1(CLBLM_L_X72Y105_SLICE_X108Y105_CQ),
.I2(CLBLM_L_X72Y105_SLICE_X108Y105_BQ),
.I3(1'b1),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X72Y103_SLICE_X109Y103_CO6),
.O5(CLBLM_L_X72Y105_SLICE_X108Y105_CO5),
.O6(CLBLM_L_X72Y105_SLICE_X108Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he4ccf0f0ccccf0f0)
  ) CLBLM_L_X72Y105_SLICE_X108Y105_BLUT (
.I0(CLBLM_L_X72Y103_SLICE_X108Y103_A5Q),
.I1(CLBLM_L_X72Y105_SLICE_X108Y105_BQ),
.I2(CLBLM_L_X72Y105_SLICE_X108Y105_DQ),
.I3(CLBLL_R_X73Y104_SLICE_X110Y104_BQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X72Y104_SLICE_X109Y104_A5Q),
.O5(CLBLM_L_X72Y105_SLICE_X108Y105_BO5),
.O6(CLBLM_L_X72Y105_SLICE_X108Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h550055004e4ee4e4)
  ) CLBLM_L_X72Y105_SLICE_X108Y105_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X72Y105_SLICE_X109Y105_B5Q),
.I2(CLBLM_L_X72Y103_SLICE_X109Y103_AO6),
.I3(CLBLM_L_X72Y128_SLICE_X109Y128_AQ),
.I4(CLBLM_L_X72Y105_SLICE_X108Y105_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X72Y105_SLICE_X108Y105_AO5),
.O6(CLBLM_L_X72Y105_SLICE_X108Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y105_SLICE_X109Y105_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y105_SLICE_X109Y105_BO5),
.Q(CLBLM_L_X72Y105_SLICE_X109Y105_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y105_SLICE_X109Y105_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y105_SLICE_X109Y105_AO6),
.Q(CLBLM_L_X72Y105_SLICE_X109Y105_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y105_SLICE_X109Y105_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y105_SLICE_X109Y105_BO6),
.Q(CLBLM_L_X72Y105_SLICE_X109Y105_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y105_SLICE_X109Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y105_SLICE_X109Y105_DO5),
.O6(CLBLM_L_X72Y105_SLICE_X109Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y105_SLICE_X109Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y105_SLICE_X109Y105_CO5),
.O6(CLBLM_L_X72Y105_SLICE_X109Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccf0aac3aacc)
  ) CLBLM_L_X72Y105_SLICE_X109Y105_BLUT (
.I0(CLBLM_L_X72Y105_SLICE_X109Y105_B5Q),
.I1(CLBLM_L_X72Y105_SLICE_X109Y105_BQ),
.I2(CLBLM_L_X72Y105_SLICE_X109Y105_AQ),
.I3(CLBLM_L_X72Y103_SLICE_X109Y103_CO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLM_L_X72Y105_SLICE_X109Y105_BO5),
.O6(CLBLM_L_X72Y105_SLICE_X109Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h78f0ffff78f00000)
  ) CLBLM_L_X72Y105_SLICE_X109Y105_ALUT (
.I0(CLBLM_L_X72Y104_SLICE_X109Y104_A5Q),
.I1(CLBLM_L_X72Y103_SLICE_X108Y103_A5Q),
.I2(CLBLM_L_X72Y105_SLICE_X109Y105_AQ),
.I3(CLBLL_R_X73Y104_SLICE_X110Y104_BQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X72Y105_SLICE_X108Y105_CQ),
.O5(CLBLM_L_X72Y105_SLICE_X109Y105_AO5),
.O6(CLBLM_L_X72Y105_SLICE_X109Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y106_SLICE_X108Y106_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X78Y106_SLICE_X120Y106_AQ),
.Q(CLBLM_L_X72Y106_SLICE_X108Y106_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y106_SLICE_X108Y106_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y106_SLICE_X108Y106_AO6),
.Q(CLBLM_L_X72Y106_SLICE_X108Y106_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f000f000d000f00)
  ) CLBLM_L_X72Y106_SLICE_X108Y106_DLUT (
.I0(CLBLM_L_X72Y108_SLICE_X108Y108_AQ),
.I1(CLBLL_R_X71Y107_SLICE_X106Y107_C5Q),
.I2(CLBLL_R_X71Y107_SLICE_X107Y107_DO6),
.I3(CLBLL_R_X73Y108_SLICE_X110Y108_A5Q),
.I4(CLBLM_L_X72Y107_SLICE_X109Y107_A5Q),
.I5(CLBLL_R_X71Y107_SLICE_X106Y107_CQ),
.O5(CLBLM_L_X72Y106_SLICE_X108Y106_DO5),
.O6(CLBLM_L_X72Y106_SLICE_X108Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0c0f0c0f0f0f0d0)
  ) CLBLM_L_X72Y106_SLICE_X108Y106_CLUT (
.I0(CLBLL_R_X73Y106_SLICE_X110Y106_BO6),
.I1(CLBLM_L_X72Y106_SLICE_X109Y106_CO6),
.I2(CLBLM_L_X70Y106_SLICE_X105Y106_CO6),
.I3(CLBLM_L_X72Y107_SLICE_X108Y107_CO6),
.I4(CLBLL_R_X73Y107_SLICE_X110Y107_DO6),
.I5(CLBLM_L_X72Y106_SLICE_X108Y106_DO6),
.O5(CLBLM_L_X72Y106_SLICE_X108Y106_CO5),
.O6(CLBLM_L_X72Y106_SLICE_X108Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0004000c0cc4044)
  ) CLBLM_L_X72Y106_SLICE_X108Y106_BLUT (
.I0(CLBLM_L_X72Y107_SLICE_X109Y107_A5Q),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_L_X72Y106_SLICE_X108Y106_AQ),
.I3(CLBLM_L_X78Y106_SLICE_X120Y106_AQ),
.I4(CLBLM_L_X62Y92_SLICE_X92Y92_AQ),
.I5(CLBLM_L_X72Y106_SLICE_X108Y106_A5Q),
.O5(CLBLM_L_X72Y106_SLICE_X108Y106_BO5),
.O6(CLBLM_L_X72Y106_SLICE_X108Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h08882aaa00002222)
  ) CLBLM_L_X72Y106_SLICE_X108Y106_ALUT (
.I0(CLBLM_L_X72Y106_SLICE_X108Y106_BO6),
.I1(CLBLM_L_X62Y90_SLICE_X92Y90_AQ),
.I2(CLBLM_L_X72Y106_SLICE_X108Y106_AQ),
.I3(CLBLM_L_X78Y106_SLICE_X120Y106_AQ),
.I4(CLBLM_L_X62Y92_SLICE_X92Y92_AQ),
.I5(CLBLM_L_X72Y106_SLICE_X108Y106_A5Q),
.O5(CLBLM_L_X72Y106_SLICE_X108Y106_AO5),
.O6(CLBLM_L_X72Y106_SLICE_X108Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y106_SLICE_X109Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y106_SLICE_X109Y106_DO5),
.O6(CLBLM_L_X72Y106_SLICE_X109Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heaeaaaaa00ea00aa)
  ) CLBLM_L_X72Y106_SLICE_X109Y106_CLUT (
.I0(CLBLM_L_X72Y106_SLICE_X109Y106_AO6),
.I1(CLBLM_L_X72Y106_SLICE_X108Y106_A5Q),
.I2(CLBLM_L_X72Y107_SLICE_X109Y107_BO5),
.I3(CLBLM_L_X72Y107_SLICE_X109Y107_CO6),
.I4(CLBLM_L_X74Y107_SLICE_X112Y107_BQ),
.I5(CLBLM_L_X72Y106_SLICE_X109Y106_BO6),
.O5(CLBLM_L_X72Y106_SLICE_X109Y106_CO5),
.O6(CLBLM_L_X72Y106_SLICE_X109Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00400040ffff)
  ) CLBLM_L_X72Y106_SLICE_X109Y106_BLUT (
.I0(CLBLL_R_X71Y107_SLICE_X106Y107_C5Q),
.I1(CLBLL_R_X73Y107_SLICE_X110Y107_BQ),
.I2(CLBLM_L_X78Y106_SLICE_X120Y106_AQ),
.I3(CLBLL_R_X71Y107_SLICE_X106Y107_CQ),
.I4(CLBLM_L_X72Y106_SLICE_X108Y106_AQ),
.I5(CLBLL_R_X73Y108_SLICE_X110Y108_A5Q),
.O5(CLBLM_L_X72Y106_SLICE_X109Y106_BO5),
.O6(CLBLM_L_X72Y106_SLICE_X109Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5575aaba5555aaaa)
  ) CLBLM_L_X72Y106_SLICE_X109Y106_ALUT (
.I0(CLBLL_R_X73Y108_SLICE_X110Y108_A5Q),
.I1(CLBLL_R_X71Y107_SLICE_X106Y107_C5Q),
.I2(CLBLM_L_X62Y90_SLICE_X92Y90_AQ),
.I3(CLBLL_R_X71Y107_SLICE_X106Y107_CQ),
.I4(CLBLM_L_X72Y106_SLICE_X108Y106_AQ),
.I5(CLBLM_L_X74Y107_SLICE_X112Y107_DQ),
.O5(CLBLM_L_X72Y106_SLICE_X109Y106_AO5),
.O6(CLBLM_L_X72Y106_SLICE_X109Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y107_SLICE_X108Y107_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y107_SLICE_X109Y107_BQ),
.Q(CLBLM_L_X72Y107_SLICE_X108Y107_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y107_SLICE_X108Y107_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y107_SLICE_X108Y107_AO6),
.Q(CLBLM_L_X72Y107_SLICE_X108Y107_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y107_SLICE_X108Y107_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y107_SLICE_X108Y107_A5Q),
.Q(CLBLM_L_X72Y107_SLICE_X108Y107_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y107_SLICE_X108Y107_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y107_SLICE_X108Y107_BQ),
.Q(CLBLM_L_X72Y107_SLICE_X108Y107_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h07770fffbbbbffff)
  ) CLBLM_L_X72Y107_SLICE_X108Y107_DLUT (
.I0(CLBLM_L_X72Y106_SLICE_X108Y106_AQ),
.I1(CLBLL_R_X73Y107_SLICE_X110Y107_AQ),
.I2(CLBLM_L_X72Y107_SLICE_X108Y107_A5Q),
.I3(CLBLL_R_X71Y107_SLICE_X107Y107_BQ),
.I4(CLBLM_L_X78Y106_SLICE_X120Y106_AQ),
.I5(CLBLL_R_X73Y108_SLICE_X110Y108_A5Q),
.O5(CLBLM_L_X72Y107_SLICE_X108Y107_DO5),
.O6(CLBLM_L_X72Y107_SLICE_X108Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff5f0fdfc)
  ) CLBLM_L_X72Y107_SLICE_X108Y107_CLUT (
.I0(CLBLL_R_X71Y107_SLICE_X106Y107_BO5),
.I1(CLBLM_L_X72Y107_SLICE_X108Y107_BO5),
.I2(CLBLM_L_X72Y107_SLICE_X109Y107_BO6),
.I3(CLBLM_L_X72Y108_SLICE_X108Y108_DQ),
.I4(CLBLM_L_X72Y107_SLICE_X108Y107_DO6),
.I5(CLBLM_L_X72Y107_SLICE_X108Y107_BO6),
.O5(CLBLM_L_X72Y107_SLICE_X108Y107_CO5),
.O6(CLBLM_L_X72Y107_SLICE_X108Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1000000044444444)
  ) CLBLM_L_X72Y107_SLICE_X108Y107_BLUT (
.I0(CLBLL_R_X71Y107_SLICE_X106Y107_C5Q),
.I1(CLBLL_R_X71Y107_SLICE_X106Y107_CQ),
.I2(CLBLM_L_X72Y107_SLICE_X108Y107_AQ),
.I3(CLBLL_R_X73Y108_SLICE_X110Y108_A5Q),
.I4(CLBLM_L_X72Y107_SLICE_X108Y107_CQ),
.I5(1'b1),
.O5(CLBLM_L_X72Y107_SLICE_X108Y107_BO5),
.O6(CLBLM_L_X72Y107_SLICE_X108Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he4f0ffffe4f00000)
  ) CLBLM_L_X72Y107_SLICE_X108Y107_ALUT (
.I0(CLBLL_R_X71Y109_SLICE_X106Y109_CO6),
.I1(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I2(CLBLM_L_X72Y107_SLICE_X108Y107_AQ),
.I3(CLBLM_L_X72Y108_SLICE_X109Y108_A5Q),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X72Y108_SLICE_X108Y108_CQ),
.O5(CLBLM_L_X72Y107_SLICE_X108Y107_AO5),
.O6(CLBLM_L_X72Y107_SLICE_X108Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y107_SLICE_X109Y107_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y92_SLICE_X92Y92_AQ),
.Q(CLBLM_L_X72Y107_SLICE_X109Y107_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y107_SLICE_X109Y107_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y107_SLICE_X109Y107_AO6),
.Q(CLBLM_L_X72Y107_SLICE_X109Y107_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y107_SLICE_X109Y107_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y107_SLICE_X109Y107_A5Q),
.Q(CLBLM_L_X72Y107_SLICE_X109Y107_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8080808000000000)
  ) CLBLM_L_X72Y107_SLICE_X109Y107_DLUT (
.I0(CLBLM_L_X72Y106_SLICE_X108Y106_AQ),
.I1(CLBLM_L_X72Y106_SLICE_X108Y106_A5Q),
.I2(CLBLM_L_X62Y90_SLICE_X92Y90_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X78Y106_SLICE_X120Y106_AQ),
.O5(CLBLM_L_X72Y107_SLICE_X109Y107_DO5),
.O6(CLBLM_L_X72Y107_SLICE_X109Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbffbbff5f5fffff)
  ) CLBLM_L_X72Y107_SLICE_X109Y107_CLUT (
.I0(CLBLL_R_X71Y107_SLICE_X106Y107_CQ),
.I1(CLBLM_L_X72Y106_SLICE_X108Y106_A5Q),
.I2(CLBLM_L_X72Y108_SLICE_X109Y108_DQ),
.I3(CLBLL_R_X73Y108_SLICE_X110Y108_BQ),
.I4(CLBLM_L_X62Y90_SLICE_X92Y90_AQ),
.I5(CLBLL_R_X71Y107_SLICE_X106Y107_C5Q),
.O5(CLBLM_L_X72Y107_SLICE_X109Y107_CO5),
.O6(CLBLM_L_X72Y107_SLICE_X109Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h20000000cc00cc00)
  ) CLBLM_L_X72Y107_SLICE_X109Y107_BLUT (
.I0(CLBLL_R_X73Y108_SLICE_X110Y108_A5Q),
.I1(CLBLL_R_X71Y107_SLICE_X106Y107_CQ),
.I2(CLBLM_L_X72Y107_SLICE_X109Y107_AQ),
.I3(CLBLL_R_X71Y107_SLICE_X106Y107_C5Q),
.I4(CLBLM_L_X72Y106_SLICE_X108Y106_AQ),
.I5(1'b1),
.O5(CLBLM_L_X72Y107_SLICE_X109Y107_BO5),
.O6(CLBLM_L_X72Y107_SLICE_X109Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f7a0a2f5d5a080)
  ) CLBLM_L_X72Y107_SLICE_X109Y107_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X72Y108_SLICE_X109Y108_CO5),
.I2(CLBLM_L_X72Y107_SLICE_X109Y107_AQ),
.I3(CLBLM_L_X72Y108_SLICE_X108Y108_BO6),
.I4(CLBLM_L_X72Y107_SLICE_X108Y107_AQ),
.I5(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.O5(CLBLM_L_X72Y107_SLICE_X109Y107_AO5),
.O6(CLBLM_L_X72Y107_SLICE_X109Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y108_SLICE_X108Y108_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y108_SLICE_X108Y108_AO6),
.Q(CLBLM_L_X72Y108_SLICE_X108Y108_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y108_SLICE_X108Y108_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y108_SLICE_X108Y108_CO6),
.Q(CLBLM_L_X72Y108_SLICE_X108Y108_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y108_SLICE_X108Y108_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y108_SLICE_X108Y108_DO6),
.Q(CLBLM_L_X72Y108_SLICE_X108Y108_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd75a820fd75a820)
  ) CLBLM_L_X72Y108_SLICE_X108Y108_DLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X71Y109_SLICE_X106Y109_CO5),
.I2(CLBLM_L_X72Y108_SLICE_X108Y108_DQ),
.I3(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I4(CLBLM_L_X72Y108_SLICE_X109Y108_DQ),
.I5(1'b1),
.O5(CLBLM_L_X72Y108_SLICE_X108Y108_DO5),
.O6(CLBLM_L_X72Y108_SLICE_X108Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccd8d8ff00ff00)
  ) CLBLM_L_X72Y108_SLICE_X108Y108_CLUT (
.I0(CLBLM_L_X72Y108_SLICE_X109Y108_CO6),
.I1(CLBLM_L_X72Y108_SLICE_X108Y108_CQ),
.I2(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I3(CLBLL_R_X71Y107_SLICE_X107Y107_BQ),
.I4(CLBLL_R_X71Y109_SLICE_X106Y109_CO6),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X72Y108_SLICE_X108Y108_CO5),
.O6(CLBLM_L_X72Y108_SLICE_X108Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafafaff5f5f5f5)
  ) CLBLM_L_X72Y108_SLICE_X108Y108_BLUT (
.I0(CLBLL_R_X71Y109_SLICE_X106Y109_B5Q),
.I1(1'b1),
.I2(CLBLL_R_X71Y109_SLICE_X106Y109_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y108_SLICE_X108Y108_BO5),
.O6(CLBLM_L_X72Y108_SLICE_X108Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ff55aa00a808)
  ) CLBLM_L_X72Y108_SLICE_X108Y108_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I2(CLBLM_L_X72Y108_SLICE_X109Y108_CO5),
.I3(CLBLM_L_X72Y108_SLICE_X108Y108_AQ),
.I4(CLBLL_R_X71Y109_SLICE_X106Y109_BQ),
.I5(CLBLL_R_X71Y109_SLICE_X106Y109_B5Q),
.O5(CLBLM_L_X72Y108_SLICE_X108Y108_AO5),
.O6(CLBLM_L_X72Y108_SLICE_X108Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y108_SLICE_X109Y108_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y108_SLICE_X109Y108_AO5),
.Q(CLBLM_L_X72Y108_SLICE_X109Y108_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y108_SLICE_X109Y108_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y108_SLICE_X109Y108_AO6),
.Q(CLBLM_L_X72Y108_SLICE_X109Y108_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y108_SLICE_X109Y108_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y108_SLICE_X109Y108_DO6),
.Q(CLBLM_L_X72Y108_SLICE_X109Y108_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4eee4e4e444)
  ) CLBLM_L_X72Y108_SLICE_X109Y108_DLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X73Y108_SLICE_X110Y108_BQ),
.I2(CLBLM_L_X72Y108_SLICE_X109Y108_DQ),
.I3(CLBLM_L_X72Y108_SLICE_X109Y108_CO6),
.I4(CLBLM_L_X72Y109_SLICE_X108Y109_BO6),
.I5(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.O5(CLBLM_L_X72Y108_SLICE_X109Y108_DO5),
.O6(CLBLM_L_X72Y108_SLICE_X109Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3ffffcfffc)
  ) CLBLM_L_X72Y108_SLICE_X109Y108_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X72Y108_SLICE_X109Y108_AQ),
.I2(CLBLL_R_X71Y111_SLICE_X106Y111_AQ),
.I3(CLBLM_L_X72Y108_SLICE_X109Y108_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y108_SLICE_X109Y108_CO5),
.O6(CLBLM_L_X72Y108_SLICE_X109Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ffffffff0f0f)
  ) CLBLM_L_X72Y108_SLICE_X109Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X72Y108_SLICE_X109Y108_AQ),
.I3(1'b1),
.I4(CLBLL_R_X71Y111_SLICE_X106Y111_AQ),
.I5(1'b1),
.O5(CLBLM_L_X72Y108_SLICE_X109Y108_BO5),
.O6(CLBLM_L_X72Y108_SLICE_X109Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff0ff003000f0f0)
  ) CLBLM_L_X72Y108_SLICE_X109Y108_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X72Y108_SLICE_X109Y108_A5Q),
.I2(CLBLM_L_X72Y108_SLICE_X109Y108_AQ),
.I3(CLBLL_R_X71Y111_SLICE_X106Y111_AQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLM_L_X72Y108_SLICE_X109Y108_AO5),
.O6(CLBLM_L_X72Y108_SLICE_X109Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y109_SLICE_X108Y109_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y109_SLICE_X105Y109_AQ),
.Q(CLBLM_L_X72Y109_SLICE_X108Y109_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y109_SLICE_X108Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y109_SLICE_X108Y109_DO5),
.O6(CLBLM_L_X72Y109_SLICE_X108Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y109_SLICE_X108Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y109_SLICE_X108Y109_CO5),
.O6(CLBLM_L_X72Y109_SLICE_X108Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0fffffffff)
  ) CLBLM_L_X72Y109_SLICE_X108Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_R_X71Y109_SLICE_X106Y109_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_R_X71Y109_SLICE_X106Y109_B5Q),
.O5(CLBLM_L_X72Y109_SLICE_X108Y109_BO5),
.O6(CLBLM_L_X72Y109_SLICE_X108Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h66cccccccccccccc)
  ) CLBLM_L_X72Y109_SLICE_X108Y109_ALUT (
.I0(CLBLM_L_X72Y109_SLICE_X109Y109_BQ),
.I1(CLBLM_L_X72Y111_SLICE_X108Y111_CQ),
.I2(1'b1),
.I3(CLBLM_L_X72Y111_SLICE_X109Y111_BQ),
.I4(CLBLM_L_X72Y109_SLICE_X109Y109_AQ),
.I5(CLBLM_L_X72Y109_SLICE_X109Y109_CQ),
.O5(CLBLM_L_X72Y109_SLICE_X108Y109_AO5),
.O6(CLBLM_L_X72Y109_SLICE_X108Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y109_SLICE_X109Y109_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y109_SLICE_X109Y109_AO5),
.Q(CLBLM_L_X72Y109_SLICE_X109Y109_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y109_SLICE_X109Y109_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y109_SLICE_X109Y109_BO5),
.Q(CLBLM_L_X72Y109_SLICE_X109Y109_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y109_SLICE_X109Y109_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y109_SLICE_X109Y109_CO5),
.Q(CLBLM_L_X72Y109_SLICE_X109Y109_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y109_SLICE_X109Y109_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y109_SLICE_X109Y109_AO6),
.Q(CLBLM_L_X72Y109_SLICE_X109Y109_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y109_SLICE_X109Y109_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y109_SLICE_X109Y109_BO6),
.Q(CLBLM_L_X72Y109_SLICE_X109Y109_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y109_SLICE_X109Y109_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y109_SLICE_X109Y109_CO6),
.Q(CLBLM_L_X72Y109_SLICE_X109Y109_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y109_SLICE_X109Y109_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y109_SLICE_X109Y109_DO6),
.Q(CLBLM_L_X72Y109_SLICE_X109Y109_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hecacacacacacacac)
  ) CLBLM_L_X72Y109_SLICE_X109Y109_DLUT (
.I0(CLBLM_L_X72Y116_SLICE_X108Y116_AQ),
.I1(CLBLM_L_X72Y109_SLICE_X109Y109_CQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X72Y109_SLICE_X109Y109_BQ),
.I4(CLBLM_L_X72Y109_SLICE_X109Y109_AQ),
.I5(CLBLM_L_X72Y111_SLICE_X109Y111_BQ),
.O5(CLBLM_L_X72Y109_SLICE_X109Y109_DO5),
.O6(CLBLM_L_X72Y109_SLICE_X109Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88dddd8888)
  ) CLBLM_L_X72Y109_SLICE_X109Y109_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(RIOB33_X105Y59_IOB_X1Y59_I),
.I2(1'b1),
.I3(CLBLM_L_X72Y109_SLICE_X109Y109_BQ),
.I4(CLBLM_L_X72Y109_SLICE_X109Y109_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X72Y109_SLICE_X109Y109_CO5),
.O6(CLBLM_L_X72Y109_SLICE_X109Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaf0ccf0cc)
  ) CLBLM_L_X72Y109_SLICE_X109Y109_BLUT (
.I0(CLBLM_L_X72Y109_SLICE_X109Y109_AQ),
.I1(CLBLM_L_X72Y109_SLICE_X109Y109_A5Q),
.I2(RIOB33_X105Y57_IOB_X1Y58_I),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y109_SLICE_X109Y109_BO5),
.O6(CLBLM_L_X72Y109_SLICE_X109Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaaccaaffaa00)
  ) CLBLM_L_X72Y109_SLICE_X109Y109_ALUT (
.I0(RIOB33_X105Y57_IOB_X1Y57_I),
.I1(CLBLM_L_X72Y111_SLICE_X109Y111_BQ),
.I2(1'b1),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X72Y109_SLICE_X108Y109_AQ),
.I5(1'b1),
.O5(CLBLM_L_X72Y109_SLICE_X109Y109_AO5),
.O6(CLBLM_L_X72Y109_SLICE_X109Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y111_SLICE_X108Y111_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y111_SLICE_X108Y111_CO5),
.Q(CLBLM_L_X72Y111_SLICE_X108Y111_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y111_SLICE_X108Y111_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y111_SLICE_X108Y111_BO6),
.Q(CLBLM_L_X72Y111_SLICE_X108Y111_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y111_SLICE_X108Y111_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y111_SLICE_X108Y111_CO6),
.Q(CLBLM_L_X72Y111_SLICE_X108Y111_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y111_SLICE_X108Y111_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y111_SLICE_X108Y111_DO6),
.Q(CLBLM_L_X72Y111_SLICE_X108Y111_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0078cccc00f0cccc)
  ) CLBLM_L_X72Y111_SLICE_X108Y111_DLUT (
.I0(CLBLM_L_X72Y111_SLICE_X109Y111_AQ),
.I1(CLBLM_L_X72Y111_SLICE_X109Y111_A5Q),
.I2(CLBLM_L_X72Y111_SLICE_X108Y111_DQ),
.I3(CLBLM_L_X72Y111_SLICE_X109Y111_CQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X70Y111_SLICE_X104Y111_BQ),
.O5(CLBLM_L_X72Y111_SLICE_X108Y111_DO5),
.O6(CLBLM_L_X72Y111_SLICE_X108Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haf00aff00c0c0c0c)
  ) CLBLM_L_X72Y111_SLICE_X108Y111_CLUT (
.I0(CLBLM_L_X72Y109_SLICE_X108Y109_AO6),
.I1(CLBLM_L_X78Y123_SLICE_X121Y123_A5Q),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X70Y112_SLICE_X104Y112_CQ),
.I4(CLBLL_R_X71Y111_SLICE_X107Y111_CO6),
.I5(1'b1),
.O5(CLBLM_L_X72Y111_SLICE_X108Y111_CO5),
.O6(CLBLM_L_X72Y111_SLICE_X108Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8888f5f5a0a0)
  ) CLBLM_L_X72Y111_SLICE_X108Y111_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X72Y111_SLICE_X108Y111_BQ),
.I2(CLBLM_L_X72Y109_SLICE_X108Y109_AO6),
.I3(1'b1),
.I4(CLBLM_L_X72Y111_SLICE_X108Y111_CQ),
.I5(CLBLM_L_X70Y112_SLICE_X104Y112_CQ),
.O5(CLBLM_L_X72Y111_SLICE_X108Y111_BO5),
.O6(CLBLM_L_X72Y111_SLICE_X108Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fffff50705050)
  ) CLBLM_L_X72Y111_SLICE_X108Y111_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X72Y111_SLICE_X109Y111_CQ),
.I2(CLBLM_L_X72Y111_SLICE_X108Y111_DQ),
.I3(CLBLM_L_X70Y111_SLICE_X104Y111_BQ),
.I4(CLBLM_L_X72Y111_SLICE_X109Y111_AQ),
.I5(1'b1),
.O5(CLBLM_L_X72Y111_SLICE_X108Y111_AO5),
.O6(CLBLM_L_X72Y111_SLICE_X108Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y111_SLICE_X109Y111_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y111_SLICE_X109Y111_AO5),
.Q(CLBLM_L_X72Y111_SLICE_X109Y111_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y111_SLICE_X109Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y111_SLICE_X109Y111_AO6),
.Q(CLBLM_L_X72Y111_SLICE_X109Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y111_SLICE_X109Y111_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y113_SLICE_X108Y113_BQ),
.Q(CLBLM_L_X72Y111_SLICE_X109Y111_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y111_SLICE_X109Y111_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y111_SLICE_X108Y111_AO5),
.Q(CLBLM_L_X72Y111_SLICE_X109Y111_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y111_SLICE_X109Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y111_SLICE_X109Y111_DO5),
.O6(CLBLM_L_X72Y111_SLICE_X109Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y111_SLICE_X109Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y111_SLICE_X109Y111_CO5),
.O6(CLBLM_L_X72Y111_SLICE_X109Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y111_SLICE_X109Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y111_SLICE_X109Y111_BO5),
.O6(CLBLM_L_X72Y111_SLICE_X109Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h446c446c507a50d0)
  ) CLBLM_L_X72Y111_SLICE_X109Y111_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X70Y111_SLICE_X104Y111_BQ),
.I2(CLBLM_L_X72Y111_SLICE_X109Y111_AQ),
.I3(CLBLM_L_X72Y111_SLICE_X109Y111_CQ),
.I4(CLBLM_L_X72Y111_SLICE_X109Y111_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X72Y111_SLICE_X109Y111_AO5),
.O6(CLBLM_L_X72Y111_SLICE_X109Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y113_SLICE_X108Y113_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y108_SLICE_X105Y108_AO5),
.Q(CLBLM_L_X72Y113_SLICE_X108Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y113_SLICE_X108Y113_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X70Y113_SLICE_X104Y113_CQ),
.Q(CLBLM_L_X72Y113_SLICE_X108Y113_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y113_SLICE_X108Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y113_SLICE_X108Y113_DO5),
.O6(CLBLM_L_X72Y113_SLICE_X108Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y113_SLICE_X108Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y113_SLICE_X108Y113_CO5),
.O6(CLBLM_L_X72Y113_SLICE_X108Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y113_SLICE_X108Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y113_SLICE_X108Y113_BO5),
.O6(CLBLM_L_X72Y113_SLICE_X108Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y113_SLICE_X108Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y113_SLICE_X108Y113_AO5),
.O6(CLBLM_L_X72Y113_SLICE_X108Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y113_SLICE_X109Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y113_SLICE_X109Y113_DO5),
.O6(CLBLM_L_X72Y113_SLICE_X109Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y113_SLICE_X109Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y113_SLICE_X109Y113_CO5),
.O6(CLBLM_L_X72Y113_SLICE_X109Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y113_SLICE_X109Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y113_SLICE_X109Y113_BO5),
.O6(CLBLM_L_X72Y113_SLICE_X109Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y113_SLICE_X109Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y113_SLICE_X109Y113_AO5),
.O6(CLBLM_L_X72Y113_SLICE_X109Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y116_SLICE_X108Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y116_SLICE_X108Y116_BQ),
.Q(CLBLM_L_X72Y116_SLICE_X108Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y116_SLICE_X108Y116_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y118_SLICE_X108Y118_BQ),
.Q(CLBLM_L_X72Y116_SLICE_X108Y116_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y116_SLICE_X108Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y116_SLICE_X108Y116_DO5),
.O6(CLBLM_L_X72Y116_SLICE_X108Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y116_SLICE_X108Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y116_SLICE_X108Y116_CO5),
.O6(CLBLM_L_X72Y116_SLICE_X108Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y116_SLICE_X108Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y116_SLICE_X108Y116_BO5),
.O6(CLBLM_L_X72Y116_SLICE_X108Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y116_SLICE_X108Y116_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y116_SLICE_X108Y116_AO5),
.O6(CLBLM_L_X72Y116_SLICE_X108Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y116_SLICE_X109Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y116_SLICE_X109Y116_DO5),
.O6(CLBLM_L_X72Y116_SLICE_X109Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y116_SLICE_X109Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y116_SLICE_X109Y116_CO5),
.O6(CLBLM_L_X72Y116_SLICE_X109Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y116_SLICE_X109Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y116_SLICE_X109Y116_BO5),
.O6(CLBLM_L_X72Y116_SLICE_X109Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y116_SLICE_X109Y116_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y116_SLICE_X109Y116_AO5),
.O6(CLBLM_L_X72Y116_SLICE_X109Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y117_SLICE_X108Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y118_SLICE_X108Y118_C5Q),
.Q(CLBLM_L_X72Y117_SLICE_X108Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y117_SLICE_X108Y117_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y117_SLICE_X108Y117_AQ),
.Q(CLBLM_L_X72Y117_SLICE_X108Y117_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y117_SLICE_X108Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y117_SLICE_X108Y117_DO5),
.O6(CLBLM_L_X72Y117_SLICE_X108Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y117_SLICE_X108Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y117_SLICE_X108Y117_CO5),
.O6(CLBLM_L_X72Y117_SLICE_X108Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y117_SLICE_X108Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y117_SLICE_X108Y117_BO5),
.O6(CLBLM_L_X72Y117_SLICE_X108Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y117_SLICE_X108Y117_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y117_SLICE_X108Y117_AO5),
.O6(CLBLM_L_X72Y117_SLICE_X108Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y117_SLICE_X109Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y117_SLICE_X109Y117_DO5),
.O6(CLBLM_L_X72Y117_SLICE_X109Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y117_SLICE_X109Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y117_SLICE_X109Y117_CO5),
.O6(CLBLM_L_X72Y117_SLICE_X109Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y117_SLICE_X109Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y117_SLICE_X109Y117_BO5),
.O6(CLBLM_L_X72Y117_SLICE_X109Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y117_SLICE_X109Y117_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y117_SLICE_X109Y117_AO5),
.O6(CLBLM_L_X72Y117_SLICE_X109Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y118_SLICE_X108Y118_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y118_SLICE_X108Y118_AO5),
.Q(CLBLM_L_X72Y118_SLICE_X108Y118_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y118_SLICE_X108Y118_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y118_SLICE_X108Y118_BO5),
.Q(CLBLM_L_X72Y118_SLICE_X108Y118_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y118_SLICE_X108Y118_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y118_SLICE_X108Y118_CO5),
.Q(CLBLM_L_X72Y118_SLICE_X108Y118_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y118_SLICE_X108Y118_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y118_SLICE_X108Y118_DO5),
.Q(CLBLM_L_X72Y118_SLICE_X108Y118_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y118_SLICE_X108Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y118_SLICE_X108Y118_AO6),
.Q(CLBLM_L_X72Y118_SLICE_X108Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y118_SLICE_X108Y118_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y118_SLICE_X108Y118_BO6),
.Q(CLBLM_L_X72Y118_SLICE_X108Y118_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y118_SLICE_X108Y118_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y118_SLICE_X108Y118_CO6),
.Q(CLBLM_L_X72Y118_SLICE_X108Y118_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y118_SLICE_X108Y118_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y118_SLICE_X108Y118_DO6),
.Q(CLBLM_L_X72Y118_SLICE_X108Y118_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55f0fff0cc00cc00)
  ) CLBLM_L_X72Y118_SLICE_X108Y118_DLUT (
.I0(CLBLM_L_X72Y117_SLICE_X108Y117_BQ),
.I1(CLBLM_L_X70Y104_SLICE_X104Y104_A5Q),
.I2(CLBLM_L_X74Y118_SLICE_X112Y118_CQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X72Y117_SLICE_X108Y117_AQ),
.I5(1'b1),
.O5(CLBLM_L_X72Y118_SLICE_X108Y118_DO5),
.O6(CLBLM_L_X72Y118_SLICE_X108Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0fff0fafffa00)
  ) CLBLM_L_X72Y118_SLICE_X108Y118_CLUT (
.I0(CLBLM_L_X72Y118_SLICE_X108Y118_C5Q),
.I1(1'b1),
.I2(CLBLM_L_X74Y119_SLICE_X112Y119_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X72Y118_SLICE_X108Y118_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X72Y118_SLICE_X108Y118_CO5),
.O6(CLBLM_L_X72Y118_SLICE_X108Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00cc00fa00fa00)
  ) CLBLM_L_X72Y118_SLICE_X108Y118_BLUT (
.I0(CLBLM_L_X72Y118_SLICE_X108Y118_B5Q),
.I1(CLBLM_L_X72Y118_SLICE_X108Y118_BQ),
.I2(CLBLM_L_X72Y118_SLICE_X108Y118_DQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLL_R_X71Y119_SLICE_X106Y119_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X72Y118_SLICE_X108Y118_BO5),
.O6(CLBLM_L_X72Y118_SLICE_X108Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcaaaa0000cccc)
  ) CLBLM_L_X72Y118_SLICE_X108Y118_ALUT (
.I0(CLBLM_L_X72Y121_SLICE_X109Y121_A5Q),
.I1(CLBLM_L_X72Y118_SLICE_X108Y118_DQ),
.I2(CLBLM_L_X72Y118_SLICE_X108Y118_AQ),
.I3(CLBLM_L_X74Y119_SLICE_X112Y119_AQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLM_L_X72Y118_SLICE_X108Y118_AO5),
.O6(CLBLM_L_X72Y118_SLICE_X108Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y118_SLICE_X109Y118_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y118_SLICE_X109Y118_AO5),
.Q(CLBLM_L_X72Y118_SLICE_X109Y118_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y118_SLICE_X109Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y118_SLICE_X109Y118_AO6),
.Q(CLBLM_L_X72Y118_SLICE_X109Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y118_SLICE_X109Y118_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y118_SLICE_X109Y118_BO6),
.Q(CLBLM_L_X72Y118_SLICE_X109Y118_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y118_SLICE_X109Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y118_SLICE_X109Y118_DO5),
.O6(CLBLM_L_X72Y118_SLICE_X109Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y118_SLICE_X109Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y118_SLICE_X109Y118_CO5),
.O6(CLBLM_L_X72Y118_SLICE_X109Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3fffff3fc0f0f0c0)
  ) CLBLM_L_X72Y118_SLICE_X109Y118_BLUT (
.I0(1'b1),
.I1(CLBLL_R_X73Y118_SLICE_X110Y118_AQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X72Y119_SLICE_X108Y119_BQ),
.I4(CLBLL_R_X73Y118_SLICE_X110Y118_BQ),
.I5(CLBLM_L_X72Y119_SLICE_X108Y119_A5Q),
.O5(CLBLM_L_X72Y118_SLICE_X109Y118_BO5),
.O6(CLBLM_L_X72Y118_SLICE_X109Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafffa00cc00cc00)
  ) CLBLM_L_X72Y118_SLICE_X109Y118_ALUT (
.I0(CLBLL_R_X83Y94_SLICE_X130Y94_AQ),
.I1(CLBLL_R_X73Y104_SLICE_X110Y104_BQ),
.I2(CLBLM_L_X72Y118_SLICE_X109Y118_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X72Y119_SLICE_X108Y119_AQ),
.I5(1'b1),
.O5(CLBLM_L_X72Y118_SLICE_X109Y118_AO5),
.O6(CLBLM_L_X72Y118_SLICE_X109Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y119_SLICE_X108Y119_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y119_SLICE_X108Y119_AO5),
.Q(CLBLM_L_X72Y119_SLICE_X108Y119_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y119_SLICE_X108Y119_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y119_SLICE_X108Y119_CO5),
.Q(CLBLM_L_X72Y119_SLICE_X108Y119_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y119_SLICE_X108Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y119_SLICE_X108Y119_AO6),
.Q(CLBLM_L_X72Y119_SLICE_X108Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y119_SLICE_X108Y119_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y119_SLICE_X108Y119_BO6),
.Q(CLBLM_L_X72Y119_SLICE_X108Y119_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y119_SLICE_X108Y119_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y119_SLICE_X108Y119_CO6),
.Q(CLBLM_L_X72Y119_SLICE_X108Y119_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000100000000)
  ) CLBLM_L_X72Y119_SLICE_X108Y119_DLUT (
.I0(CLBLM_L_X72Y119_SLICE_X109Y119_A5Q),
.I1(CLBLM_L_X72Y119_SLICE_X108Y119_CQ),
.I2(CLBLM_L_X72Y119_SLICE_X109Y119_B5Q),
.I3(CLBLM_L_X70Y119_SLICE_X105Y119_A5Q),
.I4(CLBLM_L_X72Y119_SLICE_X109Y119_BQ),
.I5(CLBLL_R_X73Y118_SLICE_X111Y118_A5Q),
.O5(CLBLM_L_X72Y119_SLICE_X108Y119_DO5),
.O6(CLBLM_L_X72Y119_SLICE_X108Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc88ccf000f000)
  ) CLBLM_L_X72Y119_SLICE_X108Y119_CLUT (
.I0(CLBLM_L_X72Y119_SLICE_X109Y119_AQ),
.I1(CLBLM_L_X70Y119_SLICE_X105Y119_A5Q),
.I2(CLBLM_L_X68Y101_SLICE_X102Y101_BQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X72Y119_SLICE_X108Y119_DO6),
.I5(1'b1),
.O5(CLBLM_L_X72Y119_SLICE_X108Y119_CO5),
.O6(CLBLM_L_X72Y119_SLICE_X108Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccfcccccccccccc)
  ) CLBLM_L_X72Y119_SLICE_X108Y119_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X72Y119_SLICE_X109Y119_B5Q),
.I2(CLBLM_L_X72Y119_SLICE_X109Y119_CO6),
.I3(CLBLL_R_X73Y118_SLICE_X111Y118_A5Q),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X72Y119_SLICE_X108Y119_A5Q),
.O5(CLBLM_L_X72Y119_SLICE_X108Y119_BO5),
.O6(CLBLM_L_X72Y119_SLICE_X108Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff00f8f8cccc)
  ) CLBLM_L_X72Y119_SLICE_X108Y119_ALUT (
.I0(CLBLM_L_X72Y119_SLICE_X108Y119_DO6),
.I1(CLBLM_L_X72Y119_SLICE_X108Y119_BQ),
.I2(CLBLM_L_X72Y119_SLICE_X109Y119_A5Q),
.I3(CLBLL_R_X71Y124_SLICE_X106Y124_BQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLM_L_X72Y119_SLICE_X108Y119_AO5),
.O6(CLBLM_L_X72Y119_SLICE_X108Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y119_SLICE_X109Y119_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y119_SLICE_X108Y119_CQ),
.Q(CLBLM_L_X72Y119_SLICE_X109Y119_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y119_SLICE_X109Y119_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y119_SLICE_X109Y119_BQ),
.Q(CLBLM_L_X72Y119_SLICE_X109Y119_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y119_SLICE_X109Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y119_SLICE_X109Y119_AO6),
.Q(CLBLM_L_X72Y119_SLICE_X109Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y119_SLICE_X109Y119_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y119_SLICE_X109Y119_BO6),
.Q(CLBLM_L_X72Y119_SLICE_X109Y119_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000003300000033)
  ) CLBLM_L_X72Y119_SLICE_X109Y119_DLUT (
.I0(1'b1),
.I1(CLBLL_R_X73Y118_SLICE_X111Y118_A5Q),
.I2(1'b1),
.I3(CLBLL_R_X73Y119_SLICE_X110Y119_B5Q),
.I4(CLBLL_R_X73Y119_SLICE_X110Y119_CO6),
.I5(1'b1),
.O5(CLBLM_L_X72Y119_SLICE_X109Y119_DO5),
.O6(CLBLM_L_X72Y119_SLICE_X109Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffefffffffe)
  ) CLBLM_L_X72Y119_SLICE_X109Y119_CLUT (
.I0(CLBLM_L_X72Y119_SLICE_X109Y119_A5Q),
.I1(CLBLM_L_X70Y119_SLICE_X105Y119_A5Q),
.I2(CLBLM_L_X72Y119_SLICE_X109Y119_BQ),
.I3(CLBLM_L_X72Y119_SLICE_X108Y119_CQ),
.I4(CLBLM_L_X72Y119_SLICE_X109Y119_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X72Y119_SLICE_X109Y119_CO5),
.O6(CLBLM_L_X72Y119_SLICE_X109Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0aff3bff0a003b00)
  ) CLBLM_L_X72Y119_SLICE_X109Y119_BLUT (
.I0(CLBLM_L_X70Y119_SLICE_X105Y119_A5Q),
.I1(CLBLL_R_X73Y118_SLICE_X111Y118_A5Q),
.I2(CLBLM_L_X72Y119_SLICE_X109Y119_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X72Y119_SLICE_X109Y119_CO6),
.I5(CLBLM_L_X72Y119_SLICE_X109Y119_A5Q),
.O5(CLBLM_L_X72Y119_SLICE_X109Y119_BO5),
.O6(CLBLM_L_X72Y119_SLICE_X109Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff3bcc08ffb3cc80)
  ) CLBLM_L_X72Y119_SLICE_X109Y119_ALUT (
.I0(CLBLL_R_X73Y119_SLICE_X110Y119_CO6),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_L_X72Y119_SLICE_X109Y119_AQ),
.I3(CLBLM_L_X72Y119_SLICE_X109Y119_DO6),
.I4(CLBLL_R_X73Y118_SLICE_X110Y118_AQ),
.I5(CLBLM_L_X72Y113_SLICE_X108Y113_AQ),
.O5(CLBLM_L_X72Y119_SLICE_X109Y119_AO5),
.O6(CLBLM_L_X72Y119_SLICE_X109Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y120_SLICE_X108Y120_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y120_SLICE_X108Y120_AO5),
.Q(CLBLM_L_X72Y120_SLICE_X108Y120_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y120_SLICE_X108Y120_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y120_SLICE_X108Y120_AO6),
.Q(CLBLM_L_X72Y120_SLICE_X108Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y120_SLICE_X108Y120_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y120_SLICE_X108Y120_BO6),
.Q(CLBLM_L_X72Y120_SLICE_X108Y120_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y120_SLICE_X108Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y120_SLICE_X108Y120_DO5),
.O6(CLBLM_L_X72Y120_SLICE_X108Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y120_SLICE_X108Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y120_SLICE_X108Y120_CO5),
.O6(CLBLM_L_X72Y120_SLICE_X108Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333333333333)
  ) CLBLM_L_X72Y120_SLICE_X108Y120_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X72Y120_SLICE_X108Y120_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y120_SLICE_X108Y120_BO5),
.O6(CLBLM_L_X72Y120_SLICE_X108Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfffc00bbf0bbf0)
  ) CLBLM_L_X72Y120_SLICE_X108Y120_ALUT (
.I0(CLBLM_L_X72Y120_SLICE_X108Y120_A5Q),
.I1(CLBLM_L_X72Y120_SLICE_X108Y120_BQ),
.I2(CLBLM_L_X72Y120_SLICE_X108Y120_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X72Y118_SLICE_X109Y118_AQ),
.I5(1'b1),
.O5(CLBLM_L_X72Y120_SLICE_X108Y120_AO5),
.O6(CLBLM_L_X72Y120_SLICE_X108Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y120_SLICE_X109Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y120_SLICE_X109Y120_DO5),
.O6(CLBLM_L_X72Y120_SLICE_X109Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y120_SLICE_X109Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y120_SLICE_X109Y120_CO5),
.O6(CLBLM_L_X72Y120_SLICE_X109Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y120_SLICE_X109Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y120_SLICE_X109Y120_BO5),
.O6(CLBLM_L_X72Y120_SLICE_X109Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y120_SLICE_X109Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y120_SLICE_X109Y120_AO5),
.O6(CLBLM_L_X72Y120_SLICE_X109Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y121_SLICE_X108Y121_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y121_SLICE_X108Y121_DQ),
.Q(CLBLM_L_X72Y121_SLICE_X108Y121_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y121_SLICE_X108Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y121_SLICE_X108Y121_AO5),
.Q(CLBLM_L_X72Y121_SLICE_X108Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y121_SLICE_X108Y121_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y120_SLICE_X108Y120_A5Q),
.Q(CLBLM_L_X72Y121_SLICE_X108Y121_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y121_SLICE_X108Y121_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y121_SLICE_X108Y121_BQ),
.Q(CLBLM_L_X72Y121_SLICE_X108Y121_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y121_SLICE_X108Y121_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y121_SLICE_X108Y121_CQ),
.Q(CLBLM_L_X72Y121_SLICE_X108Y121_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y121_SLICE_X108Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y121_SLICE_X108Y121_DO5),
.O6(CLBLM_L_X72Y121_SLICE_X108Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y121_SLICE_X108Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y121_SLICE_X108Y121_CO5),
.O6(CLBLM_L_X72Y121_SLICE_X108Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0015003f15153f3f)
  ) CLBLM_L_X72Y121_SLICE_X108Y121_BLUT (
.I0(CLBLM_L_X72Y122_SLICE_X108Y122_CQ),
.I1(CLBLM_L_X72Y121_SLICE_X108Y121_BQ),
.I2(CLBLM_L_X74Y122_SLICE_X112Y122_BQ),
.I3(CLBLM_L_X72Y118_SLICE_X108Y118_AQ),
.I4(CLBLM_L_X72Y128_SLICE_X109Y128_AQ),
.I5(CLBLM_L_X72Y121_SLICE_X108Y121_A5Q),
.O5(CLBLM_L_X72Y121_SLICE_X108Y121_BO5),
.O6(CLBLM_L_X72Y121_SLICE_X108Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeaacc00f0f0f0f0)
  ) CLBLM_L_X72Y121_SLICE_X108Y121_ALUT (
.I0(CLBLM_L_X72Y121_SLICE_X108Y121_CQ),
.I1(CLBLM_L_X72Y121_SLICE_X108Y121_DQ),
.I2(CLBLM_L_X76Y119_SLICE_X116Y119_AQ),
.I3(CLBLM_L_X72Y121_SLICE_X109Y121_A5Q),
.I4(CLBLM_L_X72Y121_SLICE_X109Y121_AQ),
.I5(1'b1),
.O5(CLBLM_L_X72Y121_SLICE_X108Y121_AO5),
.O6(CLBLM_L_X72Y121_SLICE_X108Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y121_SLICE_X109Y121_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y121_SLICE_X109Y121_AO5),
.Q(CLBLM_L_X72Y121_SLICE_X109Y121_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y121_SLICE_X109Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y121_SLICE_X109Y121_AO6),
.Q(CLBLM_L_X72Y121_SLICE_X109Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y121_SLICE_X109Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y121_SLICE_X109Y121_DO5),
.O6(CLBLM_L_X72Y121_SLICE_X109Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y121_SLICE_X109Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y121_SLICE_X109Y121_CO5),
.O6(CLBLM_L_X72Y121_SLICE_X109Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y121_SLICE_X109Y121_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y121_SLICE_X109Y121_BO5),
.O6(CLBLM_L_X72Y121_SLICE_X109Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7ffc4ccfcfcfcfc)
  ) CLBLM_L_X72Y121_SLICE_X109Y121_ALUT (
.I0(CLBLM_L_X74Y129_SLICE_X113Y129_BO5),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_L_X72Y121_SLICE_X109Y121_AQ),
.I3(CLBLL_R_X73Y132_SLICE_X111Y132_AO6),
.I4(CLBLM_L_X74Y122_SLICE_X112Y122_BQ),
.I5(1'b1),
.O5(CLBLM_L_X72Y121_SLICE_X109Y121_AO5),
.O6(CLBLM_L_X72Y121_SLICE_X109Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y122_SLICE_X108Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y121_SLICE_X108Y121_A5Q),
.Q(CLBLM_L_X72Y122_SLICE_X108Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y122_SLICE_X108Y122_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y122_SLICE_X108Y122_AQ),
.Q(CLBLM_L_X72Y122_SLICE_X108Y122_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y122_SLICE_X108Y122_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y122_SLICE_X108Y122_BQ),
.Q(CLBLM_L_X72Y122_SLICE_X108Y122_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y122_SLICE_X108Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y122_SLICE_X108Y122_DO5),
.O6(CLBLM_L_X72Y122_SLICE_X108Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y122_SLICE_X108Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y122_SLICE_X108Y122_CO5),
.O6(CLBLM_L_X72Y122_SLICE_X108Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y122_SLICE_X108Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y122_SLICE_X108Y122_BO5),
.O6(CLBLM_L_X72Y122_SLICE_X108Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000070007000700)
  ) CLBLM_L_X72Y122_SLICE_X108Y122_ALUT (
.I0(CLBLM_L_X72Y122_SLICE_X108Y122_BQ),
.I1(CLBLM_L_X72Y123_SLICE_X108Y123_BQ),
.I2(CLBLM_L_X72Y121_SLICE_X108Y121_AO6),
.I3(CLBLM_L_X72Y121_SLICE_X108Y121_BO6),
.I4(CLBLL_R_X71Y121_SLICE_X106Y121_AQ),
.I5(CLBLM_L_X72Y122_SLICE_X108Y122_AQ),
.O5(CLBLM_L_X72Y122_SLICE_X108Y122_AO5),
.O6(CLBLM_L_X72Y122_SLICE_X108Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y122_SLICE_X109Y122_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y122_SLICE_X109Y122_CO5),
.Q(CLBLM_L_X72Y122_SLICE_X109Y122_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y122_SLICE_X109Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y122_SLICE_X109Y122_AO6),
.Q(CLBLM_L_X72Y122_SLICE_X109Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y122_SLICE_X109Y122_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y122_SLICE_X109Y122_BO6),
.Q(CLBLM_L_X72Y122_SLICE_X109Y122_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y122_SLICE_X109Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y122_SLICE_X109Y122_DO5),
.O6(CLBLM_L_X72Y122_SLICE_X109Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fff0ff7d5a280)
  ) CLBLM_L_X72Y122_SLICE_X109Y122_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X71Y124_SLICE_X106Y124_CO6),
.I2(CLBLL_R_X73Y123_SLICE_X111Y123_AQ),
.I3(CLBLM_L_X72Y122_SLICE_X109Y122_A5Q),
.I4(CLBLL_R_X73Y123_SLICE_X110Y123_CQ),
.I5(1'b1),
.O5(CLBLM_L_X72Y122_SLICE_X109Y122_CO5),
.O6(CLBLM_L_X72Y122_SLICE_X109Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0f044eef0f0)
  ) CLBLM_L_X72Y122_SLICE_X109Y122_BLUT (
.I0(CLBLL_R_X71Y124_SLICE_X106Y124_CO6),
.I1(CLBLM_L_X72Y122_SLICE_X109Y122_BQ),
.I2(CLBLL_R_X73Y121_SLICE_X111Y121_AQ),
.I3(CLBLL_R_X73Y122_SLICE_X111Y122_AO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X72Y122_SLICE_X109Y122_CO6),
.O5(CLBLM_L_X72Y122_SLICE_X109Y122_BO5),
.O6(CLBLM_L_X72Y122_SLICE_X109Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5050ccccf0facccc)
  ) CLBLM_L_X72Y122_SLICE_X109Y122_ALUT (
.I0(CLBLL_R_X71Y124_SLICE_X106Y124_CO6),
.I1(CLBLM_L_X72Y122_SLICE_X109Y122_BQ),
.I2(CLBLM_L_X72Y122_SLICE_X109Y122_AQ),
.I3(CLBLL_R_X73Y123_SLICE_X111Y123_AQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X72Y122_SLICE_X109Y122_A5Q),
.O5(CLBLM_L_X72Y122_SLICE_X109Y122_AO5),
.O6(CLBLM_L_X72Y122_SLICE_X109Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y123_SLICE_X108Y123_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y123_SLICE_X108Y123_BO5),
.Q(CLBLM_L_X72Y123_SLICE_X108Y123_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y123_SLICE_X108Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y123_SLICE_X108Y123_AO6),
.Q(CLBLM_L_X72Y123_SLICE_X108Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y123_SLICE_X108Y123_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y123_SLICE_X108Y123_CO5),
.Q(CLBLM_L_X72Y123_SLICE_X108Y123_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y123_SLICE_X108Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y123_SLICE_X108Y123_DO5),
.O6(CLBLM_L_X72Y123_SLICE_X108Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffcceeffffaaaa)
  ) CLBLM_L_X72Y123_SLICE_X108Y123_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X71Y129_SLICE_X107Y129_AO6),
.I2(1'b1),
.I3(CLBLM_L_X72Y125_SLICE_X109Y125_CO6),
.I4(CLBLL_R_X71Y121_SLICE_X106Y121_AQ),
.I5(1'b1),
.O5(CLBLM_L_X72Y123_SLICE_X108Y123_CO5),
.O6(CLBLM_L_X72Y123_SLICE_X108Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ff55fcfcacfc)
  ) CLBLM_L_X72Y123_SLICE_X108Y123_BLUT (
.I0(CLBLL_R_X71Y129_SLICE_X107Y129_AO6),
.I1(CLBLL_R_X71Y121_SLICE_X106Y121_A5Q),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X72Y125_SLICE_X109Y125_CO6),
.I4(CLBLM_L_X72Y123_SLICE_X108Y123_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X72Y123_SLICE_X108Y123_BO5),
.O6(CLBLM_L_X72Y123_SLICE_X108Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaccccf0f0cccc)
  ) CLBLM_L_X72Y123_SLICE_X108Y123_ALUT (
.I0(CLBLL_R_X73Y121_SLICE_X110Y121_CO6),
.I1(CLBLM_L_X72Y122_SLICE_X109Y122_A5Q),
.I2(CLBLM_L_X72Y123_SLICE_X108Y123_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X71Y124_SLICE_X106Y124_CO6),
.O5(CLBLM_L_X72Y123_SLICE_X108Y123_AO5),
.O6(CLBLM_L_X72Y123_SLICE_X108Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y123_SLICE_X109Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y123_SLICE_X109Y123_AO6),
.Q(CLBLM_L_X72Y123_SLICE_X109Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y123_SLICE_X109Y123_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y123_SLICE_X109Y123_BO6),
.Q(CLBLM_L_X72Y123_SLICE_X109Y123_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y123_SLICE_X109Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y123_SLICE_X109Y123_DO5),
.O6(CLBLM_L_X72Y123_SLICE_X109Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc0000000000)
  ) CLBLM_L_X72Y123_SLICE_X109Y123_CLUT (
.I0(1'b1),
.I1(CLBLL_R_X71Y124_SLICE_X106Y124_CO6),
.I2(1'b1),
.I3(CLBLM_L_X72Y122_SLICE_X109Y122_AQ),
.I4(1'b1),
.I5(CLBLM_L_X72Y122_SLICE_X109Y122_A5Q),
.O5(CLBLM_L_X72Y123_SLICE_X109Y123_CO5),
.O6(CLBLM_L_X72Y123_SLICE_X109Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a5f0f0ccccf0f0)
  ) CLBLM_L_X72Y123_SLICE_X109Y123_BLUT (
.I0(CLBLL_R_X73Y123_SLICE_X111Y123_DQ),
.I1(CLBLM_L_X72Y123_SLICE_X109Y123_BQ),
.I2(CLBLM_L_X72Y123_SLICE_X109Y123_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X72Y123_SLICE_X109Y123_CO6),
.O5(CLBLM_L_X72Y123_SLICE_X109Y123_BO5),
.O6(CLBLM_L_X72Y123_SLICE_X109Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8f0aaaaf0f0aaaa)
  ) CLBLM_L_X72Y123_SLICE_X109Y123_ALUT (
.I0(CLBLL_R_X73Y123_SLICE_X111Y123_DQ),
.I1(CLBLL_R_X71Y124_SLICE_X106Y124_CO6),
.I2(CLBLM_L_X72Y123_SLICE_X109Y123_AQ),
.I3(CLBLM_L_X72Y122_SLICE_X109Y122_A5Q),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X72Y122_SLICE_X109Y122_AQ),
.O5(CLBLM_L_X72Y123_SLICE_X109Y123_AO5),
.O6(CLBLM_L_X72Y123_SLICE_X109Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y124_SLICE_X108Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y124_SLICE_X108Y124_AO6),
.Q(CLBLM_L_X72Y124_SLICE_X108Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y124_SLICE_X108Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y124_SLICE_X108Y124_DO5),
.O6(CLBLM_L_X72Y124_SLICE_X108Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y124_SLICE_X108Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y124_SLICE_X108Y124_CO5),
.O6(CLBLM_L_X72Y124_SLICE_X108Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0003000200030003)
  ) CLBLM_L_X72Y124_SLICE_X108Y124_BLUT (
.I0(CLBLL_R_X71Y126_SLICE_X107Y126_BQ),
.I1(CLBLM_L_X70Y124_SLICE_X105Y124_BO6),
.I2(CLBLL_R_X71Y126_SLICE_X107Y126_AQ),
.I3(CLBLM_L_X70Y125_SLICE_X105Y125_AQ),
.I4(CLBLM_L_X70Y123_SLICE_X104Y123_AQ),
.I5(CLBLM_L_X70Y124_SLICE_X104Y124_BQ),
.O5(CLBLM_L_X72Y124_SLICE_X108Y124_BO5),
.O6(CLBLM_L_X72Y124_SLICE_X108Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3ff3bff3c0c040c0)
  ) CLBLM_L_X72Y124_SLICE_X108Y124_ALUT (
.I0(CLBLL_R_X73Y124_SLICE_X110Y124_A5Q),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_L_X72Y124_SLICE_X108Y124_AQ),
.I3(CLBLM_L_X72Y124_SLICE_X108Y124_BO6),
.I4(CLBLM_L_X72Y124_SLICE_X109Y124_AQ),
.I5(CLBLM_L_X72Y125_SLICE_X108Y125_AQ),
.O5(CLBLM_L_X72Y124_SLICE_X108Y124_AO5),
.O6(CLBLM_L_X72Y124_SLICE_X108Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y124_SLICE_X109Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y124_SLICE_X109Y124_AO6),
.Q(CLBLM_L_X72Y124_SLICE_X109Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y124_SLICE_X109Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y124_SLICE_X109Y124_DO5),
.O6(CLBLM_L_X72Y124_SLICE_X109Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y124_SLICE_X109Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y124_SLICE_X109Y124_CO5),
.O6(CLBLM_L_X72Y124_SLICE_X109Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y124_SLICE_X109Y124_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y124_SLICE_X109Y124_BO5),
.O6(CLBLM_L_X72Y124_SLICE_X109Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3030ff00f4f4ff00)
  ) CLBLM_L_X72Y124_SLICE_X109Y124_ALUT (
.I0(CLBLL_R_X73Y124_SLICE_X110Y124_A5Q),
.I1(CLBLM_L_X72Y124_SLICE_X108Y124_BO6),
.I2(CLBLM_L_X72Y124_SLICE_X109Y124_AQ),
.I3(CLBLL_R_X73Y124_SLICE_X110Y124_AQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X73Y124_SLICE_X110Y124_BQ),
.O5(CLBLM_L_X72Y124_SLICE_X109Y124_AO5),
.O6(CLBLM_L_X72Y124_SLICE_X109Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y125_SLICE_X108Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y125_SLICE_X108Y125_AO6),
.Q(CLBLM_L_X72Y125_SLICE_X108Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y125_SLICE_X108Y125_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y125_SLICE_X108Y125_BO6),
.Q(CLBLM_L_X72Y125_SLICE_X108Y125_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y125_SLICE_X108Y125_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y125_SLICE_X108Y125_CO6),
.Q(CLBLM_L_X72Y125_SLICE_X108Y125_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0000000000)
  ) CLBLM_L_X72Y125_SLICE_X108Y125_DLUT (
.I0(CLBLM_L_X72Y124_SLICE_X109Y124_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_R_X73Y124_SLICE_X110Y124_BQ),
.I4(1'b1),
.I5(CLBLM_L_X72Y124_SLICE_X108Y124_BO6),
.O5(CLBLM_L_X72Y125_SLICE_X108Y125_DO5),
.O6(CLBLM_L_X72Y125_SLICE_X108Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf05ad8d8f05ad8d8)
  ) CLBLM_L_X72Y125_SLICE_X108Y125_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X72Y125_SLICE_X108Y125_CQ),
.I2(CLBLM_L_X72Y125_SLICE_X108Y125_BQ),
.I3(CLBLL_R_X73Y125_SLICE_X111Y125_DQ),
.I4(CLBLM_L_X72Y125_SLICE_X108Y125_DO6),
.I5(1'b1),
.O5(CLBLM_L_X72Y125_SLICE_X108Y125_CO5),
.O6(CLBLM_L_X72Y125_SLICE_X108Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hacaaccaaccaaccaa)
  ) CLBLM_L_X72Y125_SLICE_X108Y125_BLUT (
.I0(CLBLL_R_X73Y125_SLICE_X111Y125_DQ),
.I1(CLBLM_L_X72Y125_SLICE_X108Y125_BQ),
.I2(CLBLM_L_X72Y124_SLICE_X109Y124_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X72Y124_SLICE_X108Y124_BO6),
.I5(CLBLL_R_X73Y124_SLICE_X110Y124_BQ),
.O5(CLBLM_L_X72Y125_SLICE_X108Y125_BO5),
.O6(CLBLM_L_X72Y125_SLICE_X108Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfff0ffcc00f000)
  ) CLBLM_L_X72Y125_SLICE_X108Y125_ALUT (
.I0(1'b1),
.I1(CLBLL_R_X73Y125_SLICE_X110Y125_AO6),
.I2(CLBLM_L_X72Y125_SLICE_X108Y125_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X72Y124_SLICE_X108Y124_BO6),
.I5(CLBLL_R_X73Y124_SLICE_X110Y124_BQ),
.O5(CLBLM_L_X72Y125_SLICE_X108Y125_AO5),
.O6(CLBLM_L_X72Y125_SLICE_X108Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y125_SLICE_X109Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y125_SLICE_X109Y125_AO6),
.Q(CLBLM_L_X72Y125_SLICE_X109Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y125_SLICE_X109Y125_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y125_SLICE_X109Y125_BO6),
.Q(CLBLM_L_X72Y125_SLICE_X109Y125_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffeeffee)
  ) CLBLM_L_X72Y125_SLICE_X109Y125_DLUT (
.I0(CLBLM_L_X72Y123_SLICE_X109Y123_BQ),
.I1(CLBLM_L_X72Y126_SLICE_X109Y126_CQ),
.I2(1'b1),
.I3(CLBLM_L_X72Y125_SLICE_X108Y125_CQ),
.I4(1'b1),
.I5(CLBLL_R_X73Y125_SLICE_X111Y125_CQ),
.O5(CLBLM_L_X72Y125_SLICE_X109Y125_DO5),
.O6(CLBLM_L_X72Y125_SLICE_X109Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000003)
  ) CLBLM_L_X72Y125_SLICE_X109Y125_CLUT (
.I0(1'b1),
.I1(CLBLL_R_X73Y128_SLICE_X111Y128_BQ),
.I2(CLBLL_R_X75Y127_SLICE_X115Y127_CQ),
.I3(CLBLL_R_X73Y122_SLICE_X111Y122_DQ),
.I4(CLBLM_L_X72Y125_SLICE_X109Y125_DO6),
.I5(CLBLM_L_X72Y126_SLICE_X108Y126_BQ),
.O5(CLBLM_L_X72Y125_SLICE_X109Y125_CO5),
.O6(CLBLM_L_X72Y125_SLICE_X109Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cccaaaaccccaaaa)
  ) CLBLM_L_X72Y125_SLICE_X109Y125_BLUT (
.I0(CLBLM_L_X72Y125_SLICE_X109Y125_AQ),
.I1(CLBLM_L_X72Y125_SLICE_X109Y125_BQ),
.I2(CLBLM_L_X72Y124_SLICE_X109Y124_AQ),
.I3(CLBLM_L_X72Y124_SLICE_X108Y124_BO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X73Y124_SLICE_X110Y124_BQ),
.O5(CLBLM_L_X72Y125_SLICE_X109Y125_BO5),
.O6(CLBLM_L_X72Y125_SLICE_X109Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3accccca3accccc)
  ) CLBLM_L_X72Y125_SLICE_X109Y125_ALUT (
.I0(CLBLM_L_X72Y125_SLICE_X109Y125_AQ),
.I1(CLBLM_L_X72Y124_SLICE_X108Y124_AQ),
.I2(CLBLL_R_X73Y124_SLICE_X110Y124_CO5),
.I3(CLBLM_L_X74Y126_SLICE_X113Y126_CQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLM_L_X72Y125_SLICE_X109Y125_AO5),
.O6(CLBLM_L_X72Y125_SLICE_X109Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y126_SLICE_X108Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y126_SLICE_X108Y126_AO6),
.Q(CLBLM_L_X72Y126_SLICE_X108Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y126_SLICE_X108Y126_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y126_SLICE_X108Y126_BO6),
.Q(CLBLM_L_X72Y126_SLICE_X108Y126_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800880088008800)
  ) CLBLM_L_X72Y126_SLICE_X108Y126_DLUT (
.I0(CLBLM_L_X72Y127_SLICE_X108Y127_AQ),
.I1(CLBLM_L_X72Y127_SLICE_X108Y127_A5Q),
.I2(1'b1),
.I3(CLBLM_L_X72Y126_SLICE_X108Y126_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y126_SLICE_X108Y126_DO5),
.O6(CLBLM_L_X72Y126_SLICE_X108Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000e000f000)
  ) CLBLM_L_X72Y126_SLICE_X108Y126_CLUT (
.I0(CLBLM_L_X70Y123_SLICE_X104Y123_AQ),
.I1(CLBLL_R_X71Y126_SLICE_X107Y126_BQ),
.I2(CLBLL_R_X71Y126_SLICE_X107Y126_AQ),
.I3(CLBLM_L_X70Y125_SLICE_X105Y125_AQ),
.I4(CLBLL_R_X71Y126_SLICE_X106Y126_AQ),
.I5(CLBLM_L_X70Y124_SLICE_X105Y124_BO6),
.O5(CLBLM_L_X72Y126_SLICE_X108Y126_CO5),
.O6(CLBLM_L_X72Y126_SLICE_X108Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he44ee44ef0f0f0f0)
  ) CLBLM_L_X72Y126_SLICE_X108Y126_BLUT (
.I0(CLBLM_L_X72Y126_SLICE_X108Y126_DO6),
.I1(CLBLM_L_X72Y126_SLICE_X108Y126_BQ),
.I2(CLBLM_L_X72Y126_SLICE_X108Y126_AQ),
.I3(CLBLL_R_X75Y127_SLICE_X115Y127_DQ),
.I4(1'b1),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X72Y126_SLICE_X108Y126_BO5),
.O6(CLBLM_L_X72Y126_SLICE_X108Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8aaf0aaf0aaf0aa)
  ) CLBLM_L_X72Y126_SLICE_X108Y126_ALUT (
.I0(CLBLL_R_X75Y127_SLICE_X115Y127_DQ),
.I1(CLBLM_L_X72Y126_SLICE_X108Y126_CO6),
.I2(CLBLM_L_X72Y126_SLICE_X108Y126_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X72Y127_SLICE_X108Y127_AQ),
.I5(CLBLM_L_X72Y127_SLICE_X108Y127_A5Q),
.O5(CLBLM_L_X72Y126_SLICE_X108Y126_AO5),
.O6(CLBLM_L_X72Y126_SLICE_X108Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y126_SLICE_X109Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y126_SLICE_X109Y126_AO6),
.Q(CLBLM_L_X72Y126_SLICE_X109Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y126_SLICE_X109Y126_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y126_SLICE_X109Y126_BO6),
.Q(CLBLM_L_X72Y126_SLICE_X109Y126_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y126_SLICE_X109Y126_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y126_SLICE_X109Y126_CO6),
.Q(CLBLM_L_X72Y126_SLICE_X109Y126_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000000000000)
  ) CLBLM_L_X72Y126_SLICE_X109Y126_DLUT (
.I0(CLBLL_R_X71Y126_SLICE_X106Y126_CO6),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X72Y126_SLICE_X109Y126_AQ),
.I5(CLBLL_R_X73Y126_SLICE_X110Y126_A5Q),
.O5(CLBLM_L_X72Y126_SLICE_X109Y126_DO5),
.O6(CLBLM_L_X72Y126_SLICE_X109Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00dd8855aadd88)
  ) CLBLM_L_X72Y126_SLICE_X109Y126_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X72Y126_SLICE_X109Y126_CQ),
.I2(1'b1),
.I3(CLBLM_L_X72Y126_SLICE_X109Y126_BQ),
.I4(CLBLM_L_X72Y126_SLICE_X109Y126_DO6),
.I5(CLBLL_R_X73Y128_SLICE_X110Y128_AQ),
.O5(CLBLM_L_X72Y126_SLICE_X109Y126_CO5),
.O6(CLBLM_L_X72Y126_SLICE_X109Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hec4cccccff00ff00)
  ) CLBLM_L_X72Y126_SLICE_X109Y126_BLUT (
.I0(CLBLL_R_X73Y126_SLICE_X110Y126_A5Q),
.I1(CLBLM_L_X72Y126_SLICE_X109Y126_BQ),
.I2(CLBLM_L_X72Y126_SLICE_X109Y126_AQ),
.I3(CLBLL_R_X73Y128_SLICE_X110Y128_AQ),
.I4(CLBLL_R_X71Y126_SLICE_X106Y126_CO6),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X72Y126_SLICE_X109Y126_BO5),
.O6(CLBLM_L_X72Y126_SLICE_X109Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h77ff44cc37330400)
  ) CLBLM_L_X72Y126_SLICE_X109Y126_ALUT (
.I0(CLBLL_R_X73Y126_SLICE_X110Y126_A5Q),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLL_R_X71Y127_SLICE_X107Y127_AQ),
.I3(CLBLL_R_X71Y126_SLICE_X106Y126_CO6),
.I4(CLBLL_R_X73Y126_SLICE_X110Y126_BQ),
.I5(CLBLM_L_X72Y126_SLICE_X109Y126_AQ),
.O5(CLBLM_L_X72Y126_SLICE_X109Y126_AO5),
.O6(CLBLM_L_X72Y126_SLICE_X109Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y127_SLICE_X108Y127_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y127_SLICE_X108Y127_BO5),
.Q(CLBLM_L_X72Y127_SLICE_X108Y127_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y127_SLICE_X108Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y127_SLICE_X108Y127_AO6),
.Q(CLBLM_L_X72Y127_SLICE_X108Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y127_SLICE_X108Y127_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y127_SLICE_X108Y127_CO6),
.Q(CLBLM_L_X72Y127_SLICE_X108Y127_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y127_SLICE_X108Y127_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y127_SLICE_X108Y127_DO6),
.Q(CLBLM_L_X72Y127_SLICE_X108Y127_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7df5f5f528a0a0a0)
  ) CLBLM_L_X72Y127_SLICE_X108Y127_DLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X72Y127_SLICE_X108Y127_AQ),
.I2(CLBLM_L_X72Y127_SLICE_X108Y127_DQ),
.I3(CLBLM_L_X72Y127_SLICE_X108Y127_A5Q),
.I4(CLBLM_L_X72Y126_SLICE_X108Y126_CO6),
.I5(CLBLM_L_X72Y128_SLICE_X108Y128_DQ),
.O5(CLBLM_L_X72Y127_SLICE_X108Y127_DO5),
.O6(CLBLM_L_X72Y127_SLICE_X108Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcff000c0cff00)
  ) CLBLM_L_X72Y127_SLICE_X108Y127_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X72Y127_SLICE_X108Y127_CQ),
.I2(CLBLM_L_X72Y126_SLICE_X108Y126_CO6),
.I3(CLBLM_L_X72Y127_SLICE_X108Y127_A5Q),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X74Y127_SLICE_X112Y127_BO6),
.O5(CLBLM_L_X72Y127_SLICE_X108Y127_CO5),
.O6(CLBLM_L_X72Y127_SLICE_X108Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5555bf8cb380)
  ) CLBLM_L_X72Y127_SLICE_X108Y127_BLUT (
.I0(CLBLM_L_X72Y128_SLICE_X108Y128_A5Q),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_L_X72Y126_SLICE_X108Y126_CO6),
.I3(CLBLM_L_X72Y127_SLICE_X109Y127_BQ),
.I4(CLBLM_L_X72Y127_SLICE_X108Y127_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X72Y127_SLICE_X108Y127_BO5),
.O6(CLBLM_L_X72Y127_SLICE_X108Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h75752020f5fda0a8)
  ) CLBLM_L_X72Y127_SLICE_X108Y127_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X72Y126_SLICE_X108Y126_CO6),
.I2(CLBLM_L_X72Y127_SLICE_X108Y127_AQ),
.I3(CLBLM_L_X72Y128_SLICE_X108Y128_A5Q),
.I4(CLBLM_L_X72Y128_SLICE_X108Y128_AQ),
.I5(CLBLM_L_X72Y127_SLICE_X108Y127_A5Q),
.O5(CLBLM_L_X72Y127_SLICE_X108Y127_AO5),
.O6(CLBLM_L_X72Y127_SLICE_X108Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y127_SLICE_X109Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y127_SLICE_X114Y127_AQ),
.Q(CLBLM_L_X72Y127_SLICE_X109Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y127_SLICE_X109Y127_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y128_SLICE_X108Y128_A5Q),
.Q(CLBLM_L_X72Y127_SLICE_X109Y127_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y127_SLICE_X109Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y127_SLICE_X109Y127_DO5),
.O6(CLBLM_L_X72Y127_SLICE_X109Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff11ff33ff55ffff)
  ) CLBLM_L_X72Y127_SLICE_X109Y127_CLUT (
.I0(CLBLM_L_X72Y126_SLICE_X109Y126_AQ),
.I1(CLBLL_R_X73Y126_SLICE_X110Y126_A5Q),
.I2(1'b1),
.I3(CLBLL_R_X71Y127_SLICE_X107Y127_AQ),
.I4(CLBLL_R_X73Y127_SLICE_X110Y127_BQ),
.I5(CLBLL_R_X75Y127_SLICE_X114Y127_BQ),
.O5(CLBLM_L_X72Y127_SLICE_X109Y127_CO5),
.O6(CLBLM_L_X72Y127_SLICE_X109Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2f222f2200000000)
  ) CLBLM_L_X72Y127_SLICE_X109Y127_BLUT (
.I0(CLBLL_R_X73Y127_SLICE_X110Y127_DQ),
.I1(CLBLL_R_X73Y126_SLICE_X110Y126_A5Q),
.I2(CLBLM_L_X72Y126_SLICE_X109Y126_AQ),
.I3(CLBLL_R_X73Y127_SLICE_X111Y127_AQ),
.I4(1'b1),
.I5(CLBLL_R_X71Y127_SLICE_X107Y127_AQ),
.O5(CLBLM_L_X72Y127_SLICE_X109Y127_BO5),
.O6(CLBLM_L_X72Y127_SLICE_X109Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8f8f3f0ffffffff)
  ) CLBLM_L_X72Y127_SLICE_X109Y127_ALUT (
.I0(CLBLL_R_X73Y127_SLICE_X111Y127_CQ),
.I1(CLBLL_R_X73Y126_SLICE_X110Y126_A5Q),
.I2(CLBLM_L_X72Y127_SLICE_X109Y127_BO6),
.I3(CLBLL_R_X73Y127_SLICE_X110Y127_AQ),
.I4(CLBLM_L_X72Y126_SLICE_X109Y126_AQ),
.I5(CLBLM_L_X72Y127_SLICE_X109Y127_CO6),
.O5(CLBLM_L_X72Y127_SLICE_X109Y127_AO5),
.O6(CLBLM_L_X72Y127_SLICE_X109Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y128_SLICE_X108Y128_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y128_SLICE_X108Y128_BO6),
.Q(CLBLM_L_X72Y128_SLICE_X108Y128_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y128_SLICE_X108Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y128_SLICE_X108Y128_AO6),
.Q(CLBLM_L_X72Y128_SLICE_X108Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y128_SLICE_X108Y128_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y128_SLICE_X108Y128_CO6),
.Q(CLBLM_L_X72Y128_SLICE_X108Y128_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y128_SLICE_X108Y128_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y128_SLICE_X108Y128_DO6),
.Q(CLBLM_L_X72Y128_SLICE_X108Y128_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff003c3ccccccccc)
  ) CLBLM_L_X72Y128_SLICE_X108Y128_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X72Y128_SLICE_X108Y128_CQ),
.I2(CLBLM_L_X74Y128_SLICE_X113Y128_CQ),
.I3(CLBLM_L_X72Y128_SLICE_X108Y128_DQ),
.I4(CLBLM_L_X72Y128_SLICE_X108Y128_BO5),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X72Y128_SLICE_X108Y128_DO5),
.O6(CLBLM_L_X72Y128_SLICE_X108Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7c3c8cccffff0000)
  ) CLBLM_L_X72Y128_SLICE_X108Y128_CLUT (
.I0(CLBLM_L_X72Y127_SLICE_X108Y127_AQ),
.I1(CLBLM_L_X72Y128_SLICE_X108Y128_CQ),
.I2(CLBLM_L_X72Y126_SLICE_X108Y126_CO6),
.I3(CLBLM_L_X72Y128_SLICE_X108Y128_A5Q),
.I4(CLBLM_L_X72Y127_SLICE_X108Y127_CQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X72Y128_SLICE_X108Y128_CO5),
.O6(CLBLM_L_X72Y128_SLICE_X108Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ccf0f3f3ffff)
  ) CLBLM_L_X72Y128_SLICE_X108Y128_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X72Y128_SLICE_X108Y128_A5Q),
.I2(CLBLM_L_X72Y127_SLICE_X108Y127_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X72Y126_SLICE_X108Y126_CO6),
.I5(1'b1),
.O5(CLBLM_L_X72Y128_SLICE_X108Y128_BO5),
.O6(CLBLM_L_X72Y128_SLICE_X108Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf033f0f0aaaaaaaa)
  ) CLBLM_L_X72Y128_SLICE_X108Y128_ALUT (
.I0(CLBLM_L_X74Y128_SLICE_X112Y128_CQ),
.I1(CLBLM_L_X74Y127_SLICE_X112Y127_AO6),
.I2(CLBLM_L_X72Y128_SLICE_X108Y128_AQ),
.I3(CLBLM_L_X72Y127_SLICE_X108Y127_BO6),
.I4(CLBLM_L_X72Y126_SLICE_X108Y126_CO6),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X72Y128_SLICE_X108Y128_AO5),
.O6(CLBLM_L_X72Y128_SLICE_X108Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y128_SLICE_X109Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y128_SLICE_X109Y128_AO5),
.Q(CLBLM_L_X72Y128_SLICE_X109Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y128_SLICE_X109Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y128_SLICE_X109Y128_DO5),
.O6(CLBLM_L_X72Y128_SLICE_X109Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y128_SLICE_X109Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y128_SLICE_X109Y128_CO5),
.O6(CLBLM_L_X72Y128_SLICE_X109Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y128_SLICE_X109Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y128_SLICE_X109Y128_BO5),
.O6(CLBLM_L_X72Y128_SLICE_X109Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaafffff5ffcccc)
  ) CLBLM_L_X72Y128_SLICE_X109Y128_ALUT (
.I0(CLBLM_L_X74Y134_SLICE_X112Y134_DQ),
.I1(CLBLM_L_X72Y123_SLICE_X108Y123_BQ),
.I2(CLBLM_L_X72Y128_SLICE_X109Y128_AQ),
.I3(CLBLL_R_X77Y128_SLICE_X119Y128_AQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLM_L_X72Y128_SLICE_X109Y128_AO5),
.O6(CLBLM_L_X72Y128_SLICE_X109Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y129_SLICE_X108Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y129_SLICE_X108Y129_AO6),
.Q(CLBLM_L_X72Y129_SLICE_X108Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y129_SLICE_X108Y129_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y129_SLICE_X108Y129_BO6),
.Q(CLBLM_L_X72Y129_SLICE_X108Y129_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y129_SLICE_X108Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y129_SLICE_X108Y129_DO5),
.O6(CLBLM_L_X72Y129_SLICE_X108Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y129_SLICE_X108Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y129_SLICE_X108Y129_CO5),
.O6(CLBLM_L_X72Y129_SLICE_X108Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafcfcfa0a0c0c0)
  ) CLBLM_L_X72Y129_SLICE_X108Y129_BLUT (
.I0(CLBLL_R_X71Y130_SLICE_X107Y130_AO6),
.I1(CLBLM_L_X72Y129_SLICE_X108Y129_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(1'b1),
.I4(CLBLL_R_X71Y125_SLICE_X107Y125_BO6),
.I5(CLBLL_R_X71Y129_SLICE_X106Y129_AQ),
.O5(CLBLM_L_X72Y129_SLICE_X108Y129_BO5),
.O6(CLBLM_L_X72Y129_SLICE_X108Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfd0808ffff3f3f)
  ) CLBLM_L_X72Y129_SLICE_X108Y129_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X72Y129_SLICE_X108Y129_AQ),
.I2(CLBLL_R_X71Y125_SLICE_X107Y125_BO6),
.I3(1'b1),
.I4(CLBLL_R_X71Y130_SLICE_X106Y130_BQ),
.I5(1'b1),
.O5(CLBLM_L_X72Y129_SLICE_X108Y129_AO5),
.O6(CLBLM_L_X72Y129_SLICE_X108Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y129_SLICE_X109Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y129_SLICE_X109Y129_DO5),
.O6(CLBLM_L_X72Y129_SLICE_X109Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y129_SLICE_X109Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y129_SLICE_X109Y129_CO5),
.O6(CLBLM_L_X72Y129_SLICE_X109Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y129_SLICE_X109Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y129_SLICE_X109Y129_BO5),
.O6(CLBLM_L_X72Y129_SLICE_X109Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y129_SLICE_X109Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y129_SLICE_X109Y129_AO5),
.O6(CLBLM_L_X72Y129_SLICE_X109Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y130_SLICE_X108Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y130_SLICE_X108Y130_AO5),
.Q(CLBLM_L_X72Y130_SLICE_X108Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y130_SLICE_X108Y130_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y130_SLICE_X108Y130_BO6),
.Q(CLBLM_L_X72Y130_SLICE_X108Y130_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y130_SLICE_X108Y130_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y130_SLICE_X108Y130_CO6),
.Q(CLBLM_L_X72Y130_SLICE_X108Y130_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y130_SLICE_X108Y130_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y130_SLICE_X108Y130_DO6),
.Q(CLBLM_L_X72Y130_SLICE_X108Y130_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5af0ccccf0f0cccc)
  ) CLBLM_L_X72Y130_SLICE_X108Y130_DLUT (
.I0(CLBLL_R_X71Y130_SLICE_X106Y130_BQ),
.I1(CLBLM_L_X72Y130_SLICE_X108Y130_CQ),
.I2(CLBLM_L_X72Y130_SLICE_X108Y130_DQ),
.I3(CLBLL_R_X71Y125_SLICE_X107Y125_BO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X71Y129_SLICE_X106Y129_AQ),
.O5(CLBLM_L_X72Y130_SLICE_X108Y130_DO5),
.O6(CLBLM_L_X72Y130_SLICE_X108Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd5f88a0dd5f88a0)
  ) CLBLM_L_X72Y130_SLICE_X108Y130_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X72Y130_SLICE_X108Y130_CQ),
.I2(CLBLM_L_X72Y131_SLICE_X109Y131_DQ),
.I3(CLBLM_L_X72Y129_SLICE_X108Y129_AO5),
.I4(CLBLM_L_X72Y130_SLICE_X108Y130_BQ),
.I5(1'b1),
.O5(CLBLM_L_X72Y130_SLICE_X108Y130_CO5),
.O6(CLBLM_L_X72Y130_SLICE_X108Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3bc4ff00ccccff00)
  ) CLBLM_L_X72Y130_SLICE_X108Y130_BLUT (
.I0(CLBLM_L_X72Y129_SLICE_X108Y129_AQ),
.I1(CLBLM_L_X72Y130_SLICE_X108Y130_BQ),
.I2(CLBLL_R_X71Y130_SLICE_X106Y130_BQ),
.I3(CLBLM_L_X72Y129_SLICE_X108Y129_BQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X71Y125_SLICE_X107Y125_BO6),
.O5(CLBLM_L_X72Y130_SLICE_X108Y130_BO5),
.O6(CLBLM_L_X72Y130_SLICE_X108Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000f0f0e4eee444)
  ) CLBLM_L_X72Y130_SLICE_X108Y130_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X71Y130_SLICE_X107Y130_AQ),
.I2(CLBLM_L_X72Y130_SLICE_X108Y130_AQ),
.I3(CLBLM_L_X72Y133_SLICE_X109Y133_DO6),
.I4(CLBLM_L_X72Y131_SLICE_X108Y131_AQ),
.I5(1'b1),
.O5(CLBLM_L_X72Y130_SLICE_X108Y130_AO5),
.O6(CLBLM_L_X72Y130_SLICE_X108Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y130_SLICE_X109Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y130_SLICE_X109Y130_AO6),
.Q(CLBLM_L_X72Y130_SLICE_X109Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y130_SLICE_X109Y130_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y130_SLICE_X109Y130_BO6),
.Q(CLBLM_L_X72Y130_SLICE_X109Y130_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y130_SLICE_X109Y130_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y130_SLICE_X109Y130_CO6),
.Q(CLBLM_L_X72Y130_SLICE_X109Y130_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y130_SLICE_X109Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y130_SLICE_X109Y130_DO5),
.O6(CLBLM_L_X72Y130_SLICE_X109Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefeff000101ff00)
  ) CLBLM_L_X72Y130_SLICE_X109Y130_CLUT (
.I0(CLBLM_L_X72Y131_SLICE_X108Y131_AQ),
.I1(CLBLM_L_X72Y133_SLICE_X109Y133_DO6),
.I2(CLBLM_L_X72Y131_SLICE_X108Y131_A5Q),
.I3(CLBLM_L_X72Y130_SLICE_X109Y130_BQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X72Y130_SLICE_X109Y130_CQ),
.O5(CLBLM_L_X72Y130_SLICE_X109Y130_CO5),
.O6(CLBLM_L_X72Y130_SLICE_X109Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5f0a5f0ccf0ccf0)
  ) CLBLM_L_X72Y130_SLICE_X109Y130_BLUT (
.I0(CLBLM_L_X72Y130_SLICE_X108Y130_DQ),
.I1(CLBLM_L_X72Y130_SLICE_X109Y130_BQ),
.I2(CLBLM_L_X72Y130_SLICE_X109Y130_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(1'b1),
.I5(CLBLM_L_X72Y131_SLICE_X109Y131_AO5),
.O5(CLBLM_L_X72Y130_SLICE_X109Y130_BO5),
.O6(CLBLM_L_X72Y130_SLICE_X109Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0e2aaaaaaaa)
  ) CLBLM_L_X72Y130_SLICE_X109Y130_ALUT (
.I0(CLBLM_L_X72Y130_SLICE_X108Y130_DQ),
.I1(CLBLM_L_X72Y133_SLICE_X109Y133_DO6),
.I2(CLBLM_L_X72Y130_SLICE_X109Y130_AQ),
.I3(CLBLM_L_X72Y131_SLICE_X108Y131_A5Q),
.I4(CLBLM_L_X72Y131_SLICE_X108Y131_AQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X72Y130_SLICE_X109Y130_AO5),
.O6(CLBLM_L_X72Y130_SLICE_X109Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y131_SLICE_X108Y131_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y131_SLICE_X108Y131_AO5),
.Q(CLBLM_L_X72Y131_SLICE_X108Y131_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y131_SLICE_X108Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y131_SLICE_X108Y131_AO6),
.Q(CLBLM_L_X72Y131_SLICE_X108Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y131_SLICE_X108Y131_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y131_SLICE_X108Y131_BO6),
.Q(CLBLM_L_X72Y131_SLICE_X108Y131_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y131_SLICE_X108Y131_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y131_SLICE_X108Y131_CO6),
.Q(CLBLM_L_X72Y131_SLICE_X108Y131_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff00aaffaaff)
  ) CLBLM_L_X72Y131_SLICE_X108Y131_DLUT (
.I0(CLBLM_L_X72Y130_SLICE_X108Y130_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X72Y131_SLICE_X108Y131_A5Q),
.I4(CLBLM_L_X72Y133_SLICE_X109Y133_DO6),
.I5(1'b1),
.O5(CLBLM_L_X72Y131_SLICE_X108Y131_DO5),
.O6(CLBLM_L_X72Y131_SLICE_X108Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccee44f0f0f0f0)
  ) CLBLM_L_X72Y131_SLICE_X108Y131_CLUT (
.I0(CLBLM_L_X72Y130_SLICE_X108Y130_AQ),
.I1(CLBLM_L_X72Y131_SLICE_X108Y131_CQ),
.I2(CLBLM_L_X72Y131_SLICE_X108Y131_BQ),
.I3(CLBLM_L_X72Y134_SLICE_X109Y134_AO5),
.I4(CLBLM_L_X72Y131_SLICE_X108Y131_DO6),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X72Y131_SLICE_X108Y131_CO5),
.O6(CLBLM_L_X72Y131_SLICE_X108Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefeff000202ff00)
  ) CLBLM_L_X72Y131_SLICE_X108Y131_BLUT (
.I0(CLBLM_L_X72Y134_SLICE_X109Y134_AO5),
.I1(CLBLM_L_X72Y130_SLICE_X108Y130_AQ),
.I2(CLBLM_L_X72Y131_SLICE_X109Y131_AO6),
.I3(CLBLM_L_X72Y131_SLICE_X109Y131_BQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X72Y131_SLICE_X108Y131_BQ),
.O5(CLBLM_L_X72Y131_SLICE_X108Y131_BO5),
.O6(CLBLM_L_X72Y131_SLICE_X108Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8080a0a2ff887700)
  ) CLBLM_L_X72Y131_SLICE_X108Y131_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X72Y133_SLICE_X109Y133_DO6),
.I2(CLBLM_L_X72Y131_SLICE_X108Y131_AQ),
.I3(CLBLM_L_X72Y130_SLICE_X108Y130_AQ),
.I4(CLBLM_L_X72Y131_SLICE_X108Y131_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X72Y131_SLICE_X108Y131_AO5),
.O6(CLBLM_L_X72Y131_SLICE_X108Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y131_SLICE_X109Y131_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y131_SLICE_X109Y131_BO6),
.Q(CLBLM_L_X72Y131_SLICE_X109Y131_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y131_SLICE_X109Y131_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y131_SLICE_X109Y131_CO6),
.Q(CLBLM_L_X72Y131_SLICE_X109Y131_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y131_SLICE_X109Y131_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y131_SLICE_X109Y131_DO6),
.Q(CLBLM_L_X72Y131_SLICE_X109Y131_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0ccf0cce4cc)
  ) CLBLM_L_X72Y131_SLICE_X109Y131_DLUT (
.I0(CLBLM_L_X72Y131_SLICE_X108Y131_AQ),
.I1(CLBLM_L_X72Y131_SLICE_X109Y131_CQ),
.I2(CLBLM_L_X72Y131_SLICE_X109Y131_DQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X72Y131_SLICE_X108Y131_A5Q),
.I5(CLBLM_L_X72Y133_SLICE_X109Y133_DO6),
.O5(CLBLM_L_X72Y131_SLICE_X109Y131_DO5),
.O6(CLBLM_L_X72Y131_SLICE_X109Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc003cff7800)
  ) CLBLM_L_X72Y131_SLICE_X109Y131_CLUT (
.I0(CLBLM_L_X72Y131_SLICE_X108Y131_AQ),
.I1(CLBLM_L_X72Y131_SLICE_X109Y131_CQ),
.I2(CLBLM_L_X72Y134_SLICE_X109Y134_BO5),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X72Y131_SLICE_X108Y131_A5Q),
.I5(CLBLM_L_X72Y133_SLICE_X109Y133_DO6),
.O5(CLBLM_L_X72Y131_SLICE_X109Y131_CO5),
.O6(CLBLM_L_X72Y131_SLICE_X109Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00ccffcc00)
  ) CLBLM_L_X72Y131_SLICE_X109Y131_BLUT (
.I0(CLBLM_L_X72Y134_SLICE_X109Y134_AO5),
.I1(CLBLM_L_X72Y131_SLICE_X109Y131_BQ),
.I2(1'b1),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X72Y131_SLICE_X109Y131_DQ),
.I5(CLBLM_L_X72Y131_SLICE_X109Y131_AO5),
.O5(CLBLM_L_X72Y131_SLICE_X109Y131_BO5),
.O6(CLBLM_L_X72Y131_SLICE_X109Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ffff00000055)
  ) CLBLM_L_X72Y131_SLICE_X109Y131_ALUT (
.I0(CLBLM_L_X72Y131_SLICE_X108Y131_A5Q),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X72Y133_SLICE_X109Y133_DO6),
.I4(CLBLM_L_X72Y131_SLICE_X108Y131_AQ),
.I5(1'b1),
.O5(CLBLM_L_X72Y131_SLICE_X109Y131_AO5),
.O6(CLBLM_L_X72Y131_SLICE_X109Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y132_SLICE_X108Y132_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y132_SLICE_X108Y132_AO6),
.Q(CLBLM_L_X72Y132_SLICE_X108Y132_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y132_SLICE_X108Y132_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y132_SLICE_X108Y132_BO6),
.Q(CLBLM_L_X72Y132_SLICE_X108Y132_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y132_SLICE_X108Y132_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y132_SLICE_X108Y132_CO6),
.Q(CLBLM_L_X72Y132_SLICE_X108Y132_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y132_SLICE_X108Y132_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y132_SLICE_X108Y132_DO6),
.Q(CLBLM_L_X72Y132_SLICE_X108Y132_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f7d5a0a0a280)
  ) CLBLM_L_X72Y132_SLICE_X108Y132_DLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X72Y133_SLICE_X108Y133_DO5),
.I2(CLBLM_L_X72Y132_SLICE_X108Y132_DQ),
.I3(CLBLL_R_X73Y132_SLICE_X110Y132_AO6),
.I4(CLBLL_R_X73Y132_SLICE_X110Y132_BO6),
.I5(CLBLM_L_X72Y133_SLICE_X108Y133_CQ),
.O5(CLBLM_L_X72Y132_SLICE_X108Y132_DO5),
.O6(CLBLM_L_X72Y132_SLICE_X108Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfad8fafa72505050)
  ) CLBLM_L_X72Y132_SLICE_X108Y132_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X73Y132_SLICE_X110Y132_BO6),
.I2(CLBLM_L_X72Y132_SLICE_X108Y132_DQ),
.I3(CLBLL_R_X73Y132_SLICE_X110Y132_AO6),
.I4(CLBLL_R_X71Y132_SLICE_X107Y132_AO6),
.I5(CLBLM_L_X72Y132_SLICE_X108Y132_CQ),
.O5(CLBLM_L_X72Y132_SLICE_X108Y132_CO5),
.O6(CLBLM_L_X72Y132_SLICE_X108Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaf0f0ccccf0f0)
  ) CLBLM_L_X72Y132_SLICE_X108Y132_BLUT (
.I0(CLBLL_R_X73Y132_SLICE_X110Y132_AO6),
.I1(CLBLM_L_X72Y132_SLICE_X108Y132_BQ),
.I2(CLBLM_L_X72Y132_SLICE_X108Y132_CQ),
.I3(CLBLM_L_X72Y133_SLICE_X108Y133_BO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X72Y133_SLICE_X108Y133_A5Q),
.O5(CLBLM_L_X72Y132_SLICE_X108Y132_BO5),
.O6(CLBLM_L_X72Y132_SLICE_X108Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f5ccccf0a0cccc)
  ) CLBLM_L_X72Y132_SLICE_X108Y132_ALUT (
.I0(CLBLL_R_X71Y132_SLICE_X107Y132_AQ),
.I1(CLBLM_L_X72Y134_SLICE_X108Y134_AQ),
.I2(CLBLM_L_X72Y132_SLICE_X108Y132_AQ),
.I3(CLBLM_L_X72Y133_SLICE_X108Y133_BO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X73Y132_SLICE_X110Y132_AO6),
.O5(CLBLM_L_X72Y132_SLICE_X108Y132_AO5),
.O6(CLBLM_L_X72Y132_SLICE_X108Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y132_SLICE_X109Y132_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y133_SLICE_X108Y133_AQ),
.Q(CLBLM_L_X72Y132_SLICE_X109Y132_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33bb00aa00000000)
  ) CLBLM_L_X72Y132_SLICE_X109Y132_DLUT (
.I0(CLBLM_L_X72Y132_SLICE_X108Y132_AQ),
.I1(CLBLL_R_X71Y131_SLICE_X107Y131_A5Q),
.I2(1'b1),
.I3(CLBLL_R_X71Y131_SLICE_X106Y131_AQ),
.I4(CLBLM_L_X72Y132_SLICE_X108Y132_DQ),
.I5(CLBLL_R_X71Y132_SLICE_X106Y132_AQ),
.O5(CLBLM_L_X72Y132_SLICE_X109Y132_DO5),
.O6(CLBLM_L_X72Y132_SLICE_X109Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000eeaacc00)
  ) CLBLM_L_X72Y132_SLICE_X109Y132_CLUT (
.I0(CLBLM_L_X72Y132_SLICE_X108Y132_CQ),
.I1(CLBLM_L_X72Y133_SLICE_X108Y133_CQ),
.I2(1'b1),
.I3(CLBLL_R_X71Y131_SLICE_X107Y131_A5Q),
.I4(CLBLL_R_X71Y131_SLICE_X106Y131_AQ),
.I5(CLBLL_R_X71Y132_SLICE_X106Y132_AQ),
.O5(CLBLM_L_X72Y132_SLICE_X109Y132_CO5),
.O6(CLBLM_L_X72Y132_SLICE_X109Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefeeeeeefeeefee)
  ) CLBLM_L_X72Y132_SLICE_X109Y132_BLUT (
.I0(CLBLM_L_X72Y132_SLICE_X109Y132_DO6),
.I1(CLBLM_L_X72Y132_SLICE_X109Y132_CO6),
.I2(CLBLL_R_X71Y131_SLICE_X106Y131_AQ),
.I3(CLBLM_L_X72Y132_SLICE_X108Y132_BQ),
.I4(CLBLM_L_X72Y134_SLICE_X108Y134_AQ),
.I5(CLBLL_R_X71Y131_SLICE_X107Y131_A5Q),
.O5(CLBLM_L_X72Y132_SLICE_X109Y132_BO5),
.O6(CLBLM_L_X72Y132_SLICE_X109Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7333333300000000)
  ) CLBLM_L_X72Y132_SLICE_X109Y132_ALUT (
.I0(CLBLM_L_X74Y134_SLICE_X113Y134_CQ),
.I1(CLBLM_L_X60Y92_SLICE_X90Y92_AQ),
.I2(CLBLL_R_X73Y133_SLICE_X110Y133_A5Q),
.I3(CLBLM_L_X74Y134_SLICE_X113Y134_A5Q),
.I4(CLBLM_L_X70Y136_SLICE_X105Y136_CO6),
.I5(CLBLL_R_X73Y132_SLICE_X111Y132_BO6),
.O5(CLBLM_L_X72Y132_SLICE_X109Y132_AO5),
.O6(CLBLM_L_X72Y132_SLICE_X109Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y133_SLICE_X108Y133_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y133_SLICE_X108Y133_AO5),
.Q(CLBLM_L_X72Y133_SLICE_X108Y133_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y133_SLICE_X108Y133_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y133_SLICE_X108Y133_AO6),
.Q(CLBLM_L_X72Y133_SLICE_X108Y133_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y133_SLICE_X108Y133_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y133_SLICE_X108Y133_CO6),
.Q(CLBLM_L_X72Y133_SLICE_X108Y133_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0fff0aaffaaff)
  ) CLBLM_L_X72Y133_SLICE_X108Y133_DLUT (
.I0(CLBLL_R_X71Y132_SLICE_X107Y132_AQ),
.I1(1'b1),
.I2(CLBLL_R_X73Y132_SLICE_X110Y132_BO6),
.I3(CLBLM_L_X72Y133_SLICE_X108Y133_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y133_SLICE_X108Y133_DO5),
.O6(CLBLM_L_X72Y133_SLICE_X108Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0afcfa0c0)
  ) CLBLM_L_X72Y133_SLICE_X108Y133_CLUT (
.I0(CLBLL_R_X73Y132_SLICE_X110Y132_AO6),
.I1(CLBLM_L_X72Y133_SLICE_X108Y133_CQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLL_R_X71Y132_SLICE_X107Y132_AQ),
.I4(CLBLM_L_X72Y132_SLICE_X108Y132_AQ),
.I5(CLBLM_L_X72Y133_SLICE_X108Y133_DO6),
.O5(CLBLM_L_X72Y133_SLICE_X108Y133_CO5),
.O6(CLBLM_L_X72Y133_SLICE_X108Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfcfcf01010101)
  ) CLBLM_L_X72Y133_SLICE_X108Y133_BLUT (
.I0(CLBLM_L_X72Y133_SLICE_X108Y133_A5Q),
.I1(CLBLL_R_X73Y132_SLICE_X110Y132_BO6),
.I2(CLBLM_L_X72Y133_SLICE_X108Y133_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y133_SLICE_X108Y133_BO5),
.O6(CLBLM_L_X72Y133_SLICE_X108Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc040c044bbff8800)
  ) CLBLM_L_X72Y133_SLICE_X108Y133_ALUT (
.I0(CLBLM_L_X72Y133_SLICE_X108Y133_A5Q),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_L_X72Y133_SLICE_X108Y133_AQ),
.I3(CLBLL_R_X73Y132_SLICE_X110Y132_BO6),
.I4(CLBLL_R_X71Y132_SLICE_X107Y132_AQ),
.I5(1'b1),
.O5(CLBLM_L_X72Y133_SLICE_X108Y133_AO5),
.O6(CLBLM_L_X72Y133_SLICE_X108Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y133_SLICE_X109Y133_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y133_SLICE_X109Y133_BO6),
.Q(CLBLM_L_X72Y133_SLICE_X109Y133_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd500550055005500)
  ) CLBLM_L_X72Y133_SLICE_X109Y133_DLUT (
.I0(CLBLM_L_X60Y94_SLICE_X90Y94_AQ),
.I1(CLBLM_L_X70Y136_SLICE_X105Y136_CO6),
.I2(CLBLM_L_X74Y134_SLICE_X113Y134_CQ),
.I3(CLBLL_R_X73Y133_SLICE_X111Y133_CO6),
.I4(CLBLL_R_X73Y133_SLICE_X110Y133_A5Q),
.I5(CLBLM_L_X74Y134_SLICE_X113Y134_A5Q),
.O5(CLBLM_L_X72Y133_SLICE_X109Y133_DO5),
.O6(CLBLM_L_X72Y133_SLICE_X109Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55005500d5005500)
  ) CLBLM_L_X72Y133_SLICE_X109Y133_CLUT (
.I0(CLBLL_R_X71Y134_SLICE_X106Y134_AQ),
.I1(CLBLM_L_X70Y136_SLICE_X105Y136_CO6),
.I2(CLBLM_L_X74Y134_SLICE_X113Y134_CQ),
.I3(CLBLL_R_X73Y133_SLICE_X111Y133_BO6),
.I4(CLBLL_R_X73Y133_SLICE_X110Y133_A5Q),
.I5(CLBLM_L_X74Y134_SLICE_X113Y134_A5Q),
.O5(CLBLM_L_X72Y133_SLICE_X109Y133_CO5),
.O6(CLBLM_L_X72Y133_SLICE_X109Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfcfdfc0c0c080)
  ) CLBLM_L_X72Y133_SLICE_X109Y133_BLUT (
.I0(CLBLM_L_X72Y133_SLICE_X108Y133_A5Q),
.I1(CLBLM_L_X72Y133_SLICE_X109Y133_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLL_R_X73Y132_SLICE_X110Y132_BO6),
.I4(CLBLM_L_X72Y133_SLICE_X108Y133_AQ),
.I5(CLBLL_R_X73Y133_SLICE_X110Y133_BQ),
.O5(CLBLM_L_X72Y133_SLICE_X109Y133_BO5),
.O6(CLBLM_L_X72Y133_SLICE_X109Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcfffcfffccffff)
  ) CLBLM_L_X72Y133_SLICE_X109Y133_ALUT (
.I0(1'b1),
.I1(CLBLL_R_X73Y132_SLICE_X111Y132_AO5),
.I2(CLBLL_R_X73Y131_SLICE_X110Y131_AQ),
.I3(CLBLM_L_X74Y133_SLICE_X112Y133_AQ),
.I4(CLBLM_L_X74Y132_SLICE_X112Y132_CQ),
.I5(1'b1),
.O5(CLBLM_L_X72Y133_SLICE_X109Y133_AO5),
.O6(CLBLM_L_X72Y133_SLICE_X109Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y134_SLICE_X108Y134_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y134_SLICE_X108Y134_AO6),
.Q(CLBLM_L_X72Y134_SLICE_X108Y134_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y134_SLICE_X108Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y134_SLICE_X108Y134_DO5),
.O6(CLBLM_L_X72Y134_SLICE_X108Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y134_SLICE_X108Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y134_SLICE_X108Y134_CO5),
.O6(CLBLM_L_X72Y134_SLICE_X108Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y134_SLICE_X108Y134_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y134_SLICE_X108Y134_BO5),
.O6(CLBLM_L_X72Y134_SLICE_X108Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ccccf0f0cccc)
  ) CLBLM_L_X72Y134_SLICE_X108Y134_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X72Y133_SLICE_X109Y133_BQ),
.I2(CLBLM_L_X72Y134_SLICE_X108Y134_AQ),
.I3(CLBLL_R_X73Y132_SLICE_X110Y132_AO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X72Y133_SLICE_X108Y133_BO5),
.O5(CLBLM_L_X72Y134_SLICE_X108Y134_AO5),
.O6(CLBLM_L_X72Y134_SLICE_X108Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y134_SLICE_X109Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y134_SLICE_X109Y134_DO5),
.O6(CLBLM_L_X72Y134_SLICE_X109Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y134_SLICE_X109Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y134_SLICE_X109Y134_CO5),
.O6(CLBLM_L_X72Y134_SLICE_X109Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffccffeeffee)
  ) CLBLM_L_X72Y134_SLICE_X109Y134_BLUT (
.I0(CLBLM_L_X74Y133_SLICE_X112Y133_CQ),
.I1(CLBLM_L_X74Y132_SLICE_X112Y132_CQ),
.I2(1'b1),
.I3(CLBLL_R_X73Y132_SLICE_X111Y132_AO5),
.I4(CLBLM_L_X74Y134_SLICE_X113Y134_AQ),
.I5(1'b1),
.O5(CLBLM_L_X72Y134_SLICE_X109Y134_BO5),
.O6(CLBLM_L_X72Y134_SLICE_X109Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffcfcfffffafa)
  ) CLBLM_L_X72Y134_SLICE_X109Y134_ALUT (
.I0(CLBLM_L_X74Y133_SLICE_X112Y133_CQ),
.I1(CLBLM_L_X74Y134_SLICE_X113Y134_AQ),
.I2(CLBLL_R_X73Y131_SLICE_X110Y131_AQ),
.I3(1'b1),
.I4(CLBLL_R_X73Y132_SLICE_X111Y132_AO5),
.I5(1'b1),
.O5(CLBLM_L_X72Y134_SLICE_X109Y134_AO5),
.O6(CLBLM_L_X72Y134_SLICE_X109Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y102_SLICE_X112Y102_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y102_SLICE_X112Y102_AO6),
.Q(CLBLM_L_X74Y102_SLICE_X112Y102_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y102_SLICE_X112Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y102_SLICE_X112Y102_DO5),
.O6(CLBLM_L_X74Y102_SLICE_X112Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y102_SLICE_X112Y102_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y102_SLICE_X112Y102_CO5),
.O6(CLBLM_L_X74Y102_SLICE_X112Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y102_SLICE_X112Y102_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y102_SLICE_X112Y102_BO5),
.O6(CLBLM_L_X74Y102_SLICE_X112Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1e0f1e0ffff0000)
  ) CLBLM_L_X74Y102_SLICE_X112Y102_ALUT (
.I0(CLBLM_L_X72Y103_SLICE_X108Y103_DO5),
.I1(CLBLM_L_X72Y103_SLICE_X108Y103_CO6),
.I2(CLBLM_L_X74Y102_SLICE_X112Y102_AQ),
.I3(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I4(CLBLL_R_X73Y101_SLICE_X110Y101_AQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X74Y102_SLICE_X112Y102_AO5),
.O6(CLBLM_L_X74Y102_SLICE_X112Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y102_SLICE_X113Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y102_SLICE_X113Y102_DO5),
.O6(CLBLM_L_X74Y102_SLICE_X113Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y102_SLICE_X113Y102_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y102_SLICE_X113Y102_CO5),
.O6(CLBLM_L_X74Y102_SLICE_X113Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y102_SLICE_X113Y102_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y102_SLICE_X113Y102_BO5),
.O6(CLBLM_L_X74Y102_SLICE_X113Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y102_SLICE_X113Y102_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y102_SLICE_X113Y102_AO5),
.O6(CLBLM_L_X74Y102_SLICE_X113Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y103_SLICE_X112Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y103_SLICE_X112Y103_AO6),
.Q(CLBLM_L_X74Y103_SLICE_X112Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y103_SLICE_X112Y103_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y103_SLICE_X112Y103_BO6),
.Q(CLBLM_L_X74Y103_SLICE_X112Y103_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf800000088000000)
  ) CLBLM_L_X74Y103_SLICE_X112Y103_DLUT (
.I0(CLBLM_L_X74Y103_SLICE_X113Y103_AQ),
.I1(CLBLM_L_X72Y103_SLICE_X109Y103_AQ),
.I2(CLBLL_R_X75Y103_SLICE_X115Y103_AQ),
.I3(CLBLM_L_X72Y104_SLICE_X109Y104_BQ),
.I4(CLBLM_L_X72Y104_SLICE_X109Y104_B5Q),
.I5(CLBLM_L_X74Y104_SLICE_X112Y104_AQ),
.O5(CLBLM_L_X74Y103_SLICE_X112Y103_DO5),
.O6(CLBLM_L_X74Y103_SLICE_X112Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000aa808080)
  ) CLBLM_L_X74Y103_SLICE_X112Y103_CLUT (
.I0(CLBLM_L_X72Y104_SLICE_X109Y104_BQ),
.I1(CLBLL_R_X73Y103_SLICE_X110Y103_A5Q),
.I2(CLBLM_L_X74Y103_SLICE_X112Y103_AQ),
.I3(CLBLL_R_X73Y102_SLICE_X110Y102_A5Q),
.I4(CLBLM_L_X74Y103_SLICE_X112Y103_BQ),
.I5(CLBLM_L_X72Y104_SLICE_X109Y104_B5Q),
.O5(CLBLM_L_X74Y103_SLICE_X112Y103_CO5),
.O6(CLBLM_L_X74Y103_SLICE_X112Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfd08f80cfc0cfc0)
  ) CLBLM_L_X74Y103_SLICE_X112Y103_BLUT (
.I0(CLBLL_R_X73Y104_SLICE_X110Y104_DO6),
.I1(CLBLM_L_X74Y103_SLICE_X112Y103_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLL_R_X73Y103_SLICE_X111Y103_AQ),
.I4(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I5(CLBLM_L_X72Y103_SLICE_X108Y103_A5Q),
.O5(CLBLM_L_X74Y103_SLICE_X112Y103_BO5),
.O6(CLBLM_L_X74Y103_SLICE_X112Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000e2ffe200)
  ) CLBLM_L_X74Y103_SLICE_X112Y103_ALUT (
.I0(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I1(CLBLM_L_X72Y103_SLICE_X108Y103_BO6),
.I2(CLBLM_L_X74Y103_SLICE_X112Y103_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLL_R_X73Y102_SLICE_X111Y102_AQ),
.I5(CLBLL_R_X73Y104_SLICE_X110Y104_DO6),
.O5(CLBLM_L_X74Y103_SLICE_X112Y103_AO5),
.O6(CLBLM_L_X74Y103_SLICE_X112Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y103_SLICE_X113Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y103_SLICE_X113Y103_AO6),
.Q(CLBLM_L_X74Y103_SLICE_X113Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y103_SLICE_X113Y103_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y103_SLICE_X113Y103_BO6),
.Q(CLBLM_L_X74Y103_SLICE_X113Y103_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc0ff00ff00ff00)
  ) CLBLM_L_X74Y103_SLICE_X113Y103_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X72Y104_SLICE_X109Y104_B5Q),
.I2(CLBLL_R_X73Y103_SLICE_X111Y103_A5Q),
.I3(CLBLM_L_X74Y103_SLICE_X113Y103_CO6),
.I4(CLBLL_R_X73Y101_SLICE_X110Y101_AQ),
.I5(CLBLM_L_X72Y104_SLICE_X109Y104_BQ),
.O5(CLBLM_L_X74Y103_SLICE_X113Y103_DO5),
.O6(CLBLM_L_X74Y103_SLICE_X113Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0ff0f02f0ff2f0)
  ) CLBLM_L_X74Y103_SLICE_X113Y103_CLUT (
.I0(CLBLM_L_X74Y102_SLICE_X112Y102_AQ),
.I1(CLBLM_L_X72Y104_SLICE_X109Y104_B5Q),
.I2(CLBLL_R_X73Y104_SLICE_X110Y104_A5Q),
.I3(CLBLM_L_X62Y95_SLICE_X92Y95_AQ),
.I4(CLBLL_R_X75Y103_SLICE_X115Y103_AQ),
.I5(CLBLM_L_X72Y104_SLICE_X109Y104_BQ),
.O5(CLBLM_L_X74Y103_SLICE_X113Y103_CO5),
.O6(CLBLM_L_X74Y103_SLICE_X113Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccddf0f0cc88f0f0)
  ) CLBLM_L_X74Y103_SLICE_X113Y103_BLUT (
.I0(CLBLL_R_X73Y104_SLICE_X110Y104_DO6),
.I1(CLBLM_L_X74Y103_SLICE_X113Y103_BQ),
.I2(CLBLM_L_X74Y103_SLICE_X113Y103_AQ),
.I3(CLBLM_L_X72Y103_SLICE_X108Y103_DO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.O5(CLBLM_L_X74Y103_SLICE_X113Y103_BO5),
.O6(CLBLM_L_X74Y103_SLICE_X113Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f7c0c4f3b3c080)
  ) CLBLM_L_X74Y103_SLICE_X113Y103_ALUT (
.I0(CLBLM_L_X72Y103_SLICE_X108Y103_BO5),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_L_X74Y103_SLICE_X113Y103_AQ),
.I3(CLBLL_R_X73Y104_SLICE_X110Y104_DO6),
.I4(CLBLM_L_X74Y103_SLICE_X112Y103_AQ),
.I5(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.O5(CLBLM_L_X74Y103_SLICE_X113Y103_AO5),
.O6(CLBLM_L_X74Y103_SLICE_X113Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y104_SLICE_X112Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y104_SLICE_X112Y104_AO6),
.Q(CLBLM_L_X74Y104_SLICE_X112Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y104_SLICE_X112Y104_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y104_SLICE_X112Y104_BO6),
.Q(CLBLM_L_X74Y104_SLICE_X112Y104_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y104_SLICE_X112Y104_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y104_SLICE_X112Y104_CO6),
.Q(CLBLM_L_X74Y104_SLICE_X112Y104_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y104_SLICE_X112Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y104_SLICE_X112Y104_DO5),
.O6(CLBLM_L_X74Y104_SLICE_X112Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccff00cacaff00)
  ) CLBLM_L_X74Y104_SLICE_X112Y104_CLUT (
.I0(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I1(CLBLM_L_X74Y104_SLICE_X112Y104_CQ),
.I2(CLBLL_R_X73Y104_SLICE_X110Y104_DO5),
.I3(CLBLM_L_X74Y104_SLICE_X112Y104_BQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X72Y103_SLICE_X108Y103_DO6),
.O5(CLBLM_L_X74Y104_SLICE_X112Y104_CO5),
.O6(CLBLM_L_X74Y104_SLICE_X112Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafafad8505050d8)
  ) CLBLM_L_X74Y104_SLICE_X112Y104_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I2(CLBLM_L_X74Y104_SLICE_X112Y104_AQ),
.I3(CLBLM_L_X72Y103_SLICE_X108Y103_BO5),
.I4(CLBLL_R_X73Y104_SLICE_X110Y104_DO5),
.I5(CLBLM_L_X74Y104_SLICE_X112Y104_BQ),
.O5(CLBLM_L_X74Y104_SLICE_X112Y104_BO5),
.O6(CLBLM_L_X74Y104_SLICE_X112Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a0f7d5a280)
  ) CLBLM_L_X74Y104_SLICE_X112Y104_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X72Y103_SLICE_X108Y103_BO6),
.I2(CLBLM_L_X74Y104_SLICE_X112Y104_AQ),
.I3(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I4(CLBLM_L_X74Y103_SLICE_X112Y103_BQ),
.I5(CLBLL_R_X73Y104_SLICE_X110Y104_DO5),
.O5(CLBLM_L_X74Y104_SLICE_X112Y104_AO5),
.O6(CLBLM_L_X74Y104_SLICE_X112Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y104_SLICE_X113Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y104_SLICE_X113Y104_DO5),
.O6(CLBLM_L_X74Y104_SLICE_X113Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y104_SLICE_X113Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y104_SLICE_X113Y104_CO5),
.O6(CLBLM_L_X74Y104_SLICE_X113Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y104_SLICE_X113Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y104_SLICE_X113Y104_BO5),
.O6(CLBLM_L_X74Y104_SLICE_X113Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y104_SLICE_X113Y104_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y104_SLICE_X113Y104_AO5),
.O6(CLBLM_L_X74Y104_SLICE_X113Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y107_SLICE_X112Y107_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y107_SLICE_X112Y107_AO6),
.Q(CLBLM_L_X74Y107_SLICE_X112Y107_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y107_SLICE_X112Y107_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y107_SLICE_X112Y107_BO6),
.Q(CLBLM_L_X74Y107_SLICE_X112Y107_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y107_SLICE_X112Y107_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y107_SLICE_X112Y107_CO6),
.Q(CLBLM_L_X74Y107_SLICE_X112Y107_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y107_SLICE_X112Y107_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y107_SLICE_X112Y107_DO6),
.Q(CLBLM_L_X74Y107_SLICE_X112Y107_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0f7a2d580)
  ) CLBLM_L_X74Y107_SLICE_X112Y107_DLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X72Y108_SLICE_X108Y108_BO6),
.I2(CLBLM_L_X74Y107_SLICE_X112Y107_DQ),
.I3(CLBLM_L_X74Y107_SLICE_X112Y107_BQ),
.I4(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I5(CLBLM_L_X72Y108_SLICE_X109Y108_CO6),
.O5(CLBLM_L_X74Y107_SLICE_X112Y107_DO5),
.O6(CLBLM_L_X74Y107_SLICE_X112Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccf0ddf088f0)
  ) CLBLM_L_X74Y107_SLICE_X112Y107_CLUT (
.I0(CLBLM_L_X72Y108_SLICE_X108Y108_BO5),
.I1(CLBLM_L_X74Y107_SLICE_X112Y107_CQ),
.I2(CLBLL_R_X73Y107_SLICE_X111Y107_DQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I5(CLBLM_L_X72Y108_SLICE_X109Y108_BO5),
.O5(CLBLM_L_X74Y107_SLICE_X112Y107_CO5),
.O6(CLBLM_L_X74Y107_SLICE_X112Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcdc8ffffcdc80000)
  ) CLBLM_L_X74Y107_SLICE_X112Y107_BLUT (
.I0(CLBLM_L_X72Y108_SLICE_X108Y108_BO6),
.I1(CLBLM_L_X74Y107_SLICE_X112Y107_BQ),
.I2(CLBLM_L_X72Y108_SLICE_X109Y108_BO5),
.I3(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X73Y107_SLICE_X110Y107_AQ),
.O5(CLBLM_L_X74Y107_SLICE_X112Y107_BO5),
.O6(CLBLM_L_X74Y107_SLICE_X112Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff00e4e4ff00)
  ) CLBLM_L_X74Y107_SLICE_X112Y107_ALUT (
.I0(CLBLM_L_X72Y109_SLICE_X108Y109_BO6),
.I1(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I2(CLBLM_L_X74Y107_SLICE_X112Y107_AQ),
.I3(CLBLL_R_X73Y107_SLICE_X111Y107_CQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X72Y108_SLICE_X109Y108_CO5),
.O5(CLBLM_L_X74Y107_SLICE_X112Y107_AO5),
.O6(CLBLM_L_X74Y107_SLICE_X112Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y107_SLICE_X113Y107_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y107_SLICE_X113Y107_AO6),
.Q(CLBLM_L_X74Y107_SLICE_X113Y107_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y107_SLICE_X113Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y107_SLICE_X113Y107_DO5),
.O6(CLBLM_L_X74Y107_SLICE_X113Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y107_SLICE_X113Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y107_SLICE_X113Y107_CO5),
.O6(CLBLM_L_X74Y107_SLICE_X113Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y107_SLICE_X113Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y107_SLICE_X113Y107_BO5),
.O6(CLBLM_L_X74Y107_SLICE_X113Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f5dda0a0a088)
  ) CLBLM_L_X74Y107_SLICE_X113Y107_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I2(CLBLM_L_X74Y107_SLICE_X113Y107_AQ),
.I3(CLBLM_L_X72Y108_SLICE_X109Y108_CO6),
.I4(CLBLM_L_X72Y108_SLICE_X108Y108_BO5),
.I5(CLBLM_L_X74Y107_SLICE_X112Y107_CQ),
.O5(CLBLM_L_X74Y107_SLICE_X113Y107_AO5),
.O6(CLBLM_L_X74Y107_SLICE_X113Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y109_SLICE_X112Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y109_SLICE_X112Y109_DO5),
.O6(CLBLM_L_X74Y109_SLICE_X112Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y109_SLICE_X112Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y109_SLICE_X112Y109_CO5),
.O6(CLBLM_L_X74Y109_SLICE_X112Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y109_SLICE_X112Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y109_SLICE_X112Y109_BO5),
.O6(CLBLM_L_X74Y109_SLICE_X112Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y109_SLICE_X112Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y109_SLICE_X112Y109_AO5),
.O6(CLBLM_L_X74Y109_SLICE_X112Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y109_SLICE_X113Y109_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y109_SLICE_X113Y109_AO5),
.Q(CLBLM_L_X74Y109_SLICE_X113Y109_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y109_SLICE_X113Y109_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y109_SLICE_X113Y109_AO6),
.Q(CLBLM_L_X74Y109_SLICE_X113Y109_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y109_SLICE_X113Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y109_SLICE_X113Y109_DO5),
.O6(CLBLM_L_X74Y109_SLICE_X113Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y109_SLICE_X113Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y109_SLICE_X113Y109_CO5),
.O6(CLBLM_L_X74Y109_SLICE_X113Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y109_SLICE_X113Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y109_SLICE_X113Y109_BO5),
.O6(CLBLM_L_X74Y109_SLICE_X113Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000f0066cc66cc)
  ) CLBLM_L_X74Y109_SLICE_X113Y109_ALUT (
.I0(CLBLM_L_X72Y109_SLICE_X109Y109_DQ),
.I1(CLBLL_R_X73Y109_SLICE_X110Y109_AQ),
.I2(CLBLM_L_X74Y109_SLICE_X113Y109_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLL_R_X75Y113_SLICE_X114Y113_AQ),
.I5(1'b1),
.O5(CLBLM_L_X74Y109_SLICE_X113Y109_AO5),
.O6(CLBLM_L_X74Y109_SLICE_X113Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y117_SLICE_X112Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y116_SLICE_X108Y116_AQ),
.Q(CLBLM_L_X74Y117_SLICE_X112Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y117_SLICE_X112Y117_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y117_SLICE_X112Y117_AQ),
.Q(CLBLM_L_X74Y117_SLICE_X112Y117_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y117_SLICE_X112Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y117_SLICE_X112Y117_DO5),
.O6(CLBLM_L_X74Y117_SLICE_X112Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y117_SLICE_X112Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y117_SLICE_X112Y117_CO5),
.O6(CLBLM_L_X74Y117_SLICE_X112Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y117_SLICE_X112Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y117_SLICE_X112Y117_BO5),
.O6(CLBLM_L_X74Y117_SLICE_X112Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y117_SLICE_X112Y117_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y117_SLICE_X112Y117_AO5),
.O6(CLBLM_L_X74Y117_SLICE_X112Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y117_SLICE_X113Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y117_SLICE_X113Y117_DO5),
.O6(CLBLM_L_X74Y117_SLICE_X113Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y117_SLICE_X113Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y117_SLICE_X113Y117_CO5),
.O6(CLBLM_L_X74Y117_SLICE_X113Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y117_SLICE_X113Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y117_SLICE_X113Y117_BO5),
.O6(CLBLM_L_X74Y117_SLICE_X113Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y117_SLICE_X113Y117_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y117_SLICE_X113Y117_AO5),
.O6(CLBLM_L_X74Y117_SLICE_X113Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y118_SLICE_X112Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y118_SLICE_X112Y118_AO6),
.Q(CLBLM_L_X74Y118_SLICE_X112Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y118_SLICE_X112Y118_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y118_SLICE_X112Y118_CO6),
.Q(CLBLM_L_X74Y118_SLICE_X112Y118_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y118_SLICE_X112Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y118_SLICE_X112Y118_DO5),
.O6(CLBLM_L_X74Y118_SLICE_X112Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8fad8d8d850d8)
  ) CLBLM_L_X74Y118_SLICE_X112Y118_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X74Y118_SLICE_X112Y118_CQ),
.I2(CLBLM_L_X74Y118_SLICE_X112Y118_AQ),
.I3(CLBLM_L_X74Y119_SLICE_X113Y119_AO6),
.I4(CLBLM_L_X74Y118_SLICE_X112Y118_BO5),
.I5(CLBLL_R_X75Y124_SLICE_X115Y124_BQ),
.O5(CLBLM_L_X74Y118_SLICE_X112Y118_CO5),
.O6(CLBLM_L_X74Y118_SLICE_X112Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff0ff0fff0fff)
  ) CLBLM_L_X74Y118_SLICE_X112Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X72Y118_SLICE_X108Y118_CQ),
.I3(CLBLM_R_X65Y105_SLICE_X99Y105_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y118_SLICE_X112Y118_BO5),
.O6(CLBLM_L_X74Y118_SLICE_X112Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccaaaaf0f0aaaa)
  ) CLBLM_L_X74Y118_SLICE_X112Y118_ALUT (
.I0(CLBLM_L_X74Y119_SLICE_X112Y119_DQ),
.I1(CLBLL_R_X75Y124_SLICE_X115Y124_BQ),
.I2(CLBLM_L_X74Y118_SLICE_X112Y118_AQ),
.I3(CLBLM_L_X74Y118_SLICE_X112Y118_BO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X74Y119_SLICE_X113Y119_AO6),
.O5(CLBLM_L_X74Y118_SLICE_X112Y118_AO5),
.O6(CLBLM_L_X74Y118_SLICE_X112Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y118_SLICE_X113Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y118_SLICE_X113Y118_DO5),
.O6(CLBLM_L_X74Y118_SLICE_X113Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y118_SLICE_X113Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y118_SLICE_X113Y118_CO5),
.O6(CLBLM_L_X74Y118_SLICE_X113Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y118_SLICE_X113Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y118_SLICE_X113Y118_BO5),
.O6(CLBLM_L_X74Y118_SLICE_X113Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y118_SLICE_X113Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y118_SLICE_X113Y118_AO5),
.O6(CLBLM_L_X74Y118_SLICE_X113Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y119_SLICE_X112Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y119_SLICE_X112Y119_AO6),
.Q(CLBLM_L_X74Y119_SLICE_X112Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y119_SLICE_X112Y119_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y119_SLICE_X112Y119_CO6),
.Q(CLBLM_L_X74Y119_SLICE_X112Y119_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y119_SLICE_X112Y119_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y119_SLICE_X112Y119_DO6),
.Q(CLBLM_L_X74Y119_SLICE_X112Y119_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccfaccf0cc50cc)
  ) CLBLM_L_X74Y119_SLICE_X112Y119_DLUT (
.I0(CLBLM_L_X74Y119_SLICE_X113Y119_AO6),
.I1(CLBLM_L_X74Y119_SLICE_X112Y119_CQ),
.I2(CLBLM_L_X74Y119_SLICE_X112Y119_DQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X74Y119_SLICE_X112Y119_BO5),
.I5(CLBLL_R_X75Y124_SLICE_X115Y124_BQ),
.O5(CLBLM_L_X74Y119_SLICE_X112Y119_DO5),
.O6(CLBLM_L_X74Y119_SLICE_X112Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffceffcc00c400)
  ) CLBLM_L_X74Y119_SLICE_X112Y119_CLUT (
.I0(CLBLM_L_X74Y119_SLICE_X113Y119_AO6),
.I1(CLBLM_L_X74Y119_SLICE_X112Y119_CQ),
.I2(CLBLM_L_X72Y118_SLICE_X108Y118_CQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_R_X65Y105_SLICE_X99Y105_CQ),
.I5(CLBLL_R_X75Y124_SLICE_X115Y124_BQ),
.O5(CLBLM_L_X74Y119_SLICE_X112Y119_CO5),
.O6(CLBLM_L_X74Y119_SLICE_X112Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffcccccffff)
  ) CLBLM_L_X74Y119_SLICE_X112Y119_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X65Y105_SLICE_X99Y105_CQ),
.I2(CLBLM_L_X76Y125_SLICE_X116Y125_C5Q),
.I3(CLBLM_L_X76Y122_SLICE_X116Y122_CQ),
.I4(CLBLM_L_X72Y118_SLICE_X108Y118_CQ),
.I5(1'b1),
.O5(CLBLM_L_X74Y119_SLICE_X112Y119_BO5),
.O6(CLBLM_L_X74Y119_SLICE_X112Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbfffff00000000)
  ) CLBLM_L_X74Y119_SLICE_X112Y119_ALUT (
.I0(CLBLM_L_X70Y105_SLICE_X105Y105_AQ),
.I1(CLBLL_R_X75Y122_SLICE_X115Y122_AQ),
.I2(CLBLM_L_X74Y121_SLICE_X113Y121_AQ),
.I3(CLBLM_L_X74Y119_SLICE_X112Y119_BO6),
.I4(CLBLL_R_X75Y121_SLICE_X114Y121_AQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X74Y119_SLICE_X112Y119_AO5),
.O6(CLBLM_L_X74Y119_SLICE_X112Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y119_SLICE_X113Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y119_SLICE_X113Y119_DO5),
.O6(CLBLM_L_X74Y119_SLICE_X113Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y119_SLICE_X113Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y119_SLICE_X113Y119_CO5),
.O6(CLBLM_L_X74Y119_SLICE_X113Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y119_SLICE_X113Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y119_SLICE_X113Y119_BO5),
.O6(CLBLM_L_X74Y119_SLICE_X113Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_L_X74Y119_SLICE_X113Y119_ALUT (
.I0(CLBLM_L_X70Y105_SLICE_X105Y105_AQ),
.I1(CLBLM_L_X76Y122_SLICE_X116Y122_CQ),
.I2(CLBLL_R_X75Y121_SLICE_X114Y121_AQ),
.I3(CLBLM_L_X74Y121_SLICE_X113Y121_AQ),
.I4(CLBLL_R_X75Y122_SLICE_X115Y122_AQ),
.I5(CLBLM_L_X76Y125_SLICE_X116Y125_C5Q),
.O5(CLBLM_L_X74Y119_SLICE_X113Y119_AO5),
.O6(CLBLM_L_X74Y119_SLICE_X113Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y120_SLICE_X112Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y120_SLICE_X112Y120_DO5),
.O6(CLBLM_L_X74Y120_SLICE_X112Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000ff00ff)
  ) CLBLM_L_X74Y120_SLICE_X112Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X76Y125_SLICE_X116Y125_C5Q),
.I4(1'b1),
.I5(CLBLM_L_X76Y122_SLICE_X116Y122_CQ),
.O5(CLBLM_L_X74Y120_SLICE_X112Y120_CO5),
.O6(CLBLM_L_X74Y120_SLICE_X112Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000003030303)
  ) CLBLM_L_X74Y120_SLICE_X112Y120_BLUT (
.I0(1'b1),
.I1(CLBLL_R_X75Y121_SLICE_X114Y121_AQ),
.I2(CLBLM_L_X70Y105_SLICE_X105Y105_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_R_X75Y122_SLICE_X115Y122_AQ),
.O5(CLBLM_L_X74Y120_SLICE_X112Y120_BO5),
.O6(CLBLM_L_X74Y120_SLICE_X112Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0400000005050505)
  ) CLBLM_L_X74Y120_SLICE_X112Y120_ALUT (
.I0(CLBLM_R_X65Y105_SLICE_X99Y105_CQ),
.I1(CLBLM_L_X74Y119_SLICE_X112Y119_CQ),
.I2(CLBLM_L_X72Y118_SLICE_X108Y118_CQ),
.I3(CLBLM_L_X74Y120_SLICE_X112Y120_BO6),
.I4(CLBLM_L_X74Y121_SLICE_X113Y121_AQ),
.I5(CLBLM_L_X74Y120_SLICE_X112Y120_CO6),
.O5(CLBLM_L_X74Y120_SLICE_X112Y120_AO5),
.O6(CLBLM_L_X74Y120_SLICE_X112Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y120_SLICE_X113Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y120_SLICE_X113Y120_DO5),
.O6(CLBLM_L_X74Y120_SLICE_X113Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y120_SLICE_X113Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y120_SLICE_X113Y120_CO5),
.O6(CLBLM_L_X74Y120_SLICE_X113Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y120_SLICE_X113Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y120_SLICE_X113Y120_BO5),
.O6(CLBLM_L_X74Y120_SLICE_X113Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y120_SLICE_X113Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y120_SLICE_X113Y120_AO5),
.O6(CLBLM_L_X74Y120_SLICE_X113Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y121_SLICE_X112Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y121_SLICE_X112Y121_DO5),
.O6(CLBLM_L_X74Y121_SLICE_X112Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y121_SLICE_X112Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y121_SLICE_X112Y121_CO5),
.O6(CLBLM_L_X74Y121_SLICE_X112Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y121_SLICE_X112Y121_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y121_SLICE_X112Y121_BO5),
.O6(CLBLM_L_X74Y121_SLICE_X112Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y121_SLICE_X112Y121_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y121_SLICE_X112Y121_AO5),
.O6(CLBLM_L_X74Y121_SLICE_X112Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y121_SLICE_X113Y121_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y121_SLICE_X113Y121_AO5),
.Q(CLBLM_L_X74Y121_SLICE_X113Y121_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y121_SLICE_X113Y121_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y121_SLICE_X113Y121_BO5),
.Q(CLBLM_L_X74Y121_SLICE_X113Y121_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y121_SLICE_X113Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y121_SLICE_X113Y121_AO6),
.Q(CLBLM_L_X74Y121_SLICE_X113Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y121_SLICE_X113Y121_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y121_SLICE_X113Y121_BO6),
.Q(CLBLM_L_X74Y121_SLICE_X113Y121_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y121_SLICE_X113Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y121_SLICE_X113Y121_DO5),
.O6(CLBLM_L_X74Y121_SLICE_X113Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y121_SLICE_X113Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y121_SLICE_X113Y121_CO5),
.O6(CLBLM_L_X74Y121_SLICE_X113Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3fcfc0c06cacacac)
  ) CLBLM_L_X74Y121_SLICE_X113Y121_BLUT (
.I0(CLBLM_L_X74Y121_SLICE_X113Y121_B5Q),
.I1(CLBLM_L_X74Y121_SLICE_X113Y121_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X74Y123_SLICE_X112Y123_B5Q),
.I4(CLBLM_L_X74Y121_SLICE_X113Y121_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X74Y121_SLICE_X113Y121_BO5),
.O6(CLBLM_L_X74Y121_SLICE_X113Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeeeeee55aaff00)
  ) CLBLM_L_X74Y121_SLICE_X113Y121_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X76Y122_SLICE_X116Y122_CQ),
.I2(1'b1),
.I3(CLBLM_L_X74Y123_SLICE_X112Y123_B5Q),
.I4(CLBLM_L_X74Y121_SLICE_X113Y121_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X74Y121_SLICE_X113Y121_AO5),
.O6(CLBLM_L_X74Y121_SLICE_X113Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y122_SLICE_X112Y122_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y122_SLICE_X112Y122_AO5),
.Q(CLBLM_L_X74Y122_SLICE_X112Y122_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y122_SLICE_X112Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y122_SLICE_X112Y122_AO6),
.Q(CLBLM_L_X74Y122_SLICE_X112Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y122_SLICE_X112Y122_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y122_SLICE_X112Y122_BO6),
.Q(CLBLM_L_X74Y122_SLICE_X112Y122_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y122_SLICE_X112Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y122_SLICE_X112Y122_DO5),
.O6(CLBLM_L_X74Y122_SLICE_X112Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y122_SLICE_X112Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y122_SLICE_X112Y122_CO5),
.O6(CLBLM_L_X74Y122_SLICE_X112Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffefffffffef0000)
  ) CLBLM_L_X74Y122_SLICE_X112Y122_BLUT (
.I0(CLBLM_L_X76Y130_SLICE_X116Y130_DQ),
.I1(CLBLM_L_X74Y122_SLICE_X112Y122_BQ),
.I2(CLBLM_L_X76Y125_SLICE_X117Y125_BQ),
.I3(CLBLM_L_X74Y123_SLICE_X112Y123_BQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X72Y122_SLICE_X108Y122_CQ),
.O5(CLBLM_L_X74Y122_SLICE_X112Y122_BO5),
.O6(CLBLM_L_X74Y122_SLICE_X112Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8080a0a2ff887700)
  ) CLBLM_L_X74Y122_SLICE_X112Y122_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X75Y128_SLICE_X115Y128_BO6),
.I2(CLBLM_L_X74Y122_SLICE_X112Y122_AQ),
.I3(CLBLL_R_X73Y122_SLICE_X111Y122_AQ),
.I4(CLBLM_L_X74Y122_SLICE_X112Y122_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X74Y122_SLICE_X112Y122_AO5),
.O6(CLBLM_L_X74Y122_SLICE_X112Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y122_SLICE_X113Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y122_SLICE_X113Y122_AO6),
.Q(CLBLM_L_X74Y122_SLICE_X113Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y122_SLICE_X113Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y122_SLICE_X113Y122_DO5),
.O6(CLBLM_L_X74Y122_SLICE_X113Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y122_SLICE_X113Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y122_SLICE_X113Y122_CO5),
.O6(CLBLM_L_X74Y122_SLICE_X113Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y122_SLICE_X113Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y122_SLICE_X113Y122_BO5),
.O6(CLBLM_L_X74Y122_SLICE_X113Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h78fff0f000ff0000)
  ) CLBLM_L_X74Y122_SLICE_X113Y122_ALUT (
.I0(CLBLL_R_X75Y123_SLICE_X114Y123_BQ),
.I1(CLBLM_L_X74Y123_SLICE_X113Y123_CO5),
.I2(CLBLM_L_X74Y122_SLICE_X113Y122_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X74Y123_SLICE_X113Y123_DQ),
.I5(CLBLL_R_X75Y121_SLICE_X114Y121_AO5),
.O5(CLBLM_L_X74Y122_SLICE_X113Y122_AO5),
.O6(CLBLM_L_X74Y122_SLICE_X113Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y123_SLICE_X112Y123_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y123_SLICE_X112Y123_BO5),
.Q(CLBLM_L_X74Y123_SLICE_X112Y123_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y123_SLICE_X112Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y123_SLICE_X112Y123_AO6),
.Q(CLBLM_L_X74Y123_SLICE_X112Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y123_SLICE_X112Y123_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y123_SLICE_X112Y123_BO6),
.Q(CLBLM_L_X74Y123_SLICE_X112Y123_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff7fff7fffffffff)
  ) CLBLM_L_X74Y123_SLICE_X112Y123_DLUT (
.I0(CLBLM_L_X76Y125_SLICE_X117Y125_AQ),
.I1(CLBLL_R_X75Y123_SLICE_X115Y123_DO6),
.I2(CLBLL_R_X75Y124_SLICE_X114Y124_AQ),
.I3(CLBLL_R_X77Y122_SLICE_X118Y122_CO6),
.I4(1'b1),
.I5(CLBLL_R_X75Y124_SLICE_X114Y124_BQ),
.O5(CLBLM_L_X74Y123_SLICE_X112Y123_DO5),
.O6(CLBLM_L_X74Y123_SLICE_X112Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff7fffffffffffff)
  ) CLBLM_L_X74Y123_SLICE_X112Y123_CLUT (
.I0(CLBLM_L_X76Y125_SLICE_X117Y125_AQ),
.I1(CLBLL_R_X75Y124_SLICE_X114Y124_BQ),
.I2(CLBLL_R_X75Y123_SLICE_X115Y123_DO6),
.I3(CLBLL_R_X77Y122_SLICE_X118Y122_CO6),
.I4(CLBLL_R_X75Y124_SLICE_X114Y124_AQ),
.I5(CLBLL_R_X73Y125_SLICE_X111Y125_AQ),
.O5(CLBLM_L_X74Y123_SLICE_X112Y123_CO5),
.O6(CLBLM_L_X74Y123_SLICE_X112Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h30f000f055005500)
  ) CLBLM_L_X74Y123_SLICE_X112Y123_BLUT (
.I0(CLBLM_L_X74Y123_SLICE_X112Y123_B5Q),
.I1(CLBLM_L_X74Y123_SLICE_X112Y123_CO6),
.I2(CLBLM_L_X74Y123_SLICE_X112Y123_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X74Y123_SLICE_X113Y123_AQ),
.I5(1'b1),
.O5(CLBLM_L_X74Y123_SLICE_X112Y123_BO5),
.O6(CLBLM_L_X74Y123_SLICE_X112Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h37330000b7f3c0c0)
  ) CLBLM_L_X74Y123_SLICE_X112Y123_ALUT (
.I0(CLBLM_L_X74Y123_SLICE_X112Y123_DO6),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_L_X74Y123_SLICE_X112Y123_AQ),
.I3(CLBLL_R_X73Y125_SLICE_X111Y125_AQ),
.I4(CLBLM_L_X74Y123_SLICE_X113Y123_AQ),
.I5(CLBLL_R_X77Y122_SLICE_X118Y122_CO6),
.O5(CLBLM_L_X74Y123_SLICE_X112Y123_AO5),
.O6(CLBLM_L_X74Y123_SLICE_X112Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y123_SLICE_X113Y123_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y123_SLICE_X113Y123_CO6),
.Q(CLBLM_L_X74Y123_SLICE_X113Y123_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y123_SLICE_X113Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y123_SLICE_X113Y123_AO6),
.Q(CLBLM_L_X74Y123_SLICE_X113Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y123_SLICE_X113Y123_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y123_SLICE_X113Y123_BO6),
.Q(CLBLM_L_X74Y123_SLICE_X113Y123_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y123_SLICE_X113Y123_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y123_SLICE_X113Y123_DO6),
.Q(CLBLM_L_X74Y123_SLICE_X113Y123_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h78fc78fc00cc00cc)
  ) CLBLM_L_X74Y123_SLICE_X113Y123_DLUT (
.I0(CLBLM_L_X74Y123_SLICE_X113Y123_CO5),
.I1(CLBLL_R_X75Y123_SLICE_X114Y123_BQ),
.I2(CLBLM_L_X74Y123_SLICE_X113Y123_DQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(1'b1),
.I5(CLBLL_R_X75Y121_SLICE_X114Y121_AO5),
.O5(CLBLM_L_X74Y123_SLICE_X113Y123_DO5),
.O6(CLBLM_L_X74Y123_SLICE_X113Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h30fcfc30a0000000)
  ) CLBLM_L_X74Y123_SLICE_X113Y123_CLUT (
.I0(CLBLM_L_X76Y123_SLICE_X117Y123_AQ),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_L_X74Y123_SLICE_X113Y123_BQ),
.I3(CLBLM_L_X74Y123_SLICE_X113Y123_A5Q),
.I4(CLBLL_R_X75Y113_SLICE_X114Y113_AQ),
.I5(1'b1),
.O5(CLBLM_L_X74Y123_SLICE_X113Y123_CO5),
.O6(CLBLM_L_X74Y123_SLICE_X113Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7ddd2888dddd8888)
  ) CLBLM_L_X74Y123_SLICE_X113Y123_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X74Y123_SLICE_X113Y123_BQ),
.I2(CLBLM_L_X74Y109_SLICE_X113Y109_AQ),
.I3(CLBLM_L_X76Y123_SLICE_X117Y123_AQ),
.I4(CLBLL_R_X75Y113_SLICE_X114Y113_AQ),
.I5(CLBLM_L_X74Y123_SLICE_X113Y123_A5Q),
.O5(CLBLM_L_X74Y123_SLICE_X113Y123_BO5),
.O6(CLBLM_L_X74Y123_SLICE_X113Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h50cc14cc50cc14cc)
  ) CLBLM_L_X74Y123_SLICE_X113Y123_ALUT (
.I0(CLBLL_R_X77Y122_SLICE_X118Y122_CO6),
.I1(CLBLL_R_X73Y125_SLICE_X111Y125_AQ),
.I2(CLBLM_L_X74Y123_SLICE_X113Y123_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLL_R_X75Y123_SLICE_X115Y123_BO6),
.I5(1'b1),
.O5(CLBLM_L_X74Y123_SLICE_X113Y123_AO5),
.O6(CLBLM_L_X74Y123_SLICE_X113Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y125_SLICE_X112Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y126_SLICE_X113Y126_AQ),
.Q(CLBLM_L_X74Y125_SLICE_X112Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y125_SLICE_X112Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y125_SLICE_X112Y125_DO5),
.O6(CLBLM_L_X74Y125_SLICE_X112Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y125_SLICE_X112Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y125_SLICE_X112Y125_CO5),
.O6(CLBLM_L_X74Y125_SLICE_X112Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffcfffc)
  ) CLBLM_L_X74Y125_SLICE_X112Y125_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X74Y127_SLICE_X112Y127_AQ),
.I2(CLBLM_L_X74Y125_SLICE_X112Y125_AQ),
.I3(CLBLL_R_X73Y123_SLICE_X110Y123_CQ),
.I4(1'b1),
.I5(CLBLM_L_X74Y127_SLICE_X112Y127_BQ),
.O5(CLBLM_L_X74Y125_SLICE_X112Y125_BO5),
.O6(CLBLM_L_X74Y125_SLICE_X112Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000007f80ff00)
  ) CLBLM_L_X74Y125_SLICE_X112Y125_ALUT (
.I0(CLBLL_R_X75Y123_SLICE_X115Y123_DO6),
.I1(CLBLL_R_X75Y124_SLICE_X114Y124_BQ),
.I2(CLBLM_L_X76Y125_SLICE_X117Y125_AQ),
.I3(CLBLL_R_X73Y125_SLICE_X111Y125_AQ),
.I4(CLBLL_R_X75Y124_SLICE_X114Y124_AQ),
.I5(CLBLL_R_X77Y122_SLICE_X118Y122_CO6),
.O5(CLBLM_L_X74Y125_SLICE_X112Y125_AO5),
.O6(CLBLM_L_X74Y125_SLICE_X112Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y125_SLICE_X113Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y125_SLICE_X113Y125_DO5),
.O6(CLBLM_L_X74Y125_SLICE_X113Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y125_SLICE_X113Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y125_SLICE_X113Y125_CO5),
.O6(CLBLM_L_X74Y125_SLICE_X113Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y125_SLICE_X113Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y125_SLICE_X113Y125_BO5),
.O6(CLBLM_L_X74Y125_SLICE_X113Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y125_SLICE_X113Y125_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y125_SLICE_X113Y125_AO5),
.O6(CLBLM_L_X74Y125_SLICE_X113Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y126_SLICE_X112Y126_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y126_SLICE_X112Y126_CO5),
.Q(CLBLM_L_X74Y126_SLICE_X112Y126_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y126_SLICE_X112Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y126_SLICE_X112Y126_AO6),
.Q(CLBLM_L_X74Y126_SLICE_X112Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y126_SLICE_X112Y126_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y126_SLICE_X112Y126_DO6),
.Q(CLBLM_L_X74Y126_SLICE_X112Y126_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44ee44e4e4)
  ) CLBLM_L_X74Y126_SLICE_X112Y126_DLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X74Y126_SLICE_X112Y126_AQ),
.I2(CLBLL_R_X75Y128_SLICE_X114Y128_AO6),
.I3(CLBLM_L_X74Y126_SLICE_X112Y126_DQ),
.I4(CLBLM_L_X74Y126_SLICE_X112Y126_BO5),
.I5(CLBLL_R_X75Y128_SLICE_X115Y128_AO6),
.O5(CLBLM_L_X74Y126_SLICE_X112Y126_DO5),
.O6(CLBLM_L_X74Y126_SLICE_X112Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33003300fa50d8d8)
  ) CLBLM_L_X74Y126_SLICE_X112Y126_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X74Y126_SLICE_X113Y126_AQ),
.I2(CLBLM_L_X74Y125_SLICE_X112Y125_AQ),
.I3(CLBLM_L_X74Y126_SLICE_X112Y126_A5Q),
.I4(CLBLL_R_X75Y128_SLICE_X115Y128_AO6),
.I5(1'b1),
.O5(CLBLM_L_X74Y126_SLICE_X112Y126_CO5),
.O6(CLBLM_L_X74Y126_SLICE_X112Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaffaadddddddd)
  ) CLBLM_L_X74Y126_SLICE_X112Y126_BLUT (
.I0(CLBLM_L_X74Y126_SLICE_X113Y126_A5Q),
.I1(CLBLM_L_X74Y126_SLICE_X112Y126_A5Q),
.I2(1'b1),
.I3(CLBLL_R_X75Y128_SLICE_X115Y128_AO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y126_SLICE_X112Y126_BO5),
.O6(CLBLM_L_X74Y126_SLICE_X112Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0b8fffff0b80000)
  ) CLBLM_L_X74Y126_SLICE_X112Y126_ALUT (
.I0(CLBLL_R_X75Y128_SLICE_X114Y128_AO6),
.I1(CLBLM_L_X74Y126_SLICE_X112Y126_A5Q),
.I2(CLBLM_L_X74Y126_SLICE_X112Y126_AQ),
.I3(CLBLM_L_X74Y126_SLICE_X112Y126_BO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X73Y126_SLICE_X111Y126_AQ),
.O5(CLBLM_L_X74Y126_SLICE_X112Y126_AO5),
.O6(CLBLM_L_X74Y126_SLICE_X112Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y126_SLICE_X113Y126_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y126_SLICE_X113Y126_AO5),
.Q(CLBLM_L_X74Y126_SLICE_X113Y126_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y126_SLICE_X113Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y126_SLICE_X113Y126_AO6),
.Q(CLBLM_L_X74Y126_SLICE_X113Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y126_SLICE_X113Y126_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y126_SLICE_X113Y126_BO6),
.Q(CLBLM_L_X74Y126_SLICE_X113Y126_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y126_SLICE_X113Y126_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y126_SLICE_X113Y126_CO6),
.Q(CLBLM_L_X74Y126_SLICE_X113Y126_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y126_SLICE_X113Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y126_SLICE_X113Y126_DO5),
.O6(CLBLM_L_X74Y126_SLICE_X113Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaaaacccaaaaa)
  ) CLBLM_L_X74Y126_SLICE_X113Y126_CLUT (
.I0(CLBLM_L_X74Y126_SLICE_X113Y126_BQ),
.I1(CLBLM_L_X74Y126_SLICE_X113Y126_CQ),
.I2(CLBLM_L_X74Y126_SLICE_X113Y126_AQ),
.I3(CLBLM_L_X74Y126_SLICE_X113Y126_A5Q),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X75Y128_SLICE_X115Y128_AO6),
.O5(CLBLM_L_X74Y126_SLICE_X113Y126_CO5),
.O6(CLBLM_L_X74Y126_SLICE_X113Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd77dddd882a8880)
  ) CLBLM_L_X74Y126_SLICE_X113Y126_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X74Y126_SLICE_X113Y126_BQ),
.I2(CLBLM_L_X74Y126_SLICE_X113Y126_AQ),
.I3(CLBLL_R_X75Y128_SLICE_X115Y128_AO6),
.I4(CLBLM_L_X74Y128_SLICE_X113Y128_AO6),
.I5(CLBLM_L_X74Y126_SLICE_X113Y126_A5Q),
.O5(CLBLM_L_X74Y126_SLICE_X113Y126_BO5),
.O6(CLBLM_L_X74Y126_SLICE_X113Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8080a0a2ff887700)
  ) CLBLM_L_X74Y126_SLICE_X113Y126_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X75Y128_SLICE_X115Y128_AO6),
.I2(CLBLM_L_X74Y126_SLICE_X113Y126_AQ),
.I3(CLBLM_L_X74Y126_SLICE_X112Y126_A5Q),
.I4(CLBLM_L_X74Y126_SLICE_X113Y126_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X74Y126_SLICE_X113Y126_AO5),
.O6(CLBLM_L_X74Y126_SLICE_X113Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y127_SLICE_X112Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X71Y127_SLICE_X107Y127_AQ),
.Q(CLBLM_L_X74Y127_SLICE_X112Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y127_SLICE_X112Y127_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y129_SLICE_X112Y129_AQ),
.Q(CLBLM_L_X74Y127_SLICE_X112Y127_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7755000033000000)
  ) CLBLM_L_X74Y127_SLICE_X112Y127_DLUT (
.I0(CLBLM_L_X72Y127_SLICE_X108Y127_AQ),
.I1(CLBLM_L_X72Y127_SLICE_X108Y127_A5Q),
.I2(1'b1),
.I3(CLBLM_L_X74Y127_SLICE_X113Y127_CQ),
.I4(CLBLM_L_X72Y128_SLICE_X108Y128_A5Q),
.I5(CLBLM_L_X74Y128_SLICE_X112Y128_AQ),
.O5(CLBLM_L_X74Y127_SLICE_X112Y127_DO5),
.O6(CLBLM_L_X74Y127_SLICE_X112Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000eca0eca0)
  ) CLBLM_L_X74Y127_SLICE_X112Y127_CLUT (
.I0(CLBLM_L_X72Y127_SLICE_X108Y127_AQ),
.I1(CLBLM_L_X74Y127_SLICE_X113Y127_AQ),
.I2(CLBLM_L_X74Y128_SLICE_X112Y128_DQ),
.I3(CLBLM_L_X72Y127_SLICE_X108Y127_A5Q),
.I4(1'b1),
.I5(CLBLM_L_X72Y128_SLICE_X108Y128_A5Q),
.O5(CLBLM_L_X74Y127_SLICE_X112Y127_CO5),
.O6(CLBLM_L_X74Y127_SLICE_X112Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffaaaffffaeae)
  ) CLBLM_L_X74Y127_SLICE_X112Y127_BLUT (
.I0(CLBLM_L_X74Y127_SLICE_X112Y127_DO6),
.I1(CLBLM_L_X74Y128_SLICE_X112Y128_CQ),
.I2(CLBLM_L_X72Y127_SLICE_X108Y127_AQ),
.I3(CLBLM_L_X74Y128_SLICE_X112Y128_BQ),
.I4(CLBLM_L_X74Y127_SLICE_X112Y127_CO6),
.I5(CLBLM_L_X72Y127_SLICE_X108Y127_A5Q),
.O5(CLBLM_L_X74Y127_SLICE_X112Y127_BO5),
.O6(CLBLM_L_X74Y127_SLICE_X112Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ff00fc5cac0c)
  ) CLBLM_L_X74Y127_SLICE_X112Y127_ALUT (
.I0(CLBLL_R_X75Y128_SLICE_X115Y128_DO6),
.I1(CLBLM_L_X74Y127_SLICE_X112Y127_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X74Y127_SLICE_X113Y127_A5Q),
.I4(CLBLM_L_X74Y129_SLICE_X112Y129_AQ),
.I5(1'b1),
.O5(CLBLM_L_X74Y127_SLICE_X112Y127_AO5),
.O6(CLBLM_L_X74Y127_SLICE_X112Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y127_SLICE_X113Y127_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y127_SLICE_X112Y127_AO5),
.Q(CLBLM_L_X74Y127_SLICE_X113Y127_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y127_SLICE_X113Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y127_SLICE_X113Y127_AO6),
.Q(CLBLM_L_X74Y127_SLICE_X113Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y127_SLICE_X113Y127_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y127_SLICE_X113Y127_CO6),
.Q(CLBLM_L_X74Y127_SLICE_X113Y127_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y127_SLICE_X113Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y127_SLICE_X113Y127_DO5),
.O6(CLBLM_L_X74Y127_SLICE_X113Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88df8add88d580)
  ) CLBLM_L_X74Y127_SLICE_X113Y127_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X74Y127_SLICE_X113Y127_CQ),
.I2(CLBLL_R_X75Y128_SLICE_X115Y128_DO6),
.I3(CLBLM_L_X74Y127_SLICE_X113Y127_AQ),
.I4(CLBLM_L_X74Y127_SLICE_X113Y127_BO5),
.I5(CLBLL_R_X75Y128_SLICE_X114Y128_DO6),
.O5(CLBLM_L_X74Y127_SLICE_X113Y127_CO5),
.O6(CLBLM_L_X74Y127_SLICE_X113Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaffaaccffccff)
  ) CLBLM_L_X74Y127_SLICE_X113Y127_BLUT (
.I0(CLBLL_R_X75Y128_SLICE_X115Y128_DO6),
.I1(CLBLM_L_X74Y127_SLICE_X113Y127_A5Q),
.I2(1'b1),
.I3(CLBLM_L_X74Y129_SLICE_X112Y129_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y127_SLICE_X113Y127_BO5),
.O6(CLBLM_L_X74Y127_SLICE_X113Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0ccccaaaacccc)
  ) CLBLM_L_X74Y127_SLICE_X113Y127_ALUT (
.I0(CLBLM_L_X74Y127_SLICE_X113Y127_AQ),
.I1(CLBLM_L_X74Y128_SLICE_X112Y128_AQ),
.I2(CLBLL_R_X75Y128_SLICE_X114Y128_DO6),
.I3(CLBLM_L_X74Y127_SLICE_X113Y127_BO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X74Y127_SLICE_X113Y127_A5Q),
.O5(CLBLM_L_X74Y127_SLICE_X113Y127_AO5),
.O6(CLBLM_L_X74Y127_SLICE_X113Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y128_SLICE_X112Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y128_SLICE_X112Y128_AO6),
.Q(CLBLM_L_X74Y128_SLICE_X112Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y128_SLICE_X112Y128_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y128_SLICE_X112Y128_BO6),
.Q(CLBLM_L_X74Y128_SLICE_X112Y128_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y128_SLICE_X112Y128_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y128_SLICE_X112Y128_CO6),
.Q(CLBLM_L_X74Y128_SLICE_X112Y128_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y128_SLICE_X112Y128_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y128_SLICE_X112Y128_DO6),
.Q(CLBLM_L_X74Y128_SLICE_X112Y128_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he4eee4e4e444e4e4)
  ) CLBLM_L_X74Y128_SLICE_X112Y128_DLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X74Y127_SLICE_X113Y127_CQ),
.I2(CLBLM_L_X74Y128_SLICE_X112Y128_DQ),
.I3(CLBLL_R_X75Y128_SLICE_X115Y128_DO6),
.I4(CLBLM_L_X74Y127_SLICE_X112Y127_AO6),
.I5(CLBLL_R_X75Y128_SLICE_X114Y128_DO6),
.O5(CLBLM_L_X74Y128_SLICE_X112Y128_DO5),
.O6(CLBLM_L_X74Y128_SLICE_X112Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaeeaa22f0f0f0f0)
  ) CLBLM_L_X74Y128_SLICE_X112Y128_CLUT (
.I0(CLBLM_L_X74Y128_SLICE_X112Y128_CQ),
.I1(CLBLM_L_X74Y129_SLICE_X112Y129_A5Q),
.I2(CLBLM_L_X74Y128_SLICE_X112Y128_DQ),
.I3(CLBLM_L_X74Y128_SLICE_X113Y128_BO6),
.I4(CLBLL_R_X75Y128_SLICE_X114Y128_DO6),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X74Y128_SLICE_X112Y128_CO5),
.O6(CLBLM_L_X74Y128_SLICE_X112Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacffffacac0000)
  ) CLBLM_L_X74Y128_SLICE_X112Y128_BLUT (
.I0(CLBLL_R_X75Y128_SLICE_X114Y128_DO6),
.I1(CLBLM_L_X74Y128_SLICE_X112Y128_BQ),
.I2(CLBLM_L_X74Y128_SLICE_X113Y128_BO5),
.I3(1'b1),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X74Y128_SLICE_X113Y128_CQ),
.O5(CLBLM_L_X74Y128_SLICE_X112Y128_BO5),
.O6(CLBLM_L_X74Y128_SLICE_X112Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ccccf0aacccc)
  ) CLBLM_L_X74Y128_SLICE_X112Y128_ALUT (
.I0(CLBLL_R_X75Y128_SLICE_X114Y128_DO6),
.I1(CLBLM_L_X74Y128_SLICE_X112Y128_BQ),
.I2(CLBLM_L_X74Y128_SLICE_X112Y128_AQ),
.I3(CLBLM_L_X74Y127_SLICE_X113Y127_A5Q),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X74Y128_SLICE_X113Y128_BO6),
.O5(CLBLM_L_X74Y128_SLICE_X112Y128_AO5),
.O6(CLBLM_L_X74Y128_SLICE_X112Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y128_SLICE_X113Y128_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y128_SLICE_X113Y128_CO6),
.Q(CLBLM_L_X74Y128_SLICE_X113Y128_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y128_SLICE_X113Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y128_SLICE_X113Y128_DO5),
.O6(CLBLM_L_X74Y128_SLICE_X113Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0cfdfc080)
  ) CLBLM_L_X74Y128_SLICE_X113Y128_CLUT (
.I0(CLBLM_L_X74Y129_SLICE_X112Y129_AQ),
.I1(CLBLM_L_X74Y128_SLICE_X113Y128_CQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLL_R_X75Y128_SLICE_X115Y128_DO6),
.I4(CLBLM_L_X74Y129_SLICE_X113Y129_AQ),
.I5(CLBLM_L_X74Y129_SLICE_X112Y129_A5Q),
.O5(CLBLM_L_X74Y128_SLICE_X113Y128_CO5),
.O6(CLBLM_L_X74Y128_SLICE_X113Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaffff00000505)
  ) CLBLM_L_X74Y128_SLICE_X113Y128_BLUT (
.I0(CLBLL_R_X75Y128_SLICE_X115Y128_DO6),
.I1(1'b1),
.I2(CLBLM_L_X74Y129_SLICE_X112Y129_A5Q),
.I3(1'b1),
.I4(CLBLM_L_X74Y129_SLICE_X112Y129_AQ),
.I5(1'b1),
.O5(CLBLM_L_X74Y128_SLICE_X113Y128_BO5),
.O6(CLBLM_L_X74Y128_SLICE_X113Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeeeefdfdfdfd)
  ) CLBLM_L_X74Y128_SLICE_X113Y128_ALUT (
.I0(CLBLL_R_X77Y128_SLICE_X118Y128_B5Q),
.I1(CLBLM_L_X74Y129_SLICE_X113Y129_CO6),
.I2(CLBLL_R_X75Y130_SLICE_X115Y130_AQ),
.I3(1'b1),
.I4(CLBLL_R_X75Y129_SLICE_X114Y129_DQ),
.I5(1'b1),
.O5(CLBLM_L_X74Y128_SLICE_X113Y128_AO5),
.O6(CLBLM_L_X74Y128_SLICE_X113Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y129_SLICE_X112Y129_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y129_SLICE_X112Y129_AO5),
.Q(CLBLM_L_X74Y129_SLICE_X112Y129_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y129_SLICE_X112Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y129_SLICE_X112Y129_AO6),
.Q(CLBLM_L_X74Y129_SLICE_X112Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y129_SLICE_X112Y129_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y133_SLICE_X114Y133_AQ),
.Q(CLBLM_L_X74Y129_SLICE_X112Y129_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y129_SLICE_X112Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y129_SLICE_X112Y129_DO5),
.O6(CLBLM_L_X74Y129_SLICE_X112Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y129_SLICE_X112Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y129_SLICE_X112Y129_CO5),
.O6(CLBLM_L_X74Y129_SLICE_X112Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y129_SLICE_X112Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y129_SLICE_X112Y129_BO5),
.O6(CLBLM_L_X74Y129_SLICE_X112Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha000a0a2eecc44cc)
  ) CLBLM_L_X74Y129_SLICE_X112Y129_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X74Y127_SLICE_X113Y127_A5Q),
.I2(CLBLM_L_X74Y129_SLICE_X112Y129_AQ),
.I3(CLBLL_R_X75Y128_SLICE_X115Y128_DO6),
.I4(CLBLM_L_X74Y129_SLICE_X112Y129_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X74Y129_SLICE_X112Y129_AO5),
.O6(CLBLM_L_X74Y129_SLICE_X112Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y129_SLICE_X113Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y129_SLICE_X113Y129_AO6),
.Q(CLBLM_L_X74Y129_SLICE_X113Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y129_SLICE_X113Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y129_SLICE_X113Y129_DO5),
.O6(CLBLM_L_X74Y129_SLICE_X113Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5f5fffff5fff)
  ) CLBLM_L_X74Y129_SLICE_X113Y129_CLUT (
.I0(CLBLL_R_X77Y129_SLICE_X119Y129_BQ),
.I1(1'b1),
.I2(CLBLM_L_X76Y125_SLICE_X117Y125_BQ),
.I3(CLBLM_L_X78Y131_SLICE_X120Y131_AQ),
.I4(CLBLM_L_X76Y130_SLICE_X116Y130_DQ),
.I5(CLBLL_R_X77Y130_SLICE_X118Y130_AQ),
.O5(CLBLM_L_X74Y129_SLICE_X113Y129_CO5),
.O6(CLBLM_L_X74Y129_SLICE_X113Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff5d5f0c0f0c0)
  ) CLBLM_L_X74Y129_SLICE_X113Y129_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X78Y131_SLICE_X120Y131_AQ),
.I2(CLBLL_R_X77Y129_SLICE_X119Y129_BQ),
.I3(CLBLL_R_X77Y130_SLICE_X118Y130_AQ),
.I4(CLBLL_R_X73Y132_SLICE_X111Y132_AO6),
.I5(1'b1),
.O5(CLBLM_L_X74Y129_SLICE_X113Y129_BO5),
.O6(CLBLM_L_X74Y129_SLICE_X113Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8fadaf872507250)
  ) CLBLM_L_X74Y129_SLICE_X113Y129_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X75Y128_SLICE_X115Y128_DO6),
.I2(CLBLM_L_X74Y129_SLICE_X112Y129_A5Q),
.I3(CLBLL_R_X75Y128_SLICE_X114Y128_DO5),
.I4(CLBLM_L_X74Y129_SLICE_X112Y129_AQ),
.I5(CLBLM_L_X74Y129_SLICE_X113Y129_AQ),
.O5(CLBLM_L_X74Y129_SLICE_X113Y129_AO5),
.O6(CLBLM_L_X74Y129_SLICE_X113Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y131_SLICE_X112Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X73Y131_SLICE_X111Y131_AQ),
.Q(CLBLM_L_X74Y131_SLICE_X112Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y131_SLICE_X112Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y131_SLICE_X112Y131_DO5),
.O6(CLBLM_L_X74Y131_SLICE_X112Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y131_SLICE_X112Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y131_SLICE_X112Y131_CO5),
.O6(CLBLM_L_X74Y131_SLICE_X112Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y131_SLICE_X112Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y131_SLICE_X112Y131_BO5),
.O6(CLBLM_L_X74Y131_SLICE_X112Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y131_SLICE_X112Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y131_SLICE_X112Y131_AO5),
.O6(CLBLM_L_X74Y131_SLICE_X112Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y131_SLICE_X113Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y131_SLICE_X113Y131_DO5),
.O6(CLBLM_L_X74Y131_SLICE_X113Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y131_SLICE_X113Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y131_SLICE_X113Y131_CO5),
.O6(CLBLM_L_X74Y131_SLICE_X113Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y131_SLICE_X113Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y131_SLICE_X113Y131_BO5),
.O6(CLBLM_L_X74Y131_SLICE_X113Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y131_SLICE_X113Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y131_SLICE_X113Y131_AO5),
.O6(CLBLM_L_X74Y131_SLICE_X113Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y132_SLICE_X112Y132_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y132_SLICE_X112Y132_BO5),
.Q(CLBLM_L_X74Y132_SLICE_X112Y132_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y132_SLICE_X112Y132_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y132_SLICE_X112Y132_CO5),
.Q(CLBLM_L_X74Y132_SLICE_X112Y132_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y132_SLICE_X112Y132_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y132_SLICE_X112Y132_AO6),
.Q(CLBLM_L_X74Y132_SLICE_X112Y132_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y132_SLICE_X112Y132_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y132_SLICE_X112Y132_CO6),
.Q(CLBLM_L_X74Y132_SLICE_X112Y132_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y132_SLICE_X112Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y132_SLICE_X112Y132_DO5),
.O6(CLBLM_L_X74Y132_SLICE_X112Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc30fc30ee22ee22)
  ) CLBLM_L_X74Y132_SLICE_X112Y132_CLUT (
.I0(CLBLM_L_X74Y131_SLICE_X112Y131_AQ),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLL_R_X73Y131_SLICE_X110Y131_AQ),
.I3(CLBLM_L_X70Y136_SLICE_X105Y136_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y132_SLICE_X112Y132_CO5),
.O6(CLBLM_L_X74Y132_SLICE_X112Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000f0f7f000c00)
  ) CLBLM_L_X74Y132_SLICE_X112Y132_BLUT (
.I0(CLBLM_L_X74Y134_SLICE_X113Y134_BQ),
.I1(CLBLM_L_X74Y133_SLICE_X112Y133_DO5),
.I2(CLBLM_L_X74Y132_SLICE_X112Y132_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X74Y132_SLICE_X112Y132_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X74Y132_SLICE_X112Y132_BO5),
.O6(CLBLM_L_X74Y132_SLICE_X112Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0e2f0aaaaaaaa)
  ) CLBLM_L_X74Y132_SLICE_X112Y132_ALUT (
.I0(CLBLM_L_X74Y134_SLICE_X113Y134_BQ),
.I1(CLBLM_L_X74Y134_SLICE_X113Y134_CQ),
.I2(CLBLM_L_X74Y132_SLICE_X112Y132_AQ),
.I3(CLBLM_L_X74Y129_SLICE_X112Y129_BQ),
.I4(CLBLM_L_X74Y134_SLICE_X113Y134_A5Q),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X74Y132_SLICE_X112Y132_AO5),
.O6(CLBLM_L_X74Y132_SLICE_X112Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y132_SLICE_X113Y132_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y132_SLICE_X113Y132_AO6),
.Q(CLBLM_L_X74Y132_SLICE_X113Y132_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y132_SLICE_X113Y132_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y132_SLICE_X113Y132_BO6),
.Q(CLBLM_L_X74Y132_SLICE_X113Y132_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y132_SLICE_X113Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y132_SLICE_X113Y132_DO5),
.O6(CLBLM_L_X74Y132_SLICE_X113Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffffffef)
  ) CLBLM_L_X74Y132_SLICE_X113Y132_CLUT (
.I0(CLBLM_L_X74Y132_SLICE_X112Y132_AQ),
.I1(CLBLM_L_X74Y132_SLICE_X112Y132_A5Q),
.I2(CLBLM_L_X74Y129_SLICE_X112Y129_BQ),
.I3(CLBLM_L_X74Y134_SLICE_X113Y134_A5Q),
.I4(CLBLM_L_X74Y134_SLICE_X113Y134_CQ),
.I5(CLBLM_L_X74Y132_SLICE_X113Y132_AQ),
.O5(CLBLM_L_X74Y132_SLICE_X113Y132_CO5),
.O6(CLBLM_L_X74Y132_SLICE_X113Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc6cccccf0f0f0f0)
  ) CLBLM_L_X74Y132_SLICE_X113Y132_BLUT (
.I0(CLBLM_L_X74Y133_SLICE_X112Y133_DO5),
.I1(CLBLM_L_X74Y132_SLICE_X113Y132_BQ),
.I2(CLBLM_L_X74Y132_SLICE_X113Y132_AQ),
.I3(CLBLM_L_X74Y134_SLICE_X113Y134_BQ),
.I4(CLBLM_L_X74Y132_SLICE_X112Y132_AQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X74Y132_SLICE_X113Y132_BO5),
.O6(CLBLM_L_X74Y132_SLICE_X113Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a0a0a3afacafa)
  ) CLBLM_L_X74Y132_SLICE_X113Y132_ALUT (
.I0(CLBLM_L_X74Y133_SLICE_X112Y133_CQ),
.I1(CLBLM_L_X74Y133_SLICE_X113Y133_AO6),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X74Y133_SLICE_X112Y133_DO5),
.I4(CLBLM_L_X74Y132_SLICE_X113Y132_BQ),
.I5(CLBLM_L_X74Y132_SLICE_X113Y132_CO6),
.O5(CLBLM_L_X74Y132_SLICE_X113Y132_AO5),
.O6(CLBLM_L_X74Y132_SLICE_X113Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y133_SLICE_X112Y133_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y133_SLICE_X112Y133_AO6),
.Q(CLBLM_L_X74Y133_SLICE_X112Y133_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y133_SLICE_X112Y133_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y133_SLICE_X112Y133_BO6),
.Q(CLBLM_L_X74Y133_SLICE_X112Y133_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y133_SLICE_X112Y133_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y133_SLICE_X112Y133_CO6),
.Q(CLBLM_L_X74Y133_SLICE_X112Y133_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800880000220022)
  ) CLBLM_L_X74Y133_SLICE_X112Y133_DLUT (
.I0(CLBLM_L_X74Y129_SLICE_X112Y129_BQ),
.I1(CLBLM_L_X74Y134_SLICE_X113Y134_A5Q),
.I2(1'b1),
.I3(CLBLM_L_X74Y134_SLICE_X113Y134_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y133_SLICE_X112Y133_DO5),
.O6(CLBLM_L_X74Y133_SLICE_X112Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdff0fff02f000f00)
  ) CLBLM_L_X74Y133_SLICE_X112Y133_CLUT (
.I0(CLBLM_L_X74Y132_SLICE_X112Y132_AQ),
.I1(CLBLM_L_X74Y134_SLICE_X113Y134_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X74Y133_SLICE_X112Y133_BQ),
.I4(CLBLM_L_X74Y133_SLICE_X112Y133_DO6),
.I5(CLBLM_L_X74Y133_SLICE_X112Y133_CQ),
.O5(CLBLM_L_X74Y133_SLICE_X112Y133_CO5),
.O6(CLBLM_L_X74Y133_SLICE_X112Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeccf0f04444f0f0)
  ) CLBLM_L_X74Y133_SLICE_X112Y133_BLUT (
.I0(CLBLM_L_X74Y133_SLICE_X112Y133_DO6),
.I1(CLBLM_L_X74Y133_SLICE_X112Y133_BQ),
.I2(CLBLM_L_X74Y133_SLICE_X112Y133_AQ),
.I3(CLBLM_L_X74Y132_SLICE_X112Y132_BO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X74Y133_SLICE_X113Y133_AO5),
.O5(CLBLM_L_X74Y133_SLICE_X112Y133_BO5),
.O6(CLBLM_L_X74Y133_SLICE_X112Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd2fff0fff000f000)
  ) CLBLM_L_X74Y133_SLICE_X112Y133_ALUT (
.I0(CLBLM_L_X74Y134_SLICE_X112Y134_AO5),
.I1(CLBLM_L_X74Y134_SLICE_X113Y134_BQ),
.I2(CLBLM_L_X74Y133_SLICE_X112Y133_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X74Y132_SLICE_X112Y132_AQ),
.I5(CLBLL_R_X73Y133_SLICE_X111Y133_AQ),
.O5(CLBLM_L_X74Y133_SLICE_X112Y133_AO5),
.O6(CLBLM_L_X74Y133_SLICE_X112Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y133_SLICE_X113Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y133_SLICE_X113Y133_DO5),
.O6(CLBLM_L_X74Y133_SLICE_X113Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y133_SLICE_X113Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y133_SLICE_X113Y133_CO5),
.O6(CLBLM_L_X74Y133_SLICE_X113Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y133_SLICE_X113Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y133_SLICE_X113Y133_BO5),
.O6(CLBLM_L_X74Y133_SLICE_X113Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h32003200cdff3200)
  ) CLBLM_L_X74Y133_SLICE_X113Y133_ALUT (
.I0(CLBLM_L_X76Y133_SLICE_X116Y133_BQ),
.I1(CLBLL_R_X73Y133_SLICE_X110Y133_CQ),
.I2(CLBLL_R_X75Y133_SLICE_X115Y133_AQ),
.I3(CLBLM_L_X74Y135_SLICE_X113Y135_BQ),
.I4(CLBLM_L_X74Y133_SLICE_X112Y133_CQ),
.I5(1'b1),
.O5(CLBLM_L_X74Y133_SLICE_X113Y133_AO5),
.O6(CLBLM_L_X74Y133_SLICE_X113Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y134_SLICE_X112Y134_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y134_SLICE_X112Y134_BO6),
.Q(CLBLM_L_X74Y134_SLICE_X112Y134_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y134_SLICE_X112Y134_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y134_SLICE_X112Y134_CO6),
.Q(CLBLM_L_X74Y134_SLICE_X112Y134_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y134_SLICE_X112Y134_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y134_SLICE_X112Y134_DO6),
.Q(CLBLM_L_X74Y134_SLICE_X112Y134_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8f0f0ff00ff00)
  ) CLBLM_L_X74Y134_SLICE_X112Y134_DLUT (
.I0(CLBLM_L_X74Y134_SLICE_X113Y134_DO5),
.I1(CLBLM_L_X74Y132_SLICE_X112Y132_C5Q),
.I2(CLBLM_L_X74Y134_SLICE_X112Y134_DQ),
.I3(CLBLM_L_X74Y134_SLICE_X112Y134_BQ),
.I4(CLBLM_L_X74Y134_SLICE_X113Y134_A5Q),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X74Y134_SLICE_X112Y134_DO5),
.O6(CLBLM_L_X74Y134_SLICE_X112Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc00ccf0f0f0f0)
  ) CLBLM_L_X74Y134_SLICE_X112Y134_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X74Y134_SLICE_X112Y134_CQ),
.I2(CLBLM_L_X74Y134_SLICE_X112Y134_DQ),
.I3(CLBLL_R_X75Y133_SLICE_X114Y133_BQ),
.I4(CLBLM_L_X74Y134_SLICE_X112Y134_BQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X74Y134_SLICE_X112Y134_CO5),
.O6(CLBLM_L_X74Y134_SLICE_X112Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaaccf0f0f0f0)
  ) CLBLM_L_X74Y134_SLICE_X112Y134_BLUT (
.I0(CLBLM_L_X74Y132_SLICE_X112Y132_C5Q),
.I1(CLBLM_L_X74Y134_SLICE_X112Y134_BQ),
.I2(CLBLM_L_X74Y134_SLICE_X113Y134_A5Q),
.I3(CLBLL_R_X75Y133_SLICE_X114Y133_BQ),
.I4(1'b1),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X74Y134_SLICE_X112Y134_BO5),
.O6(CLBLM_L_X74Y134_SLICE_X112Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4400440022002200)
  ) CLBLM_L_X74Y134_SLICE_X112Y134_ALUT (
.I0(CLBLM_L_X74Y134_SLICE_X113Y134_A5Q),
.I1(CLBLM_L_X74Y134_SLICE_X113Y134_CQ),
.I2(1'b1),
.I3(CLBLM_L_X74Y129_SLICE_X112Y129_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y134_SLICE_X112Y134_AO5),
.O6(CLBLM_L_X74Y134_SLICE_X112Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y134_SLICE_X113Y134_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y134_SLICE_X113Y134_DO6),
.Q(CLBLM_L_X74Y134_SLICE_X113Y134_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y134_SLICE_X113Y134_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y134_SLICE_X113Y134_AO6),
.Q(CLBLM_L_X74Y134_SLICE_X113Y134_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y134_SLICE_X113Y134_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y134_SLICE_X113Y134_BO6),
.Q(CLBLM_L_X74Y134_SLICE_X113Y134_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y134_SLICE_X113Y134_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y134_SLICE_X113Y134_CO6),
.Q(CLBLM_L_X74Y134_SLICE_X113Y134_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3fcfaa0acccc0000)
  ) CLBLM_L_X74Y134_SLICE_X113Y134_DLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X75Y133_SLICE_X114Y133_BQ),
.I2(CLBLM_L_X74Y135_SLICE_X113Y135_DO6),
.I3(CLBLM_L_X74Y134_SLICE_X113Y134_A5Q),
.I4(CLBLM_L_X74Y134_SLICE_X113Y134_CQ),
.I5(1'b1),
.O5(CLBLM_L_X74Y134_SLICE_X113Y134_DO5),
.O6(CLBLM_L_X74Y134_SLICE_X113Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h22a82288aaaa2288)
  ) CLBLM_L_X74Y134_SLICE_X113Y134_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X74Y134_SLICE_X113Y134_CQ),
.I2(CLBLM_L_X74Y134_SLICE_X113Y134_A5Q),
.I3(CLBLL_R_X75Y133_SLICE_X114Y133_BQ),
.I4(CLBLL_R_X75Y134_SLICE_X115Y134_CO6),
.I5(CLBLM_L_X74Y135_SLICE_X113Y135_BQ),
.O5(CLBLM_L_X74Y134_SLICE_X113Y134_CO5),
.O6(CLBLM_L_X74Y134_SLICE_X113Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfdfcfcfc080c0c0)
  ) CLBLM_L_X74Y134_SLICE_X113Y134_BLUT (
.I0(CLBLM_L_X74Y134_SLICE_X113Y134_CQ),
.I1(CLBLM_L_X74Y134_SLICE_X113Y134_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X74Y134_SLICE_X113Y134_A5Q),
.I4(CLBLM_L_X74Y129_SLICE_X112Y129_BQ),
.I5(CLBLM_L_X74Y132_SLICE_X112Y132_A5Q),
.O5(CLBLM_L_X74Y134_SLICE_X113Y134_BO5),
.O6(CLBLM_L_X74Y134_SLICE_X113Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h9affaaffaa00aa00)
  ) CLBLM_L_X74Y134_SLICE_X113Y134_ALUT (
.I0(CLBLM_L_X74Y134_SLICE_X113Y134_AQ),
.I1(CLBLM_L_X74Y134_SLICE_X113Y134_BQ),
.I2(CLBLM_L_X74Y134_SLICE_X112Y134_AO6),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X74Y132_SLICE_X112Y132_AQ),
.I5(CLBLL_R_X73Y134_SLICE_X111Y134_AQ),
.O5(CLBLM_L_X74Y134_SLICE_X113Y134_AO5),
.O6(CLBLM_L_X74Y134_SLICE_X113Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y135_SLICE_X112Y135_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y135_SLICE_X112Y135_AO6),
.Q(CLBLM_L_X74Y135_SLICE_X112Y135_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y135_SLICE_X112Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y135_SLICE_X112Y135_DO5),
.O6(CLBLM_L_X74Y135_SLICE_X112Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y135_SLICE_X112Y135_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y135_SLICE_X112Y135_CO5),
.O6(CLBLM_L_X74Y135_SLICE_X112Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd0f0000000000000)
  ) CLBLM_L_X74Y135_SLICE_X112Y135_BLUT (
.I0(CLBLM_L_X74Y132_SLICE_X112Y132_C5Q),
.I1(CLBLM_L_X74Y134_SLICE_X112Y134_CQ),
.I2(CLBLM_L_X74Y135_SLICE_X112Y135_AQ),
.I3(CLBLM_L_X74Y134_SLICE_X112Y134_BQ),
.I4(CLBLL_R_X73Y134_SLICE_X110Y134_AO6),
.I5(CLBLL_R_X75Y133_SLICE_X114Y133_BQ),
.O5(CLBLM_L_X74Y135_SLICE_X112Y135_BO5),
.O6(CLBLM_L_X74Y135_SLICE_X112Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4848ff484848ff48)
  ) CLBLM_L_X74Y135_SLICE_X112Y135_ALUT (
.I0(CLBLM_L_X74Y135_SLICE_X113Y135_CO6),
.I1(CLBLM_L_X74Y135_SLICE_X113Y135_DO6),
.I2(CLBLM_L_X74Y135_SLICE_X112Y135_AQ),
.I3(CLBLM_L_X74Y135_SLICE_X113Y135_BQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLM_L_X74Y135_SLICE_X112Y135_AO5),
.O6(CLBLM_L_X74Y135_SLICE_X112Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y135_SLICE_X113Y135_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y135_SLICE_X113Y135_AO6),
.Q(CLBLM_L_X74Y135_SLICE_X113Y135_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X74Y135_SLICE_X113Y135_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X74Y135_SLICE_X113Y135_BO6),
.Q(CLBLM_L_X74Y135_SLICE_X113Y135_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3737300000000)
  ) CLBLM_L_X74Y135_SLICE_X113Y135_DLUT (
.I0(CLBLM_L_X74Y134_SLICE_X113Y134_A5Q),
.I1(CLBLL_R_X75Y134_SLICE_X115Y134_CO6),
.I2(CLBLM_L_X74Y135_SLICE_X113Y135_BQ),
.I3(1'b1),
.I4(CLBLM_L_X74Y134_SLICE_X113Y134_CQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X74Y135_SLICE_X113Y135_DO5),
.O6(CLBLM_L_X74Y135_SLICE_X113Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2200220002002200)
  ) CLBLM_L_X74Y135_SLICE_X113Y135_CLUT (
.I0(CLBLM_L_X74Y134_SLICE_X113Y134_A5Q),
.I1(CLBLM_L_X74Y134_SLICE_X113Y134_CQ),
.I2(CLBLM_L_X74Y132_SLICE_X112Y132_C5Q),
.I3(CLBLL_R_X75Y133_SLICE_X114Y133_BQ),
.I4(CLBLM_L_X74Y134_SLICE_X112Y134_BQ),
.I5(CLBLM_L_X74Y134_SLICE_X112Y134_CQ),
.O5(CLBLM_L_X74Y135_SLICE_X113Y135_CO5),
.O6(CLBLM_L_X74Y135_SLICE_X113Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f7f2a2aff55aa00)
  ) CLBLM_L_X74Y135_SLICE_X113Y135_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X74Y135_SLICE_X112Y135_BO6),
.I2(CLBLM_L_X74Y135_SLICE_X113Y135_AQ),
.I3(CLBLL_R_X75Y134_SLICE_X115Y134_CO6),
.I4(CLBLM_L_X74Y134_SLICE_X112Y134_CQ),
.I5(CLBLM_L_X74Y135_SLICE_X113Y135_BQ),
.O5(CLBLM_L_X74Y135_SLICE_X113Y135_BO5),
.O6(CLBLM_L_X74Y135_SLICE_X113Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3b3ba0a0b3b3a0a0)
  ) CLBLM_L_X74Y135_SLICE_X113Y135_ALUT (
.I0(CLBLM_L_X74Y135_SLICE_X113Y135_DO6),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_L_X74Y135_SLICE_X113Y135_AQ),
.I3(1'b1),
.I4(CLBLM_L_X74Y135_SLICE_X112Y135_AQ),
.I5(CLBLM_L_X74Y135_SLICE_X113Y135_CO6),
.O5(CLBLM_L_X74Y135_SLICE_X113Y135_AO5),
.O6(CLBLM_L_X74Y135_SLICE_X113Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y109_SLICE_X116Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y109_SLICE_X116Y109_DO5),
.O6(CLBLM_L_X76Y109_SLICE_X116Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y109_SLICE_X116Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y109_SLICE_X116Y109_CO5),
.O6(CLBLM_L_X76Y109_SLICE_X116Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y109_SLICE_X116Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y109_SLICE_X116Y109_BO5),
.O6(CLBLM_L_X76Y109_SLICE_X116Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00ff00ff)
  ) CLBLM_L_X76Y109_SLICE_X116Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y109_SLICE_X116Y109_AO5),
.O6(CLBLM_L_X76Y109_SLICE_X116Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y109_SLICE_X117Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y109_SLICE_X117Y109_DO5),
.O6(CLBLM_L_X76Y109_SLICE_X117Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y109_SLICE_X117Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y109_SLICE_X117Y109_CO5),
.O6(CLBLM_L_X76Y109_SLICE_X117Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y109_SLICE_X117Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y109_SLICE_X117Y109_BO5),
.O6(CLBLM_L_X76Y109_SLICE_X117Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y109_SLICE_X117Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y109_SLICE_X117Y109_AO5),
.O6(CLBLM_L_X76Y109_SLICE_X117Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y111_SLICE_X116Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y111_SLICE_X98Y111_AQ),
.Q(CLBLM_L_X76Y111_SLICE_X116Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y111_SLICE_X116Y111_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y99_SLICE_X93Y99_AQ),
.Q(CLBLM_L_X76Y111_SLICE_X116Y111_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y111_SLICE_X116Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y111_SLICE_X116Y111_DO5),
.O6(CLBLM_L_X76Y111_SLICE_X116Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y111_SLICE_X116Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y111_SLICE_X116Y111_CO5),
.O6(CLBLM_L_X76Y111_SLICE_X116Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y111_SLICE_X116Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y111_SLICE_X116Y111_BO5),
.O6(CLBLM_L_X76Y111_SLICE_X116Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y111_SLICE_X116Y111_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y111_SLICE_X116Y111_AO5),
.O6(CLBLM_L_X76Y111_SLICE_X116Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y111_SLICE_X117Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y111_SLICE_X117Y111_DO5),
.O6(CLBLM_L_X76Y111_SLICE_X117Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y111_SLICE_X117Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y111_SLICE_X117Y111_CO5),
.O6(CLBLM_L_X76Y111_SLICE_X117Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y111_SLICE_X117Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y111_SLICE_X117Y111_BO5),
.O6(CLBLM_L_X76Y111_SLICE_X117Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y111_SLICE_X117Y111_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y111_SLICE_X117Y111_AO5),
.O6(CLBLM_L_X76Y111_SLICE_X117Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y118_SLICE_X116Y118_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y118_SLICE_X116Y118_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y118_SLICE_X116Y118_BQ),
.Q(CLBLM_L_X76Y118_SLICE_X116Y118_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y118_SLICE_X116Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y118_SLICE_X116Y118_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y118_SLICE_X116Y118_AO5),
.Q(CLBLM_L_X76Y118_SLICE_X116Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y118_SLICE_X116Y118_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y118_SLICE_X116Y118_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y118_SLICE_X116Y118_DQ),
.Q(CLBLM_L_X76Y118_SLICE_X116Y118_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y118_SLICE_X116Y118_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y118_SLICE_X116Y118_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y119_SLICE_X116Y119_A5Q),
.Q(CLBLM_L_X76Y118_SLICE_X116Y118_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y118_SLICE_X116Y118_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y118_SLICE_X116Y118_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y118_SLICE_X116Y118_AQ),
.Q(CLBLM_L_X76Y118_SLICE_X116Y118_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y118_SLICE_X116Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y118_SLICE_X116Y118_DO5),
.O6(CLBLM_L_X76Y118_SLICE_X116Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y118_SLICE_X116Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y118_SLICE_X116Y118_CO5),
.O6(CLBLM_L_X76Y118_SLICE_X116Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffbfffffffefff)
  ) CLBLM_L_X76Y118_SLICE_X116Y118_BLUT (
.I0(CLBLM_L_X76Y119_SLICE_X116Y119_A5Q),
.I1(CLBLM_L_X76Y118_SLICE_X116Y118_BQ),
.I2(CLBLM_L_X76Y118_SLICE_X116Y118_CQ),
.I3(CLBLM_L_X76Y118_SLICE_X117Y118_BQ),
.I4(CLBLM_L_X76Y118_SLICE_X117Y118_AQ),
.I5(CLBLM_L_X76Y118_SLICE_X116Y118_A5Q),
.O5(CLBLM_L_X76Y118_SLICE_X116Y118_BO5),
.O6(CLBLM_L_X76Y118_SLICE_X116Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafafafffff0000)
  ) CLBLM_L_X76Y118_SLICE_X116Y118_ALUT (
.I0(CLBLM_L_X76Y123_SLICE_X117Y123_DO6),
.I1(1'b1),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(1'b1),
.I4(CLBLM_L_X76Y118_SLICE_X117Y118_AQ),
.I5(1'b1),
.O5(CLBLM_L_X76Y118_SLICE_X116Y118_AO5),
.O6(CLBLM_L_X76Y118_SLICE_X116Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y118_SLICE_X117Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y118_SLICE_X117Y118_AO6),
.Q(CLBLM_L_X76Y118_SLICE_X117Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y118_SLICE_X117Y118_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y118_SLICE_X117Y118_BO6),
.Q(CLBLM_L_X76Y118_SLICE_X117Y118_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y118_SLICE_X117Y118_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y118_SLICE_X117Y118_CO6),
.Q(CLBLM_L_X76Y118_SLICE_X117Y118_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y118_SLICE_X117Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y118_SLICE_X117Y118_DO5),
.O6(CLBLM_L_X76Y118_SLICE_X117Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeee4e4cecec4c4)
  ) CLBLM_L_X76Y118_SLICE_X117Y118_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X76Y118_SLICE_X116Y118_A5Q),
.I2(CLBLL_R_X77Y123_SLICE_X118Y123_DO6),
.I3(1'b1),
.I4(CLBLM_L_X76Y118_SLICE_X117Y118_CQ),
.I5(CLBLM_L_X76Y118_SLICE_X116Y118_BQ),
.O5(CLBLM_L_X76Y118_SLICE_X117Y118_CO5),
.O6(CLBLM_L_X76Y118_SLICE_X117Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafefefa0a0e0e0)
  ) CLBLM_L_X76Y118_SLICE_X117Y118_BLUT (
.I0(CLBLM_L_X76Y123_SLICE_X117Y123_DO6),
.I1(CLBLM_L_X76Y118_SLICE_X117Y118_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(1'b1),
.I4(CLBLM_L_X74Y123_SLICE_X113Y123_CO5),
.I5(CLBLM_L_X76Y118_SLICE_X116Y118_CQ),
.O5(CLBLM_L_X76Y118_SLICE_X117Y118_BO5),
.O6(CLBLM_L_X76Y118_SLICE_X117Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafacccc5050cccc)
  ) CLBLM_L_X76Y118_SLICE_X117Y118_ALUT (
.I0(CLBLM_L_X76Y123_SLICE_X117Y123_DO6),
.I1(CLBLM_L_X76Y118_SLICE_X117Y118_BQ),
.I2(CLBLM_L_X76Y118_SLICE_X117Y118_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X76Y118_SLICE_X116Y118_CQ),
.O5(CLBLM_L_X76Y118_SLICE_X117Y118_AO5),
.O6(CLBLM_L_X76Y118_SLICE_X117Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y119_SLICE_X116Y119_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y119_SLICE_X116Y119_AO5),
.Q(CLBLM_L_X76Y119_SLICE_X116Y119_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y119_SLICE_X116Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y119_SLICE_X116Y119_AO6),
.Q(CLBLM_L_X76Y119_SLICE_X116Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y119_SLICE_X116Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y119_SLICE_X116Y119_DO5),
.O6(CLBLM_L_X76Y119_SLICE_X116Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y119_SLICE_X116Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y119_SLICE_X116Y119_CO5),
.O6(CLBLM_L_X76Y119_SLICE_X116Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hddeeddeeddeeddee)
  ) CLBLM_L_X76Y119_SLICE_X116Y119_BLUT (
.I0(CLBLM_L_X76Y118_SLICE_X116Y118_AQ),
.I1(CLBLM_L_X76Y118_SLICE_X116Y118_BO6),
.I2(1'b1),
.I3(CLBLM_L_X76Y118_SLICE_X116Y118_DQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y119_SLICE_X116Y119_BO5),
.O6(CLBLM_L_X76Y119_SLICE_X116Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcfcfcf050a000)
  ) CLBLM_L_X76Y119_SLICE_X116Y119_ALUT (
.I0(CLBLM_L_X76Y123_SLICE_X117Y123_DO6),
.I1(CLBLM_L_X74Y117_SLICE_X112Y117_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLL_R_X77Y127_SLICE_X118Y127_AQ),
.I4(CLBLM_L_X76Y119_SLICE_X116Y119_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X76Y119_SLICE_X116Y119_AO5),
.O6(CLBLM_L_X76Y119_SLICE_X116Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y119_SLICE_X117Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y119_SLICE_X117Y119_DO5),
.O6(CLBLM_L_X76Y119_SLICE_X117Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y119_SLICE_X117Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y119_SLICE_X117Y119_CO5),
.O6(CLBLM_L_X76Y119_SLICE_X117Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y119_SLICE_X117Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y119_SLICE_X117Y119_BO5),
.O6(CLBLM_L_X76Y119_SLICE_X117Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y119_SLICE_X117Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y119_SLICE_X117Y119_AO5),
.O6(CLBLM_L_X76Y119_SLICE_X117Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y122_SLICE_X116Y122_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y122_SLICE_X116Y122_AO5),
.Q(CLBLM_L_X76Y122_SLICE_X116Y122_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y122_SLICE_X116Y122_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y122_SLICE_X116Y122_CO5),
.Q(CLBLM_L_X76Y122_SLICE_X116Y122_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y122_SLICE_X116Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y122_SLICE_X116Y122_AO6),
.Q(CLBLM_L_X76Y122_SLICE_X116Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y122_SLICE_X116Y122_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y122_SLICE_X116Y122_BO6),
.Q(CLBLM_L_X76Y122_SLICE_X116Y122_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y122_SLICE_X116Y122_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y122_SLICE_X116Y122_CO6),
.Q(CLBLM_L_X76Y122_SLICE_X116Y122_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y122_SLICE_X116Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y122_SLICE_X116Y122_DO5),
.O6(CLBLM_L_X76Y122_SLICE_X116Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0fff0e0e02020)
  ) CLBLM_L_X76Y122_SLICE_X116Y122_CLUT (
.I0(CLBLM_L_X76Y122_SLICE_X116Y122_C5Q),
.I1(CLBLM_L_X74Y123_SLICE_X113Y123_CO5),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X76Y125_SLICE_X116Y125_C5Q),
.I4(CLBLL_R_X77Y127_SLICE_X118Y127_AQ),
.I5(1'b1),
.O5(CLBLM_L_X76Y122_SLICE_X116Y122_CO5),
.O6(CLBLM_L_X76Y122_SLICE_X116Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaff00ccccff00)
  ) CLBLM_L_X76Y122_SLICE_X116Y122_BLUT (
.I0(CLBLL_R_X77Y127_SLICE_X118Y127_AQ),
.I1(CLBLM_L_X76Y122_SLICE_X116Y122_BQ),
.I2(1'b1),
.I3(CLBLM_L_X76Y124_SLICE_X116Y124_BQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X75Y123_SLICE_X114Y123_AO6),
.O5(CLBLM_L_X76Y122_SLICE_X116Y122_BO5),
.O6(CLBLM_L_X76Y122_SLICE_X116Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff500a0cceecc44)
  ) CLBLM_L_X76Y122_SLICE_X116Y122_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X76Y122_SLICE_X116Y122_BQ),
.I2(CLBLM_L_X76Y122_SLICE_X116Y122_AQ),
.I3(CLBLL_R_X75Y123_SLICE_X114Y123_AO6),
.I4(CLBLM_L_X76Y122_SLICE_X116Y122_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X76Y122_SLICE_X116Y122_AO5),
.O6(CLBLM_L_X76Y122_SLICE_X116Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y122_SLICE_X117Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y113_SLICE_X118Y113_AQ),
.Q(CLBLM_L_X76Y122_SLICE_X117Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y122_SLICE_X117Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y122_SLICE_X117Y122_DO5),
.O6(CLBLM_L_X76Y122_SLICE_X117Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y122_SLICE_X117Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y122_SLICE_X117Y122_CO5),
.O6(CLBLM_L_X76Y122_SLICE_X117Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y122_SLICE_X117Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y122_SLICE_X117Y122_BO5),
.O6(CLBLM_L_X76Y122_SLICE_X117Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y122_SLICE_X117Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y122_SLICE_X117Y122_AO5),
.O6(CLBLM_L_X76Y122_SLICE_X117Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y123_SLICE_X116Y123_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y123_SLICE_X115Y123_AO6),
.Q(CLBLM_L_X76Y123_SLICE_X116Y123_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y123_SLICE_X116Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y123_SLICE_X116Y123_AO6),
.Q(CLBLM_L_X76Y123_SLICE_X116Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y123_SLICE_X116Y123_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y123_SLICE_X116Y123_BO6),
.Q(CLBLM_L_X76Y123_SLICE_X116Y123_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y123_SLICE_X116Y123_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y123_SLICE_X116Y123_CO6),
.Q(CLBLM_L_X76Y123_SLICE_X116Y123_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h80ff80ff00ff00ff)
  ) CLBLM_L_X76Y123_SLICE_X116Y123_DLUT (
.I0(CLBLM_L_X76Y123_SLICE_X117Y123_AQ),
.I1(CLBLM_L_X74Y123_SLICE_X113Y123_A5Q),
.I2(CLBLL_R_X75Y113_SLICE_X114Y113_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(1'b1),
.I5(CLBLM_L_X74Y123_SLICE_X113Y123_BQ),
.O5(CLBLM_L_X76Y123_SLICE_X116Y123_DO5),
.O6(CLBLM_L_X76Y123_SLICE_X116Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6f006f00cf00cf00)
  ) CLBLM_L_X76Y123_SLICE_X116Y123_CLUT (
.I0(CLBLM_L_X74Y123_SLICE_X113Y123_CO5),
.I1(CLBLM_L_X76Y123_SLICE_X116Y123_CQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLL_R_X75Y121_SLICE_X114Y121_BQ),
.I4(1'b1),
.I5(CLBLL_R_X75Y123_SLICE_X115Y123_AQ),
.O5(CLBLM_L_X76Y123_SLICE_X116Y123_CO5),
.O6(CLBLM_L_X76Y123_SLICE_X116Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6acacaca0a0a0a0a)
  ) CLBLM_L_X76Y123_SLICE_X116Y123_BLUT (
.I0(CLBLM_L_X76Y123_SLICE_X116Y123_CQ),
.I1(CLBLM_L_X76Y123_SLICE_X116Y123_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLL_R_X75Y123_SLICE_X115Y123_AQ),
.I4(CLBLM_L_X74Y123_SLICE_X113Y123_CO5),
.I5(CLBLL_R_X75Y121_SLICE_X114Y121_BQ),
.O5(CLBLM_L_X76Y123_SLICE_X116Y123_BO5),
.O6(CLBLM_L_X76Y123_SLICE_X116Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0c0c00000000000)
  ) CLBLM_L_X76Y123_SLICE_X116Y123_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X76Y122_SLICE_X116Y122_A5Q),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X76Y122_SLICE_X116Y122_AQ),
.I4(CLBLM_L_X76Y122_SLICE_X116Y122_BQ),
.I5(CLBLL_R_X75Y123_SLICE_X115Y123_DO6),
.O5(CLBLM_L_X76Y123_SLICE_X116Y123_AO5),
.O6(CLBLM_L_X76Y123_SLICE_X116Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y123_SLICE_X117Y123_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y123_SLICE_X117Y123_BO5),
.Q(CLBLM_L_X76Y123_SLICE_X117Y123_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y123_SLICE_X117Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y123_SLICE_X117Y123_AO6),
.Q(CLBLM_L_X76Y123_SLICE_X117Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y123_SLICE_X117Y123_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y123_SLICE_X117Y123_BO6),
.Q(CLBLM_L_X76Y123_SLICE_X117Y123_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y123_SLICE_X117Y123_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y123_SLICE_X117Y123_CO6),
.Q(CLBLM_L_X76Y123_SLICE_X117Y123_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3030303a00000000)
  ) CLBLM_L_X76Y123_SLICE_X117Y123_DLUT (
.I0(CLBLM_L_X76Y122_SLICE_X116Y122_C5Q),
.I1(CLBLL_R_X77Y123_SLICE_X119Y123_BO6),
.I2(CLBLM_L_X76Y125_SLICE_X117Y125_BQ),
.I3(CLBLM_L_X76Y124_SLICE_X116Y124_CQ),
.I4(CLBLM_L_X76Y124_SLICE_X117Y124_AQ),
.I5(CLBLL_R_X75Y123_SLICE_X114Y123_AO6),
.O5(CLBLM_L_X76Y123_SLICE_X117Y123_DO5),
.O6(CLBLM_L_X76Y123_SLICE_X117Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdf558a00dfdf8a8a)
  ) CLBLM_L_X76Y123_SLICE_X117Y123_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X76Y123_SLICE_X117Y123_CQ),
.I2(CLBLM_L_X76Y125_SLICE_X117Y125_BQ),
.I3(CLBLM_L_X76Y122_SLICE_X117Y122_AQ),
.I4(CLBLM_L_X76Y123_SLICE_X117Y123_B5Q),
.I5(CLBLL_R_X77Y113_SLICE_X118Y113_AQ),
.O5(CLBLM_L_X76Y123_SLICE_X117Y123_CO5),
.O6(CLBLM_L_X76Y123_SLICE_X117Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0c0c0acfcacfc)
  ) CLBLM_L_X76Y123_SLICE_X117Y123_BLUT (
.I0(CLBLM_L_X76Y123_SLICE_X117Y123_B5Q),
.I1(CLBLM_L_X76Y123_SLICE_X117Y123_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X76Y125_SLICE_X117Y125_BQ),
.I4(CLBLM_L_X76Y130_SLICE_X116Y130_DQ),
.I5(1'b1),
.O5(CLBLM_L_X76Y123_SLICE_X117Y123_BO5),
.O6(CLBLM_L_X76Y123_SLICE_X117Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5af0ff00ff5f0000)
  ) CLBLM_L_X76Y123_SLICE_X117Y123_ALUT (
.I0(CLBLL_R_X75Y113_SLICE_X114Y113_AQ),
.I1(1'b1),
.I2(CLBLM_L_X76Y123_SLICE_X117Y123_AQ),
.I3(CLBLM_L_X74Y123_SLICE_X113Y123_A5Q),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLM_L_X76Y123_SLICE_X117Y123_AO5),
.O6(CLBLM_L_X76Y123_SLICE_X117Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y124_SLICE_X116Y124_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y123_SLICE_X116Y123_DO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y124_SLICE_X116Y124_B5Q),
.Q(CLBLM_L_X76Y124_SLICE_X116Y124_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y124_SLICE_X116Y124_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y123_SLICE_X116Y123_DO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y124_SLICE_X115Y124_DQ),
.Q(CLBLM_L_X76Y124_SLICE_X116Y124_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y124_SLICE_X116Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y123_SLICE_X116Y123_DO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y124_SLICE_X116Y124_AO5),
.Q(CLBLM_L_X76Y124_SLICE_X116Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y124_SLICE_X116Y124_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y123_SLICE_X116Y123_DO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y124_SLICE_X116Y124_BO5),
.Q(CLBLM_L_X76Y124_SLICE_X116Y124_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y124_SLICE_X116Y124_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y123_SLICE_X116Y123_DO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y124_SLICE_X117Y124_AQ),
.Q(CLBLM_L_X76Y124_SLICE_X116Y124_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y124_SLICE_X116Y124_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y123_SLICE_X116Y123_DO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X75Y124_SLICE_X115Y124_CQ),
.Q(CLBLM_L_X76Y124_SLICE_X116Y124_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y124_SLICE_X116Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y124_SLICE_X116Y124_DO5),
.O6(CLBLM_L_X76Y124_SLICE_X116Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc8ffc4ff32ff31)
  ) CLBLM_L_X76Y124_SLICE_X116Y124_CLUT (
.I0(CLBLM_L_X76Y124_SLICE_X116Y124_AO6),
.I1(CLBLM_L_X76Y122_SLICE_X116Y122_C5Q),
.I2(CLBLM_L_X76Y124_SLICE_X117Y124_DO6),
.I3(CLBLL_R_X75Y123_SLICE_X115Y123_AO5),
.I4(CLBLM_L_X76Y122_SLICE_X116Y122_BQ),
.I5(CLBLM_L_X76Y124_SLICE_X116Y124_BO6),
.O5(CLBLM_L_X76Y124_SLICE_X116Y124_CO5),
.O6(CLBLM_L_X76Y124_SLICE_X116Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1d441d77ff00ff00)
  ) CLBLM_L_X76Y124_SLICE_X116Y124_BLUT (
.I0(CLBLM_L_X76Y124_SLICE_X116Y124_A5Q),
.I1(CLBLM_L_X76Y124_SLICE_X116Y124_BQ),
.I2(CLBLM_L_X76Y124_SLICE_X116Y124_AQ),
.I3(CLBLL_R_X75Y124_SLICE_X115Y124_AQ),
.I4(CLBLM_L_X76Y124_SLICE_X116Y124_CQ),
.I5(1'b1),
.O5(CLBLM_L_X76Y124_SLICE_X116Y124_BO5),
.O6(CLBLM_L_X76Y124_SLICE_X116Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000cccccccc)
  ) CLBLM_L_X76Y124_SLICE_X116Y124_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X76Y124_SLICE_X116Y124_DQ),
.I2(CLBLL_R_X75Y122_SLICE_X115Y122_A5Q),
.I3(CLBLL_R_X75Y124_SLICE_X115Y124_AQ),
.I4(CLBLM_L_X76Y122_SLICE_X116Y122_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X76Y124_SLICE_X116Y124_AO5),
.O6(CLBLM_L_X76Y124_SLICE_X116Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y124_SLICE_X117Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y124_SLICE_X117Y124_AO6),
.Q(CLBLM_L_X76Y124_SLICE_X117Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y124_SLICE_X117Y124_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y124_SLICE_X117Y124_BO6),
.Q(CLBLM_L_X76Y124_SLICE_X117Y124_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff0ffffffcc)
  ) CLBLM_L_X76Y124_SLICE_X117Y124_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X76Y124_SLICE_X117Y124_AQ),
.I2(CLBLM_L_X76Y124_SLICE_X116Y124_B5Q),
.I3(CLBLM_L_X76Y125_SLICE_X117Y125_BQ),
.I4(CLBLM_L_X76Y122_SLICE_X116Y122_C5Q),
.I5(CLBLL_R_X75Y124_SLICE_X115Y124_AQ),
.O5(CLBLM_L_X76Y124_SLICE_X117Y124_DO5),
.O6(CLBLM_L_X76Y124_SLICE_X117Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00df00ff00df)
  ) CLBLM_L_X76Y124_SLICE_X117Y124_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X76Y119_SLICE_X116Y119_BO6),
.I2(CLBLL_R_X75Y122_SLICE_X114Y122_AQ),
.I3(CLBLM_L_X76Y123_SLICE_X117Y123_AO5),
.I4(CLBLM_L_X76Y125_SLICE_X117Y125_BQ),
.I5(1'b1),
.O5(CLBLM_L_X76Y124_SLICE_X117Y124_CO5),
.O6(CLBLM_L_X76Y124_SLICE_X117Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaccaaacaaccaa)
  ) CLBLM_L_X76Y124_SLICE_X117Y124_BLUT (
.I0(CLBLL_R_X77Y123_SLICE_X119Y123_CQ),
.I1(CLBLM_L_X76Y124_SLICE_X117Y124_BQ),
.I2(CLBLL_R_X75Y113_SLICE_X114Y113_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X76Y123_SLICE_X117Y123_AQ),
.I5(CLBLM_L_X74Y123_SLICE_X113Y123_A5Q),
.O5(CLBLM_L_X76Y124_SLICE_X117Y124_BO5),
.O6(CLBLM_L_X76Y124_SLICE_X117Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacafa0acacafa0a)
  ) CLBLM_L_X76Y124_SLICE_X117Y124_ALUT (
.I0(CLBLM_L_X76Y122_SLICE_X116Y122_C5Q),
.I1(CLBLM_L_X76Y124_SLICE_X116Y124_BO6),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X76Y124_SLICE_X117Y124_AQ),
.I4(CLBLM_L_X74Y123_SLICE_X113Y123_CO5),
.I5(1'b1),
.O5(CLBLM_L_X76Y124_SLICE_X117Y124_AO5),
.O6(CLBLM_L_X76Y124_SLICE_X117Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y125_SLICE_X116Y125_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y125_SLICE_X116Y125_AO5),
.Q(CLBLM_L_X76Y125_SLICE_X116Y125_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y125_SLICE_X116Y125_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y125_SLICE_X116Y125_CO5),
.Q(CLBLM_L_X76Y125_SLICE_X116Y125_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y125_SLICE_X116Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y125_SLICE_X116Y125_AO6),
.Q(CLBLM_L_X76Y125_SLICE_X116Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y125_SLICE_X116Y125_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y125_SLICE_X116Y125_BO6),
.Q(CLBLM_L_X76Y125_SLICE_X116Y125_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y125_SLICE_X116Y125_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y125_SLICE_X116Y125_CO6),
.Q(CLBLM_L_X76Y125_SLICE_X116Y125_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y125_SLICE_X116Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y125_SLICE_X116Y125_DO5),
.O6(CLBLM_L_X76Y125_SLICE_X116Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f0f33000a0a0a0a)
  ) CLBLM_L_X76Y125_SLICE_X116Y125_CLUT (
.I0(CLBLM_R_X65Y105_SLICE_X99Y105_CQ),
.I1(CLBLM_L_X76Y125_SLICE_X116Y125_CQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLL_R_X77Y127_SLICE_X119Y127_AO5),
.I4(CLBLL_R_X77Y127_SLICE_X119Y127_AQ),
.I5(1'b1),
.O5(CLBLM_L_X76Y125_SLICE_X116Y125_CO5),
.O6(CLBLM_L_X76Y125_SLICE_X116Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hba30ba3030303030)
  ) CLBLM_L_X76Y125_SLICE_X116Y125_BLUT (
.I0(CLBLM_L_X76Y126_SLICE_X116Y126_AO6),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_L_X74Y123_SLICE_X112Y123_BQ),
.I3(CLBLM_L_X76Y126_SLICE_X117Y126_AQ),
.I4(1'b1),
.I5(CLBLL_R_X77Y127_SLICE_X119Y127_AO5),
.O5(CLBLM_L_X76Y125_SLICE_X116Y125_BO5),
.O6(CLBLM_L_X76Y125_SLICE_X116Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbb8888fc30fc30)
  ) CLBLM_L_X76Y125_SLICE_X116Y125_ALUT (
.I0(CLBLL_R_X79Y127_SLICE_X122Y127_BQ),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_L_X76Y125_SLICE_X116Y125_AQ),
.I3(CLBLL_R_X79Y127_SLICE_X122Y127_CQ),
.I4(CLBLM_L_X76Y123_SLICE_X116Y123_AQ),
.I5(1'b1),
.O5(CLBLM_L_X76Y125_SLICE_X116Y125_AO5),
.O6(CLBLM_L_X76Y125_SLICE_X116Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y125_SLICE_X117Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y125_SLICE_X117Y125_AO6),
.Q(CLBLM_L_X76Y125_SLICE_X117Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y125_SLICE_X117Y125_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y125_SLICE_X117Y125_BO6),
.Q(CLBLM_L_X76Y125_SLICE_X117Y125_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7555200075552000)
  ) CLBLM_L_X76Y125_SLICE_X117Y125_DLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X77Y124_SLICE_X119Y124_CQ),
.I2(CLBLL_R_X75Y122_SLICE_X114Y122_AQ),
.I3(CLBLM_L_X76Y125_SLICE_X117Y125_BQ),
.I4(CLBLM_L_X76Y118_SLICE_X117Y118_CQ),
.I5(1'b1),
.O5(CLBLM_L_X76Y125_SLICE_X117Y125_DO5),
.O6(CLBLM_L_X76Y125_SLICE_X117Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff57575757575757)
  ) CLBLM_L_X76Y125_SLICE_X117Y125_CLUT (
.I0(CLBLL_R_X77Y125_SLICE_X118Y125_BQ),
.I1(CLBLM_L_X76Y124_SLICE_X116Y124_CO6),
.I2(CLBLL_R_X75Y122_SLICE_X114Y122_AQ),
.I3(CLBLM_L_X74Y123_SLICE_X113Y123_A5Q),
.I4(CLBLM_L_X76Y123_SLICE_X117Y123_AQ),
.I5(CLBLM_L_X74Y109_SLICE_X113Y109_AQ),
.O5(CLBLM_L_X76Y125_SLICE_X117Y125_CO5),
.O6(CLBLM_L_X76Y125_SLICE_X117Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaeeeeaaaafeee)
  ) CLBLM_L_X76Y125_SLICE_X117Y125_BLUT (
.I0(CLBLM_L_X76Y125_SLICE_X117Y125_DO6),
.I1(CLBLM_L_X76Y125_SLICE_X117Y125_BQ),
.I2(CLBLM_L_X76Y123_SLICE_X117Y123_AQ),
.I3(CLBLL_R_X75Y113_SLICE_X114Y113_AQ),
.I4(CLBLM_L_X76Y124_SLICE_X117Y124_CO6),
.I5(CLBLM_L_X74Y123_SLICE_X113Y123_A5Q),
.O5(CLBLM_L_X76Y125_SLICE_X117Y125_BO5),
.O6(CLBLM_L_X76Y125_SLICE_X117Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00a0cccc0fa0cccc)
  ) CLBLM_L_X76Y125_SLICE_X117Y125_ALUT (
.I0(CLBLL_R_X77Y123_SLICE_X119Y123_DO6),
.I1(CLBLM_L_X76Y126_SLICE_X117Y126_AQ),
.I2(CLBLM_L_X76Y125_SLICE_X117Y125_AQ),
.I3(CLBLL_R_X75Y123_SLICE_X115Y123_DO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X77Y122_SLICE_X118Y122_CO6),
.O5(CLBLM_L_X76Y125_SLICE_X117Y125_AO5),
.O6(CLBLM_L_X76Y125_SLICE_X117Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y126_SLICE_X116Y126_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y126_SLICE_X116Y126_BO5),
.Q(CLBLM_L_X76Y126_SLICE_X116Y126_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y126_SLICE_X116Y126_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y126_SLICE_X116Y126_BO6),
.Q(CLBLM_L_X76Y126_SLICE_X116Y126_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y126_SLICE_X116Y126_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y126_SLICE_X116Y126_CO6),
.Q(CLBLM_L_X76Y126_SLICE_X116Y126_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y126_SLICE_X116Y126_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y126_SLICE_X116Y126_DO6),
.Q(CLBLM_L_X76Y126_SLICE_X116Y126_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7cf4f4f444444444)
  ) CLBLM_L_X76Y126_SLICE_X116Y126_DLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X76Y126_SLICE_X116Y126_CQ),
.I2(CLBLM_L_X76Y126_SLICE_X116Y126_DQ),
.I3(CLBLM_L_X76Y126_SLICE_X116Y126_AO5),
.I4(CLBLM_L_X76Y126_SLICE_X116Y126_B5Q),
.I5(CLBLL_R_X77Y127_SLICE_X119Y127_AO5),
.O5(CLBLM_L_X76Y126_SLICE_X116Y126_DO5),
.O6(CLBLM_L_X76Y126_SLICE_X116Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f55ff00d5550000)
  ) CLBLM_L_X76Y126_SLICE_X116Y126_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X76Y125_SLICE_X116Y125_CQ),
.I2(CLBLM_L_X76Y126_SLICE_X116Y126_BQ),
.I3(CLBLL_R_X77Y127_SLICE_X119Y127_AO5),
.I4(CLBLM_L_X76Y126_SLICE_X116Y126_B5Q),
.I5(CLBLM_L_X76Y126_SLICE_X116Y126_CQ),
.O5(CLBLM_L_X76Y126_SLICE_X116Y126_CO5),
.O6(CLBLM_L_X76Y126_SLICE_X116Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c00fcf06a00eecc)
  ) CLBLM_L_X76Y126_SLICE_X116Y126_BLUT (
.I0(CLBLM_L_X76Y126_SLICE_X116Y126_B5Q),
.I1(CLBLM_L_X76Y126_SLICE_X116Y126_BQ),
.I2(CLBLM_L_X76Y125_SLICE_X116Y125_CQ),
.I3(CLBLL_R_X77Y127_SLICE_X119Y127_AO5),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLM_L_X76Y126_SLICE_X116Y126_BO5),
.O6(CLBLM_L_X76Y126_SLICE_X116Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000f0f00000)
  ) CLBLM_L_X76Y126_SLICE_X116Y126_ALUT (
.I0(CLBLM_L_X76Y126_SLICE_X116Y126_B5Q),
.I1(CLBLM_L_X76Y126_SLICE_X116Y126_DQ),
.I2(CLBLM_L_X76Y125_SLICE_X116Y125_CQ),
.I3(CLBLM_L_X76Y126_SLICE_X116Y126_CQ),
.I4(CLBLM_L_X76Y126_SLICE_X116Y126_BQ),
.I5(1'b1),
.O5(CLBLM_L_X76Y126_SLICE_X116Y126_AO5),
.O6(CLBLM_L_X76Y126_SLICE_X116Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y126_SLICE_X117Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y126_SLICE_X117Y126_AO6),
.Q(CLBLM_L_X76Y126_SLICE_X117Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y126_SLICE_X117Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y126_SLICE_X117Y126_DO5),
.O6(CLBLM_L_X76Y126_SLICE_X117Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y126_SLICE_X117Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y126_SLICE_X117Y126_CO5),
.O6(CLBLM_L_X76Y126_SLICE_X117Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y126_SLICE_X117Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y126_SLICE_X117Y126_BO5),
.O6(CLBLM_L_X76Y126_SLICE_X117Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0cae0caec0eac0ea)
  ) CLBLM_L_X76Y126_SLICE_X117Y126_ALUT (
.I0(CLBLM_L_X76Y126_SLICE_X116Y126_DQ),
.I1(CLBLL_R_X77Y127_SLICE_X119Y127_AO5),
.I2(CLBLM_L_X76Y126_SLICE_X117Y126_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(1'b1),
.I5(CLBLM_L_X76Y126_SLICE_X116Y126_AO6),
.O5(CLBLM_L_X76Y126_SLICE_X117Y126_AO5),
.O6(CLBLM_L_X76Y126_SLICE_X117Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y127_SLICE_X116Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y129_SLICE_X118Y129_AQ),
.Q(CLBLM_L_X76Y127_SLICE_X116Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y127_SLICE_X116Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y127_SLICE_X116Y127_DO5),
.O6(CLBLM_L_X76Y127_SLICE_X116Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y127_SLICE_X116Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y127_SLICE_X116Y127_CO5),
.O6(CLBLM_L_X76Y127_SLICE_X116Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y127_SLICE_X116Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y127_SLICE_X116Y127_BO5),
.O6(CLBLM_L_X76Y127_SLICE_X116Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y127_SLICE_X116Y127_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y127_SLICE_X116Y127_AO5),
.O6(CLBLM_L_X76Y127_SLICE_X116Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y127_SLICE_X117Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y127_SLICE_X117Y127_DO5),
.O6(CLBLM_L_X76Y127_SLICE_X117Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y127_SLICE_X117Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y127_SLICE_X117Y127_CO5),
.O6(CLBLM_L_X76Y127_SLICE_X117Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y127_SLICE_X117Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y127_SLICE_X117Y127_BO5),
.O6(CLBLM_L_X76Y127_SLICE_X117Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y127_SLICE_X117Y127_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y127_SLICE_X117Y127_AO5),
.O6(CLBLM_L_X76Y127_SLICE_X117Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y128_SLICE_X116Y128_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y128_SLICE_X116Y128_CQ),
.Q(CLBLM_L_X76Y128_SLICE_X116Y128_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y128_SLICE_X116Y128_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y128_SLICE_X116Y128_CO5),
.Q(CLBLM_L_X76Y128_SLICE_X116Y128_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y128_SLICE_X116Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y128_SLICE_X116Y128_AO6),
.Q(CLBLM_L_X76Y128_SLICE_X116Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y128_SLICE_X116Y128_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y128_SLICE_X116Y128_BO6),
.Q(CLBLM_L_X76Y128_SLICE_X116Y128_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y128_SLICE_X116Y128_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y128_SLICE_X116Y128_CO6),
.Q(CLBLM_L_X76Y128_SLICE_X116Y128_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000200000002)
  ) CLBLM_L_X76Y128_SLICE_X116Y128_DLUT (
.I0(CLBLL_R_X77Y128_SLICE_X118Y128_AQ),
.I1(CLBLL_R_X77Y126_SLICE_X118Y126_BQ),
.I2(CLBLM_L_X76Y128_SLICE_X116Y128_AQ),
.I3(CLBLM_L_X76Y128_SLICE_X116Y128_BQ),
.I4(CLBLM_L_X76Y128_SLICE_X117Y128_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X76Y128_SLICE_X116Y128_DO5),
.O6(CLBLM_L_X76Y128_SLICE_X116Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaacc0fff0f00)
  ) CLBLM_L_X76Y128_SLICE_X116Y128_CLUT (
.I0(CLBLM_L_X76Y125_SLICE_X116Y125_A5Q),
.I1(CLBLM_L_X76Y128_SLICE_X116Y128_AQ),
.I2(CLBLM_L_X76Y129_SLICE_X116Y129_B5Q),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X76Y130_SLICE_X116Y130_DQ),
.I5(1'b1),
.O5(CLBLM_L_X76Y128_SLICE_X116Y128_CO5),
.O6(CLBLM_L_X76Y128_SLICE_X116Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h77aaffaa08aa00aa)
  ) CLBLM_L_X76Y128_SLICE_X116Y128_BLUT (
.I0(CLBLM_L_X76Y128_SLICE_X117Y128_A5Q),
.I1(CLBLL_R_X77Y126_SLICE_X118Y126_AQ),
.I2(CLBLM_L_X76Y128_SLICE_X116Y128_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLL_R_X77Y126_SLICE_X118Y126_BQ),
.I5(CLBLM_L_X76Y128_SLICE_X116Y128_BQ),
.O5(CLBLM_L_X76Y128_SLICE_X116Y128_BO5),
.O6(CLBLM_L_X76Y128_SLICE_X116Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h58f0f0f0cccccccc)
  ) CLBLM_L_X76Y128_SLICE_X116Y128_ALUT (
.I0(CLBLM_L_X76Y128_SLICE_X117Y128_A5Q),
.I1(CLBLM_L_X76Y128_SLICE_X116Y128_BQ),
.I2(CLBLM_L_X76Y128_SLICE_X116Y128_AQ),
.I3(CLBLL_R_X77Y126_SLICE_X118Y126_AQ),
.I4(CLBLL_R_X77Y126_SLICE_X118Y126_BQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X76Y128_SLICE_X116Y128_AO5),
.O6(CLBLM_L_X76Y128_SLICE_X116Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y128_SLICE_X117Y128_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y128_SLICE_X117Y128_CO5),
.Q(CLBLM_L_X76Y128_SLICE_X117Y128_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y128_SLICE_X117Y128_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y128_SLICE_X117Y128_BO5),
.Q(CLBLM_L_X76Y128_SLICE_X117Y128_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y128_SLICE_X117Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y128_SLICE_X117Y128_AO6),
.Q(CLBLM_L_X76Y128_SLICE_X117Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y128_SLICE_X117Y128_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y128_SLICE_X117Y128_BO6),
.Q(CLBLM_L_X76Y128_SLICE_X117Y128_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y128_SLICE_X117Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y128_SLICE_X117Y128_DO5),
.O6(CLBLM_L_X76Y128_SLICE_X117Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha000000077bbcc00)
  ) CLBLM_L_X76Y128_SLICE_X117Y128_CLUT (
.I0(CLBLL_R_X77Y126_SLICE_X118Y126_AQ),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_L_X76Y128_SLICE_X116Y128_AQ),
.I3(CLBLM_L_X76Y128_SLICE_X117Y128_A5Q),
.I4(CLBLL_R_X77Y126_SLICE_X118Y126_BQ),
.I5(1'b1),
.O5(CLBLM_L_X76Y128_SLICE_X117Y128_CO5),
.O6(CLBLM_L_X76Y128_SLICE_X117Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000030c00c0c6cac)
  ) CLBLM_L_X76Y128_SLICE_X117Y128_BLUT (
.I0(CLBLM_L_X76Y128_SLICE_X117Y128_B5Q),
.I1(CLBLM_L_X76Y128_SLICE_X117Y128_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLL_R_X77Y128_SLICE_X118Y128_CO6),
.I4(CLBLL_R_X77Y128_SLICE_X118Y128_AQ),
.I5(1'b1),
.O5(CLBLM_L_X76Y128_SLICE_X117Y128_BO5),
.O6(CLBLM_L_X76Y128_SLICE_X117Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeff55ffaaaaaaaa)
  ) CLBLM_L_X76Y128_SLICE_X117Y128_ALUT (
.I0(CLBLM_L_X76Y128_SLICE_X117Y128_B5Q),
.I1(CLBLM_L_X76Y128_SLICE_X117Y128_BQ),
.I2(1'b1),
.I3(CLBLL_R_X77Y129_SLICE_X118Y129_AQ),
.I4(CLBLM_L_X76Y128_SLICE_X116Y128_CQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X76Y128_SLICE_X117Y128_AO5),
.O6(CLBLM_L_X76Y128_SLICE_X117Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y129_SLICE_X116Y129_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y128_SLICE_X116Y128_C5Q),
.Q(CLBLM_L_X76Y129_SLICE_X116Y129_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y129_SLICE_X116Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y129_SLICE_X116Y129_CQ),
.Q(CLBLM_L_X76Y129_SLICE_X116Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y129_SLICE_X116Y129_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y129_SLICE_X116Y129_BO6),
.Q(CLBLM_L_X76Y129_SLICE_X116Y129_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y129_SLICE_X116Y129_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y129_SLICE_X116Y129_CO6),
.Q(CLBLM_L_X76Y129_SLICE_X116Y129_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffff0000fffd)
  ) CLBLM_L_X76Y129_SLICE_X116Y129_DLUT (
.I0(CLBLM_L_X76Y127_SLICE_X116Y127_AQ),
.I1(CLBLM_L_X76Y130_SLICE_X116Y130_BQ),
.I2(CLBLL_R_X77Y129_SLICE_X118Y129_CQ),
.I3(CLBLM_L_X76Y130_SLICE_X116Y130_A5Q),
.I4(CLBLM_L_X76Y129_SLICE_X116Y129_BQ),
.I5(CLBLL_R_X77Y128_SLICE_X118Y128_CQ),
.O5(CLBLM_L_X76Y129_SLICE_X116Y129_DO5),
.O6(CLBLM_L_X76Y129_SLICE_X116Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5fdddddd0a888888)
  ) CLBLM_L_X76Y129_SLICE_X116Y129_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X76Y129_SLICE_X116Y129_CQ),
.I2(CLBLM_L_X76Y129_SLICE_X116Y129_AQ),
.I3(CLBLM_L_X76Y128_SLICE_X116Y128_C5Q),
.I4(CLBLM_L_X76Y129_SLICE_X116Y129_B5Q),
.I5(CLBLM_L_X76Y125_SLICE_X116Y125_BQ),
.O5(CLBLM_L_X76Y129_SLICE_X116Y129_CO5),
.O6(CLBLM_L_X76Y129_SLICE_X116Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h337f004c33f700c4)
  ) CLBLM_L_X76Y129_SLICE_X116Y129_BLUT (
.I0(CLBLL_R_X75Y130_SLICE_X115Y130_BO5),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_L_X76Y130_SLICE_X116Y130_AQ),
.I3(CLBLM_L_X76Y129_SLICE_X116Y129_DO6),
.I4(CLBLL_R_X75Y129_SLICE_X114Y129_BQ),
.I5(CLBLM_L_X76Y129_SLICE_X116Y129_AO5),
.O5(CLBLM_L_X76Y129_SLICE_X116Y129_BO5),
.O6(CLBLM_L_X76Y129_SLICE_X116Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafbf504050405040)
  ) CLBLM_L_X76Y129_SLICE_X116Y129_ALUT (
.I0(CLBLM_L_X76Y128_SLICE_X117Y128_AQ),
.I1(CLBLM_L_X78Y131_SLICE_X120Y131_AQ),
.I2(CLBLL_R_X77Y129_SLICE_X119Y129_BQ),
.I3(CLBLL_R_X77Y130_SLICE_X118Y130_AQ),
.I4(CLBLL_R_X75Y129_SLICE_X114Y129_BQ),
.I5(1'b1),
.O5(CLBLM_L_X76Y129_SLICE_X116Y129_AO5),
.O6(CLBLM_L_X76Y129_SLICE_X116Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y129_SLICE_X117Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y129_SLICE_X117Y129_DO5),
.O6(CLBLM_L_X76Y129_SLICE_X117Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y129_SLICE_X117Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y129_SLICE_X117Y129_CO5),
.O6(CLBLM_L_X76Y129_SLICE_X117Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y129_SLICE_X117Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y129_SLICE_X117Y129_BO5),
.O6(CLBLM_L_X76Y129_SLICE_X117Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y129_SLICE_X117Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y129_SLICE_X117Y129_AO5),
.O6(CLBLM_L_X76Y129_SLICE_X117Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y130_SLICE_X116Y130_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y130_SLICE_X116Y130_CO5),
.Q(CLBLM_L_X76Y130_SLICE_X116Y130_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y130_SLICE_X116Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y130_SLICE_X116Y130_AO6),
.Q(CLBLM_L_X76Y130_SLICE_X116Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y130_SLICE_X116Y130_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y130_SLICE_X116Y130_BO6),
.Q(CLBLM_L_X76Y130_SLICE_X116Y130_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y130_SLICE_X116Y130_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y130_SLICE_X116Y130_DO6),
.Q(CLBLM_L_X76Y130_SLICE_X116Y130_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h72fff0ffd800f000)
  ) CLBLM_L_X76Y130_SLICE_X116Y130_DLUT (
.I0(CLBLM_L_X76Y128_SLICE_X116Y128_C5Q),
.I1(CLBLM_L_X76Y129_SLICE_X116Y129_CQ),
.I2(CLBLM_L_X76Y130_SLICE_X116Y130_DQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X76Y129_SLICE_X116Y129_B5Q),
.I5(CLBLM_L_X76Y129_SLICE_X116Y129_AQ),
.O5(CLBLM_L_X76Y130_SLICE_X116Y130_DO5),
.O6(CLBLM_L_X76Y130_SLICE_X116Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000f000f7f0a0000)
  ) CLBLM_L_X76Y130_SLICE_X116Y130_CLUT (
.I0(CLBLL_R_X75Y130_SLICE_X115Y130_BO5),
.I1(CLBLL_R_X75Y130_SLICE_X114Y130_AQ),
.I2(CLBLM_L_X76Y130_SLICE_X116Y130_BQ),
.I3(CLBLM_L_X76Y130_SLICE_X116Y130_A5Q),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLM_L_X76Y130_SLICE_X116Y130_CO5),
.O6(CLBLM_L_X76Y130_SLICE_X116Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeaeeee222a2222)
  ) CLBLM_L_X76Y130_SLICE_X116Y130_BLUT (
.I0(CLBLL_R_X75Y130_SLICE_X114Y130_AQ),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLL_R_X77Y128_SLICE_X118Y128_CQ),
.I3(CLBLL_R_X77Y129_SLICE_X118Y129_CQ),
.I4(CLBLM_L_X76Y127_SLICE_X116Y127_AQ),
.I5(CLBLM_L_X76Y130_SLICE_X116Y130_BQ),
.O5(CLBLM_L_X76Y130_SLICE_X116Y130_BO5),
.O6(CLBLM_L_X76Y130_SLICE_X116Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb4fff000f0fff000)
  ) CLBLM_L_X76Y130_SLICE_X116Y130_ALUT (
.I0(CLBLL_R_X75Y130_SLICE_X114Y130_AQ),
.I1(CLBLM_L_X76Y130_SLICE_X116Y130_BQ),
.I2(CLBLM_L_X76Y130_SLICE_X116Y130_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X76Y129_SLICE_X116Y129_BQ),
.I5(CLBLL_R_X75Y130_SLICE_X115Y130_BO5),
.O5(CLBLM_L_X76Y130_SLICE_X116Y130_AO5),
.O6(CLBLM_L_X76Y130_SLICE_X116Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y130_SLICE_X117Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y130_SLICE_X117Y130_DO5),
.O6(CLBLM_L_X76Y130_SLICE_X117Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y130_SLICE_X117Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y130_SLICE_X117Y130_CO5),
.O6(CLBLM_L_X76Y130_SLICE_X117Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y130_SLICE_X117Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y130_SLICE_X117Y130_BO5),
.O6(CLBLM_L_X76Y130_SLICE_X117Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y130_SLICE_X117Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y130_SLICE_X117Y130_AO5),
.O6(CLBLM_L_X76Y130_SLICE_X117Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y133_SLICE_X116Y133_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y133_SLICE_X116Y133_AO6),
.Q(CLBLM_L_X76Y133_SLICE_X116Y133_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y133_SLICE_X116Y133_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y133_SLICE_X116Y133_BO6),
.Q(CLBLM_L_X76Y133_SLICE_X116Y133_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y133_SLICE_X116Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y133_SLICE_X116Y133_DO5),
.O6(CLBLM_L_X76Y133_SLICE_X116Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y133_SLICE_X116Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y133_SLICE_X116Y133_CO5),
.O6(CLBLM_L_X76Y133_SLICE_X116Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd0d050c05050d0c0)
  ) CLBLM_L_X76Y133_SLICE_X116Y133_BLUT (
.I0(CLBLM_L_X76Y134_SLICE_X116Y134_DO6),
.I1(CLBLM_L_X76Y133_SLICE_X116Y133_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLL_R_X75Y134_SLICE_X115Y134_AQ),
.I4(CLBLL_R_X75Y133_SLICE_X115Y133_BQ),
.I5(CLBLM_L_X74Y132_SLICE_X112Y132_C5Q),
.O5(CLBLM_L_X76Y133_SLICE_X116Y133_BO5),
.O6(CLBLM_L_X76Y133_SLICE_X116Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f337b730c004840)
  ) CLBLM_L_X76Y133_SLICE_X116Y133_ALUT (
.I0(CLBLL_R_X75Y134_SLICE_X115Y134_AQ),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_L_X76Y133_SLICE_X116Y133_AQ),
.I3(CLBLM_L_X76Y134_SLICE_X117Y134_CO6),
.I4(CLBLL_R_X75Y133_SLICE_X115Y133_BQ),
.I5(CLBLL_R_X75Y133_SLICE_X115Y133_AQ),
.O5(CLBLM_L_X76Y133_SLICE_X116Y133_AO5),
.O6(CLBLM_L_X76Y133_SLICE_X116Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y133_SLICE_X117Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y133_SLICE_X117Y133_DO5),
.O6(CLBLM_L_X76Y133_SLICE_X117Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y133_SLICE_X117Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y133_SLICE_X117Y133_CO5),
.O6(CLBLM_L_X76Y133_SLICE_X117Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y133_SLICE_X117Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y133_SLICE_X117Y133_BO5),
.O6(CLBLM_L_X76Y133_SLICE_X117Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y133_SLICE_X117Y133_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y133_SLICE_X117Y133_AO5),
.O6(CLBLM_L_X76Y133_SLICE_X117Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y134_SLICE_X116Y134_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y134_SLICE_X116Y134_AO6),
.Q(CLBLM_L_X76Y134_SLICE_X116Y134_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y134_SLICE_X116Y134_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y134_SLICE_X116Y134_BO6),
.Q(CLBLM_L_X76Y134_SLICE_X116Y134_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfffdf005fff5f00)
  ) CLBLM_L_X76Y134_SLICE_X116Y134_DLUT (
.I0(CLBLM_L_X76Y134_SLICE_X117Y134_AQ),
.I1(CLBLL_R_X75Y134_SLICE_X114Y134_A5Q),
.I2(CLBLM_L_X76Y134_SLICE_X116Y134_AQ),
.I3(CLBLL_R_X75Y133_SLICE_X115Y133_AQ),
.I4(CLBLL_R_X75Y134_SLICE_X115Y134_AO5),
.I5(CLBLL_R_X75Y134_SLICE_X115Y134_AO6),
.O5(CLBLM_L_X76Y134_SLICE_X116Y134_DO5),
.O6(CLBLM_L_X76Y134_SLICE_X116Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4c4ccccc4cffccff)
  ) CLBLM_L_X76Y134_SLICE_X116Y134_CLUT (
.I0(CLBLM_L_X76Y133_SLICE_X116Y133_AQ),
.I1(CLBLM_L_X76Y134_SLICE_X117Y134_CO6),
.I2(CLBLM_L_X76Y134_SLICE_X116Y134_BQ),
.I3(CLBLL_R_X75Y134_SLICE_X115Y134_AQ),
.I4(CLBLM_L_X76Y134_SLICE_X116Y134_AQ),
.I5(CLBLL_R_X75Y133_SLICE_X115Y133_BQ),
.O5(CLBLM_L_X76Y134_SLICE_X116Y134_CO5),
.O6(CLBLM_L_X76Y134_SLICE_X116Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaa60aaccaac0aa)
  ) CLBLM_L_X76Y134_SLICE_X116Y134_BLUT (
.I0(CLBLM_L_X76Y134_SLICE_X116Y134_AQ),
.I1(CLBLM_L_X76Y134_SLICE_X116Y134_BQ),
.I2(CLBLM_L_X76Y134_SLICE_X117Y134_CO6),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLL_R_X75Y134_SLICE_X115Y134_DO5),
.I5(CLBLM_L_X76Y133_SLICE_X116Y133_AQ),
.O5(CLBLM_L_X76Y134_SLICE_X116Y134_BO5),
.O6(CLBLM_L_X76Y134_SLICE_X116Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h50ffa00062ffa200)
  ) CLBLM_L_X76Y134_SLICE_X116Y134_ALUT (
.I0(CLBLM_L_X76Y134_SLICE_X116Y134_AQ),
.I1(CLBLL_R_X75Y133_SLICE_X115Y133_BQ),
.I2(CLBLM_L_X76Y134_SLICE_X117Y134_CO6),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X76Y133_SLICE_X116Y133_AQ),
.I5(CLBLL_R_X75Y134_SLICE_X115Y134_AQ),
.O5(CLBLM_L_X76Y134_SLICE_X116Y134_AO5),
.O6(CLBLM_L_X76Y134_SLICE_X116Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y134_SLICE_X117Y134_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y134_SLICE_X117Y134_AO6),
.Q(CLBLM_L_X76Y134_SLICE_X117Y134_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X76Y134_SLICE_X117Y134_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y134_SLICE_X117Y134_BO6),
.Q(CLBLM_L_X76Y134_SLICE_X117Y134_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y134_SLICE_X117Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y134_SLICE_X117Y134_DO5),
.O6(CLBLM_L_X76Y134_SLICE_X117Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0047007700330033)
  ) CLBLM_L_X76Y134_SLICE_X117Y134_CLUT (
.I0(CLBLL_R_X75Y134_SLICE_X114Y134_A5Q),
.I1(CLBLL_R_X75Y134_SLICE_X115Y134_AO6),
.I2(CLBLM_L_X76Y134_SLICE_X117Y134_AQ),
.I3(CLBLM_L_X76Y133_SLICE_X116Y133_BQ),
.I4(CLBLM_L_X76Y134_SLICE_X116Y134_AQ),
.I5(CLBLL_R_X75Y133_SLICE_X115Y133_AQ),
.O5(CLBLM_L_X76Y134_SLICE_X117Y134_CO5),
.O6(CLBLM_L_X76Y134_SLICE_X117Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9c9cf0f08888f0f0)
  ) CLBLM_L_X76Y134_SLICE_X117Y134_BLUT (
.I0(CLBLM_L_X76Y134_SLICE_X116Y134_CO6),
.I1(CLBLM_L_X76Y134_SLICE_X117Y134_BQ),
.I2(CLBLM_L_X76Y134_SLICE_X117Y134_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X76Y134_SLICE_X117Y134_CO6),
.O5(CLBLM_L_X76Y134_SLICE_X117Y134_BO5),
.O6(CLBLM_L_X76Y134_SLICE_X117Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a5ff00a0a0ff00)
  ) CLBLM_L_X76Y134_SLICE_X117Y134_ALUT (
.I0(CLBLM_L_X76Y134_SLICE_X116Y134_CO6),
.I1(1'b1),
.I2(CLBLM_L_X76Y134_SLICE_X117Y134_AQ),
.I3(CLBLM_L_X76Y134_SLICE_X116Y134_BQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X76Y134_SLICE_X117Y134_CO6),
.O5(CLBLM_L_X76Y134_SLICE_X117Y134_AO5),
.O6(CLBLM_L_X76Y134_SLICE_X117Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X78Y104_SLICE_X120Y104_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X78Y104_SLICE_X120Y104_AO5),
.Q(CLBLM_L_X78Y104_SLICE_X120Y104_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X78Y104_SLICE_X120Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X78Y104_SLICE_X120Y104_AO6),
.Q(CLBLM_L_X78Y104_SLICE_X120Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X78Y104_SLICE_X120Y104_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X78Y104_SLICE_X120Y104_A5Q),
.Q(CLBLM_L_X78Y104_SLICE_X120Y104_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y104_SLICE_X120Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y104_SLICE_X120Y104_DO5),
.O6(CLBLM_L_X78Y104_SLICE_X120Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y104_SLICE_X120Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y104_SLICE_X120Y104_CO5),
.O6(CLBLM_L_X78Y104_SLICE_X120Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y104_SLICE_X120Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y104_SLICE_X120Y104_BO5),
.O6(CLBLM_L_X78Y104_SLICE_X120Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0faa0faa00f033f0)
  ) CLBLM_L_X78Y104_SLICE_X120Y104_ALUT (
.I0(CLBLM_L_X74Y121_SLICE_X113Y121_B5Q),
.I1(CLBLM_L_X78Y104_SLICE_X120Y104_BQ),
.I2(CLBLM_L_X78Y104_SLICE_X120Y104_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X78Y104_SLICE_X120Y104_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X78Y104_SLICE_X120Y104_AO5),
.O6(CLBLM_L_X78Y104_SLICE_X120Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y104_SLICE_X121Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y104_SLICE_X121Y104_DO5),
.O6(CLBLM_L_X78Y104_SLICE_X121Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y104_SLICE_X121Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y104_SLICE_X121Y104_CO5),
.O6(CLBLM_L_X78Y104_SLICE_X121Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y104_SLICE_X121Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y104_SLICE_X121Y104_BO5),
.O6(CLBLM_L_X78Y104_SLICE_X121Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y104_SLICE_X121Y104_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y104_SLICE_X121Y104_AO5),
.O6(CLBLM_L_X78Y104_SLICE_X121Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X78Y106_SLICE_X120Y106_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X72Y106_SLICE_X108Y106_AQ),
.Q(CLBLM_L_X78Y106_SLICE_X120Y106_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y106_SLICE_X120Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y106_SLICE_X120Y106_DO5),
.O6(CLBLM_L_X78Y106_SLICE_X120Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y106_SLICE_X120Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y106_SLICE_X120Y106_CO5),
.O6(CLBLM_L_X78Y106_SLICE_X120Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y106_SLICE_X120Y106_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y106_SLICE_X120Y106_BO5),
.O6(CLBLM_L_X78Y106_SLICE_X120Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y106_SLICE_X120Y106_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y106_SLICE_X120Y106_AO5),
.O6(CLBLM_L_X78Y106_SLICE_X120Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y106_SLICE_X121Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y106_SLICE_X121Y106_DO5),
.O6(CLBLM_L_X78Y106_SLICE_X121Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y106_SLICE_X121Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y106_SLICE_X121Y106_CO5),
.O6(CLBLM_L_X78Y106_SLICE_X121Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y106_SLICE_X121Y106_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y106_SLICE_X121Y106_BO5),
.O6(CLBLM_L_X78Y106_SLICE_X121Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y106_SLICE_X121Y106_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y106_SLICE_X121Y106_AO5),
.O6(CLBLM_L_X78Y106_SLICE_X121Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X78Y120_SLICE_X120Y120_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X78Y120_SLICE_X120Y120_AO6),
.Q(CLBLM_L_X78Y120_SLICE_X120Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y120_SLICE_X120Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y120_SLICE_X120Y120_DO5),
.O6(CLBLM_L_X78Y120_SLICE_X120Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y120_SLICE_X120Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y120_SLICE_X120Y120_CO5),
.O6(CLBLM_L_X78Y120_SLICE_X120Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y120_SLICE_X120Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y120_SLICE_X120Y120_BO5),
.O6(CLBLM_L_X78Y120_SLICE_X120Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb400b4b4cccccccc)
  ) CLBLM_L_X78Y120_SLICE_X120Y120_ALUT (
.I0(CLBLM_L_X78Y121_SLICE_X120Y121_CO6),
.I1(CLBLM_L_X78Y122_SLICE_X121Y122_AQ),
.I2(CLBLM_L_X78Y120_SLICE_X120Y120_AQ),
.I3(CLBLM_L_X76Y122_SLICE_X117Y122_AQ),
.I4(CLBLL_R_X77Y113_SLICE_X118Y113_AQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X78Y120_SLICE_X120Y120_AO5),
.O6(CLBLM_L_X78Y120_SLICE_X120Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y120_SLICE_X121Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y120_SLICE_X121Y120_DO5),
.O6(CLBLM_L_X78Y120_SLICE_X121Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y120_SLICE_X121Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y120_SLICE_X121Y120_CO5),
.O6(CLBLM_L_X78Y120_SLICE_X121Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y120_SLICE_X121Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y120_SLICE_X121Y120_BO5),
.O6(CLBLM_L_X78Y120_SLICE_X121Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y120_SLICE_X121Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y120_SLICE_X121Y120_AO5),
.O6(CLBLM_L_X78Y120_SLICE_X121Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X78Y121_SLICE_X120Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X78Y121_SLICE_X120Y121_AO6),
.Q(CLBLM_L_X78Y121_SLICE_X120Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X78Y121_SLICE_X120Y121_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X78Y121_SLICE_X120Y121_BO6),
.Q(CLBLM_L_X78Y121_SLICE_X120Y121_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y121_SLICE_X120Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y121_SLICE_X120Y121_DO5),
.O6(CLBLM_L_X78Y121_SLICE_X120Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3fbf33bb33bb)
  ) CLBLM_L_X78Y121_SLICE_X120Y121_CLUT (
.I0(CLBLL_R_X77Y113_SLICE_X118Y113_AQ),
.I1(CLBLM_L_X78Y121_SLICE_X120Y121_AQ),
.I2(CLBLM_L_X78Y121_SLICE_X120Y121_BQ),
.I3(CLBLM_L_X76Y122_SLICE_X117Y122_AQ),
.I4(CLBLM_L_X78Y123_SLICE_X120Y123_BO6),
.I5(1'b1),
.O5(CLBLM_L_X78Y121_SLICE_X120Y121_CO5),
.O6(CLBLM_L_X78Y121_SLICE_X120Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9c009c9cf0f0f0f0)
  ) CLBLM_L_X78Y121_SLICE_X120Y121_BLUT (
.I0(CLBLM_L_X78Y123_SLICE_X120Y123_BO6),
.I1(CLBLM_L_X78Y121_SLICE_X120Y121_BQ),
.I2(CLBLM_L_X78Y121_SLICE_X120Y121_AQ),
.I3(CLBLM_L_X76Y122_SLICE_X117Y122_AQ),
.I4(CLBLL_R_X77Y113_SLICE_X118Y113_AQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X78Y121_SLICE_X120Y121_BO5),
.O6(CLBLM_L_X78Y121_SLICE_X120Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he44ee44e4444e44e)
  ) CLBLM_L_X78Y121_SLICE_X120Y121_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X78Y123_SLICE_X121Y123_BQ),
.I2(CLBLM_L_X78Y121_SLICE_X120Y121_AQ),
.I3(CLBLM_L_X78Y123_SLICE_X120Y123_BO6),
.I4(CLBLL_R_X77Y113_SLICE_X118Y113_AQ),
.I5(CLBLM_L_X76Y122_SLICE_X117Y122_AQ),
.O5(CLBLM_L_X78Y121_SLICE_X120Y121_AO5),
.O6(CLBLM_L_X78Y121_SLICE_X120Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y121_SLICE_X121Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y121_SLICE_X121Y121_DO5),
.O6(CLBLM_L_X78Y121_SLICE_X121Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y121_SLICE_X121Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y121_SLICE_X121Y121_CO5),
.O6(CLBLM_L_X78Y121_SLICE_X121Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y121_SLICE_X121Y121_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y121_SLICE_X121Y121_BO5),
.O6(CLBLM_L_X78Y121_SLICE_X121Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y121_SLICE_X121Y121_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y121_SLICE_X121Y121_AO5),
.O6(CLBLM_L_X78Y121_SLICE_X121Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffdfffffffff)
  ) CLBLM_L_X78Y122_SLICE_X120Y122_DLUT (
.I0(CLBLL_R_X77Y122_SLICE_X119Y122_BQ),
.I1(CLBLM_L_X78Y123_SLICE_X120Y123_CO6),
.I2(CLBLM_L_X78Y121_SLICE_X120Y121_BQ),
.I3(CLBLM_L_X78Y122_SLICE_X120Y122_AO5),
.I4(CLBLL_R_X77Y122_SLICE_X119Y122_AO5),
.I5(CLBLM_L_X78Y122_SLICE_X121Y122_BQ),
.O5(CLBLM_L_X78Y122_SLICE_X120Y122_DO5),
.O6(CLBLM_L_X78Y122_SLICE_X120Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff7fffffffff)
  ) CLBLM_L_X78Y122_SLICE_X120Y122_CLUT (
.I0(CLBLM_L_X78Y122_SLICE_X120Y122_AO6),
.I1(CLBLM_L_X78Y120_SLICE_X120Y120_AQ),
.I2(CLBLM_L_X78Y121_SLICE_X120Y121_BQ),
.I3(CLBLM_L_X78Y123_SLICE_X120Y123_CO6),
.I4(CLBLL_R_X77Y122_SLICE_X119Y122_AO5),
.I5(CLBLM_L_X78Y122_SLICE_X121Y122_BQ),
.O5(CLBLM_L_X78Y122_SLICE_X120Y122_CO5),
.O6(CLBLM_L_X78Y122_SLICE_X120Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffbfffffff)
  ) CLBLM_L_X78Y122_SLICE_X120Y122_BLUT (
.I0(CLBLM_L_X78Y123_SLICE_X121Y123_CO6),
.I1(CLBLM_L_X78Y121_SLICE_X120Y121_BQ),
.I2(CLBLM_L_X78Y120_SLICE_X120Y120_AQ),
.I3(CLBLM_L_X78Y122_SLICE_X121Y122_BQ),
.I4(CLBLM_L_X78Y122_SLICE_X121Y122_AQ),
.I5(CLBLM_L_X78Y123_SLICE_X120Y123_CO6),
.O5(CLBLM_L_X78Y122_SLICE_X120Y122_BO5),
.O6(CLBLM_L_X78Y122_SLICE_X120Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccff00003f0fffff)
  ) CLBLM_L_X78Y122_SLICE_X120Y122_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X76Y122_SLICE_X117Y122_AQ),
.I2(CLBLM_L_X78Y120_SLICE_X120Y120_AQ),
.I3(CLBLL_R_X77Y113_SLICE_X118Y113_AQ),
.I4(CLBLM_L_X78Y122_SLICE_X121Y122_AQ),
.I5(1'b1),
.O5(CLBLM_L_X78Y122_SLICE_X120Y122_AO5),
.O6(CLBLM_L_X78Y122_SLICE_X120Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X78Y122_SLICE_X121Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X78Y122_SLICE_X121Y122_AO6),
.Q(CLBLM_L_X78Y122_SLICE_X121Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X78Y122_SLICE_X121Y122_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X78Y122_SLICE_X121Y122_BO6),
.Q(CLBLM_L_X78Y122_SLICE_X121Y122_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y122_SLICE_X121Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y122_SLICE_X121Y122_DO5),
.O6(CLBLM_L_X78Y122_SLICE_X121Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y122_SLICE_X121Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y122_SLICE_X121Y122_CO5),
.O6(CLBLM_L_X78Y122_SLICE_X121Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55dd557d00880088)
  ) CLBLM_L_X78Y122_SLICE_X121Y122_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X78Y122_SLICE_X121Y122_BQ),
.I2(CLBLM_L_X78Y122_SLICE_X121Y122_AQ),
.I3(CLBLM_L_X78Y123_SLICE_X121Y123_CO6),
.I4(CLBLM_L_X78Y121_SLICE_X120Y121_CO6),
.I5(CLBLM_L_X78Y120_SLICE_X120Y120_AQ),
.O5(CLBLM_L_X78Y122_SLICE_X121Y122_BO5),
.O6(CLBLM_L_X78Y122_SLICE_X121Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha00ff00fcccccccc)
  ) CLBLM_L_X78Y122_SLICE_X121Y122_ALUT (
.I0(CLBLM_L_X76Y122_SLICE_X117Y122_AQ),
.I1(CLBLM_L_X78Y121_SLICE_X120Y121_BQ),
.I2(CLBLM_L_X78Y122_SLICE_X121Y122_AQ),
.I3(CLBLM_L_X78Y121_SLICE_X120Y121_CO6),
.I4(CLBLL_R_X77Y113_SLICE_X118Y113_AQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X78Y122_SLICE_X121Y122_AO5),
.O6(CLBLM_L_X78Y122_SLICE_X121Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffee)
  ) CLBLM_L_X78Y123_SLICE_X120Y123_DLUT (
.I0(CLBLM_L_X78Y124_SLICE_X120Y124_BQ),
.I1(CLBLM_L_X78Y124_SLICE_X120Y124_CQ),
.I2(1'b1),
.I3(CLBLM_L_X78Y124_SLICE_X120Y124_AQ),
.I4(CLBLL_R_X77Y124_SLICE_X118Y124_BQ),
.I5(CLBLL_R_X77Y123_SLICE_X118Y123_AQ),
.O5(CLBLM_L_X78Y123_SLICE_X120Y123_DO5),
.O6(CLBLM_L_X78Y123_SLICE_X120Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffefffffffff)
  ) CLBLM_L_X78Y123_SLICE_X120Y123_CLUT (
.I0(CLBLM_L_X78Y121_SLICE_X120Y121_CO5),
.I1(CLBLM_L_X78Y123_SLICE_X121Y123_CO5),
.I2(CLBLL_R_X75Y123_SLICE_X114Y123_AO6),
.I3(CLBLL_R_X77Y121_SLICE_X118Y121_AO6),
.I4(CLBLM_L_X78Y123_SLICE_X120Y123_DO6),
.I5(CLBLM_L_X78Y123_SLICE_X121Y123_BQ),
.O5(CLBLM_L_X78Y123_SLICE_X120Y123_CO5),
.O6(CLBLM_L_X78Y123_SLICE_X120Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbfffffffbfffbff)
  ) CLBLM_L_X78Y123_SLICE_X120Y123_BLUT (
.I0(CLBLM_L_X78Y123_SLICE_X120Y123_DO6),
.I1(CLBLL_R_X75Y123_SLICE_X114Y123_AO6),
.I2(CLBLL_R_X77Y121_SLICE_X118Y121_AO6),
.I3(CLBLM_L_X78Y123_SLICE_X121Y123_BQ),
.I4(CLBLL_R_X77Y113_SLICE_X118Y113_AQ),
.I5(CLBLM_L_X72Y111_SLICE_X108Y111_C5Q),
.O5(CLBLM_L_X78Y123_SLICE_X120Y123_BO5),
.O6(CLBLM_L_X78Y123_SLICE_X120Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000004)
  ) CLBLM_L_X78Y123_SLICE_X120Y123_ALUT (
.I0(CLBLM_L_X78Y124_SLICE_X120Y124_CQ),
.I1(CLBLL_R_X75Y123_SLICE_X114Y123_AO6),
.I2(CLBLL_R_X77Y124_SLICE_X118Y124_BQ),
.I3(CLBLM_L_X78Y124_SLICE_X120Y124_AQ),
.I4(CLBLM_L_X78Y124_SLICE_X120Y124_BQ),
.I5(CLBLL_R_X77Y123_SLICE_X118Y123_AQ),
.O5(CLBLM_L_X78Y123_SLICE_X120Y123_AO5),
.O6(CLBLM_L_X78Y123_SLICE_X120Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X78Y123_SLICE_X121Y123_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X78Y123_SLICE_X121Y123_AO5),
.Q(CLBLM_L_X78Y123_SLICE_X121Y123_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X78Y123_SLICE_X121Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X78Y123_SLICE_X121Y123_AO6),
.Q(CLBLM_L_X78Y123_SLICE_X121Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X78Y123_SLICE_X121Y123_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X78Y123_SLICE_X121Y123_BO6),
.Q(CLBLM_L_X78Y123_SLICE_X121Y123_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y123_SLICE_X121Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y123_SLICE_X121Y123_DO5),
.O6(CLBLM_L_X78Y123_SLICE_X121Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aaaa50505050)
  ) CLBLM_L_X78Y123_SLICE_X121Y123_CLUT (
.I0(CLBLL_R_X77Y113_SLICE_X118Y113_AQ),
.I1(1'b1),
.I2(CLBLM_L_X72Y111_SLICE_X108Y111_C5Q),
.I3(1'b1),
.I4(CLBLM_L_X76Y122_SLICE_X117Y122_AQ),
.I5(1'b1),
.O5(CLBLM_L_X78Y123_SLICE_X121Y123_CO5),
.O6(CLBLM_L_X78Y123_SLICE_X121Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8c8caaaa2c23aaaa)
  ) CLBLM_L_X78Y123_SLICE_X121Y123_BLUT (
.I0(CLBLM_L_X76Y122_SLICE_X117Y122_AQ),
.I1(CLBLM_L_X78Y123_SLICE_X121Y123_BQ),
.I2(CLBLL_R_X77Y113_SLICE_X118Y113_AQ),
.I3(CLBLM_L_X72Y111_SLICE_X108Y111_C5Q),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X77Y123_SLICE_X119Y123_BO5),
.O5(CLBLM_L_X78Y123_SLICE_X121Y123_BO5),
.O6(CLBLM_L_X78Y123_SLICE_X121Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00a0aa0af0d8f0d8)
  ) CLBLM_L_X78Y123_SLICE_X121Y123_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X78Y123_SLICE_X121Y123_A5Q),
.I2(CLBLM_L_X78Y123_SLICE_X121Y123_AQ),
.I3(CLBLM_L_X78Y123_SLICE_X120Y123_AO6),
.I4(CLBLM_L_X78Y127_SLICE_X121Y127_DO6),
.I5(1'b1),
.O5(CLBLM_L_X78Y123_SLICE_X121Y123_AO5),
.O6(CLBLM_L_X78Y123_SLICE_X121Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X78Y124_SLICE_X120Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X78Y124_SLICE_X120Y124_AO6),
.Q(CLBLM_L_X78Y124_SLICE_X120Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X78Y124_SLICE_X120Y124_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X78Y124_SLICE_X120Y124_BO6),
.Q(CLBLM_L_X78Y124_SLICE_X120Y124_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X78Y124_SLICE_X120Y124_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X78Y124_SLICE_X120Y124_CO6),
.Q(CLBLM_L_X78Y124_SLICE_X120Y124_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y124_SLICE_X120Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y124_SLICE_X120Y124_DO5),
.O6(CLBLM_L_X78Y124_SLICE_X120Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaa0accccaaaa)
  ) CLBLM_L_X78Y124_SLICE_X120Y124_CLUT (
.I0(CLBLL_R_X77Y123_SLICE_X119Y123_AQ),
.I1(CLBLM_L_X78Y124_SLICE_X120Y124_CQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLL_R_X77Y123_SLICE_X119Y123_CQ),
.I4(CLBLM_L_X76Y123_SLICE_X117Y123_AO5),
.I5(CLBLM_L_X76Y124_SLICE_X117Y124_BQ),
.O5(CLBLM_L_X78Y124_SLICE_X120Y124_CO5),
.O6(CLBLM_L_X78Y124_SLICE_X120Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6cfff0f06c6cf0f0)
  ) CLBLM_L_X78Y124_SLICE_X120Y124_BLUT (
.I0(CLBLL_R_X77Y124_SLICE_X118Y124_CO6),
.I1(CLBLM_L_X78Y124_SLICE_X120Y124_BQ),
.I2(CLBLM_L_X78Y124_SLICE_X120Y124_AQ),
.I3(CLBLL_R_X77Y123_SLICE_X119Y123_CQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X76Y124_SLICE_X117Y124_BQ),
.O5(CLBLM_L_X78Y124_SLICE_X120Y124_BO5),
.O6(CLBLM_L_X78Y124_SLICE_X120Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7d7d2828ff7daa28)
  ) CLBLM_L_X78Y124_SLICE_X120Y124_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X77Y124_SLICE_X118Y124_CO6),
.I2(CLBLM_L_X78Y124_SLICE_X120Y124_AQ),
.I3(CLBLM_L_X76Y124_SLICE_X117Y124_BQ),
.I4(CLBLL_R_X77Y124_SLICE_X118Y124_BQ),
.I5(CLBLL_R_X77Y123_SLICE_X119Y123_CQ),
.O5(CLBLM_L_X78Y124_SLICE_X120Y124_AO5),
.O6(CLBLM_L_X78Y124_SLICE_X120Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y124_SLICE_X121Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y124_SLICE_X121Y124_DO5),
.O6(CLBLM_L_X78Y124_SLICE_X121Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y124_SLICE_X121Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y124_SLICE_X121Y124_CO5),
.O6(CLBLM_L_X78Y124_SLICE_X121Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y124_SLICE_X121Y124_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y124_SLICE_X121Y124_BO5),
.O6(CLBLM_L_X78Y124_SLICE_X121Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y124_SLICE_X121Y124_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y124_SLICE_X121Y124_AO5),
.O6(CLBLM_L_X78Y124_SLICE_X121Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y127_SLICE_X120Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y127_SLICE_X120Y127_DO5),
.O6(CLBLM_L_X78Y127_SLICE_X120Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y127_SLICE_X120Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y127_SLICE_X120Y127_CO5),
.O6(CLBLM_L_X78Y127_SLICE_X120Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y127_SLICE_X120Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y127_SLICE_X120Y127_BO5),
.O6(CLBLM_L_X78Y127_SLICE_X120Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y127_SLICE_X120Y127_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y127_SLICE_X120Y127_AO5),
.O6(CLBLM_L_X78Y127_SLICE_X120Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9966996666996699)
  ) CLBLM_L_X78Y127_SLICE_X121Y127_DLUT (
.I0(CLBLL_R_X79Y127_SLICE_X122Y127_AQ),
.I1(CLBLL_R_X79Y127_SLICE_X122Y127_BQ),
.I2(1'b1),
.I3(CLBLL_R_X79Y127_SLICE_X122Y127_DO6),
.I4(1'b1),
.I5(CLBLL_R_X79Y128_SLICE_X122Y128_BQ),
.O5(CLBLM_L_X78Y127_SLICE_X121Y127_DO5),
.O6(CLBLM_L_X78Y127_SLICE_X121Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0101010100000000)
  ) CLBLM_L_X78Y127_SLICE_X121Y127_CLUT (
.I0(CLBLM_L_X78Y127_SLICE_X121Y127_AO6),
.I1(CLBLL_R_X79Y127_SLICE_X122Y127_CQ),
.I2(CLBLL_R_X79Y128_SLICE_X122Y128_DQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_R_X79Y127_SLICE_X122Y127_AQ),
.O5(CLBLM_L_X78Y127_SLICE_X121Y127_CO5),
.O6(CLBLM_L_X78Y127_SLICE_X121Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00ff003f)
  ) CLBLM_L_X78Y127_SLICE_X121Y127_BLUT (
.I0(1'b1),
.I1(CLBLL_R_X79Y127_SLICE_X122Y127_CQ),
.I2(CLBLL_R_X79Y128_SLICE_X122Y128_DQ),
.I3(CLBLL_R_X77Y127_SLICE_X119Y127_AQ),
.I4(CLBLL_R_X79Y127_SLICE_X122Y127_AQ),
.I5(CLBLM_L_X78Y127_SLICE_X121Y127_AO5),
.O5(CLBLM_L_X78Y127_SLICE_X121Y127_BO5),
.O6(CLBLM_L_X78Y127_SLICE_X121Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbffffffffffffdd)
  ) CLBLM_L_X78Y127_SLICE_X121Y127_ALUT (
.I0(CLBLL_R_X79Y128_SLICE_X122Y128_CQ),
.I1(CLBLL_R_X79Y128_SLICE_X122Y128_BQ),
.I2(1'b1),
.I3(CLBLL_R_X79Y128_SLICE_X122Y128_AQ),
.I4(CLBLL_R_X79Y127_SLICE_X122Y127_BQ),
.I5(1'b1),
.O5(CLBLM_L_X78Y127_SLICE_X121Y127_AO5),
.O6(CLBLM_L_X78Y127_SLICE_X121Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X78Y128_SLICE_X120Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X78Y128_SLICE_X120Y128_AO6),
.Q(CLBLM_L_X78Y128_SLICE_X120Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y128_SLICE_X120Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y128_SLICE_X120Y128_DO5),
.O6(CLBLM_L_X78Y128_SLICE_X120Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y128_SLICE_X120Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y128_SLICE_X120Y128_CO5),
.O6(CLBLM_L_X78Y128_SLICE_X120Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y128_SLICE_X120Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y128_SLICE_X120Y128_BO5),
.O6(CLBLM_L_X78Y128_SLICE_X120Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfacc50ccfacc50cc)
  ) CLBLM_L_X78Y128_SLICE_X120Y128_ALUT (
.I0(CLBLL_R_X77Y128_SLICE_X119Y128_BQ),
.I1(CLBLL_R_X77Y128_SLICE_X118Y128_CQ),
.I2(CLBLM_L_X78Y128_SLICE_X120Y128_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLL_R_X77Y128_SLICE_X118Y128_BQ),
.I5(1'b1),
.O5(CLBLM_L_X78Y128_SLICE_X120Y128_AO5),
.O6(CLBLM_L_X78Y128_SLICE_X120Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y128_SLICE_X121Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y128_SLICE_X121Y128_DO5),
.O6(CLBLM_L_X78Y128_SLICE_X121Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y128_SLICE_X121Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y128_SLICE_X121Y128_CO5),
.O6(CLBLM_L_X78Y128_SLICE_X121Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y128_SLICE_X121Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y128_SLICE_X121Y128_BO5),
.O6(CLBLM_L_X78Y128_SLICE_X121Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y128_SLICE_X121Y128_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y128_SLICE_X121Y128_AO5),
.O6(CLBLM_L_X78Y128_SLICE_X121Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y129_SLICE_X120Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y129_SLICE_X120Y129_DO5),
.O6(CLBLM_L_X78Y129_SLICE_X120Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y129_SLICE_X120Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y129_SLICE_X120Y129_CO5),
.O6(CLBLM_L_X78Y129_SLICE_X120Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfffffcfcfffff)
  ) CLBLM_L_X78Y129_SLICE_X120Y129_BLUT (
.I0(1'b1),
.I1(CLBLL_R_X77Y128_SLICE_X119Y128_CQ),
.I2(CLBLL_R_X77Y128_SLICE_X118Y128_BQ),
.I3(1'b1),
.I4(CLBLM_L_X78Y128_SLICE_X120Y128_AQ),
.I5(1'b1),
.O5(CLBLM_L_X78Y129_SLICE_X120Y129_BO5),
.O6(CLBLM_L_X78Y129_SLICE_X120Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0002000000000030)
  ) CLBLM_L_X78Y129_SLICE_X120Y129_ALUT (
.I0(CLBLL_R_X77Y130_SLICE_X119Y130_AQ),
.I1(CLBLM_L_X78Y131_SLICE_X120Y131_AQ),
.I2(CLBLL_R_X77Y128_SLICE_X118Y128_AQ),
.I3(CLBLL_R_X77Y130_SLICE_X118Y130_AQ),
.I4(CLBLL_R_X77Y128_SLICE_X118Y128_BQ),
.I5(CLBLL_R_X77Y128_SLICE_X119Y128_A5Q),
.O5(CLBLM_L_X78Y129_SLICE_X120Y129_AO5),
.O6(CLBLM_L_X78Y129_SLICE_X120Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y129_SLICE_X121Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y129_SLICE_X121Y129_DO5),
.O6(CLBLM_L_X78Y129_SLICE_X121Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y129_SLICE_X121Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y129_SLICE_X121Y129_CO5),
.O6(CLBLM_L_X78Y129_SLICE_X121Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y129_SLICE_X121Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y129_SLICE_X121Y129_BO5),
.O6(CLBLM_L_X78Y129_SLICE_X121Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y129_SLICE_X121Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y129_SLICE_X121Y129_AO5),
.O6(CLBLM_L_X78Y129_SLICE_X121Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X78Y130_SLICE_X120Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X78Y130_SLICE_X120Y130_AO6),
.Q(CLBLM_L_X78Y130_SLICE_X120Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X78Y130_SLICE_X120Y130_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X78Y130_SLICE_X120Y130_BO6),
.Q(CLBLM_L_X78Y130_SLICE_X120Y130_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00330000005f00ff)
  ) CLBLM_L_X78Y130_SLICE_X120Y130_DLUT (
.I0(CLBLM_L_X78Y130_SLICE_X120Y130_BQ),
.I1(CLBLL_R_X77Y130_SLICE_X118Y130_BQ),
.I2(CLBLL_R_X77Y131_SLICE_X119Y131_AQ),
.I3(CLBLM_L_X78Y131_SLICE_X120Y131_AQ),
.I4(CLBLL_R_X77Y130_SLICE_X118Y130_AQ),
.I5(CLBLL_R_X77Y130_SLICE_X119Y130_AO6),
.O5(CLBLM_L_X78Y130_SLICE_X120Y130_DO5),
.O6(CLBLM_L_X78Y130_SLICE_X120Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7fff70077ff7700)
  ) CLBLM_L_X78Y130_SLICE_X120Y130_CLUT (
.I0(CLBLM_L_X78Y130_SLICE_X120Y130_BQ),
.I1(CLBLL_R_X77Y131_SLICE_X119Y131_AQ),
.I2(CLBLL_R_X77Y130_SLICE_X118Y130_BQ),
.I3(CLBLL_R_X77Y130_SLICE_X118Y130_AQ),
.I4(CLBLL_R_X77Y130_SLICE_X119Y130_AO5),
.I5(CLBLL_R_X77Y130_SLICE_X119Y130_AO6),
.O5(CLBLM_L_X78Y130_SLICE_X120Y130_CO5),
.O6(CLBLM_L_X78Y130_SLICE_X120Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h282828ccf0f0f0f0)
  ) CLBLM_L_X78Y130_SLICE_X120Y130_BLUT (
.I0(CLBLM_L_X78Y130_SLICE_X120Y130_DO6),
.I1(CLBLM_L_X78Y130_SLICE_X120Y130_BQ),
.I2(CLBLM_L_X78Y130_SLICE_X120Y130_AQ),
.I3(CLBLL_R_X77Y130_SLICE_X119Y130_AQ),
.I4(CLBLL_R_X77Y128_SLICE_X118Y128_AQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X78Y130_SLICE_X120Y130_BO5),
.O6(CLBLM_L_X78Y130_SLICE_X120Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a3838ff00ff00)
  ) CLBLM_L_X78Y130_SLICE_X120Y130_ALUT (
.I0(CLBLM_L_X78Y130_SLICE_X120Y130_DO6),
.I1(CLBLL_R_X77Y130_SLICE_X119Y130_AQ),
.I2(CLBLM_L_X78Y130_SLICE_X120Y130_AQ),
.I3(CLBLL_R_X77Y130_SLICE_X118Y130_AQ),
.I4(CLBLL_R_X77Y128_SLICE_X118Y128_AQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_L_X78Y130_SLICE_X120Y130_AO5),
.O6(CLBLM_L_X78Y130_SLICE_X120Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y130_SLICE_X121Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y130_SLICE_X121Y130_DO5),
.O6(CLBLM_L_X78Y130_SLICE_X121Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y130_SLICE_X121Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y130_SLICE_X121Y130_CO5),
.O6(CLBLM_L_X78Y130_SLICE_X121Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y130_SLICE_X121Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y130_SLICE_X121Y130_BO5),
.O6(CLBLM_L_X78Y130_SLICE_X121Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y130_SLICE_X121Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y130_SLICE_X121Y130_AO5),
.O6(CLBLM_L_X78Y130_SLICE_X121Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X78Y131_SLICE_X120Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X78Y131_SLICE_X120Y131_AO6),
.Q(CLBLM_L_X78Y131_SLICE_X120Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y131_SLICE_X120Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y131_SLICE_X120Y131_DO5),
.O6(CLBLM_L_X78Y131_SLICE_X120Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y131_SLICE_X120Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y131_SLICE_X120Y131_CO5),
.O6(CLBLM_L_X78Y131_SLICE_X120Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y131_SLICE_X120Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y131_SLICE_X120Y131_BO5),
.O6(CLBLM_L_X78Y131_SLICE_X120Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha2a2222222a0a2a0)
  ) CLBLM_L_X78Y131_SLICE_X120Y131_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X78Y130_SLICE_X120Y130_CO6),
.I2(CLBLM_L_X78Y131_SLICE_X120Y131_AQ),
.I3(CLBLL_R_X77Y130_SLICE_X119Y130_AQ),
.I4(CLBLL_R_X77Y128_SLICE_X118Y128_BQ),
.I5(CLBLL_R_X77Y128_SLICE_X118Y128_AQ),
.O5(CLBLM_L_X78Y131_SLICE_X120Y131_AO5),
.O6(CLBLM_L_X78Y131_SLICE_X120Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y131_SLICE_X121Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y131_SLICE_X121Y131_DO5),
.O6(CLBLM_L_X78Y131_SLICE_X121Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y131_SLICE_X121Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y131_SLICE_X121Y131_CO5),
.O6(CLBLM_L_X78Y131_SLICE_X121Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y131_SLICE_X121Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y131_SLICE_X121Y131_BO5),
.O6(CLBLM_L_X78Y131_SLICE_X121Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y131_SLICE_X121Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y131_SLICE_X121Y131_AO5),
.O6(CLBLM_L_X78Y131_SLICE_X121Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X80Y132_SLICE_X124Y132_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y128_SLICE_X119Y128_BQ),
.Q(CLBLM_L_X80Y132_SLICE_X124Y132_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X80Y132_SLICE_X124Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X80Y132_SLICE_X124Y132_DO5),
.O6(CLBLM_L_X80Y132_SLICE_X124Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X80Y132_SLICE_X124Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X80Y132_SLICE_X124Y132_CO5),
.O6(CLBLM_L_X80Y132_SLICE_X124Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X80Y132_SLICE_X124Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X80Y132_SLICE_X124Y132_BO5),
.O6(CLBLM_L_X80Y132_SLICE_X124Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X80Y132_SLICE_X124Y132_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X80Y132_SLICE_X124Y132_AO5),
.O6(CLBLM_L_X80Y132_SLICE_X124Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X80Y132_SLICE_X125Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X80Y132_SLICE_X125Y132_DO5),
.O6(CLBLM_L_X80Y132_SLICE_X125Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X80Y132_SLICE_X125Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X80Y132_SLICE_X125Y132_CO5),
.O6(CLBLM_L_X80Y132_SLICE_X125Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X80Y132_SLICE_X125Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X80Y132_SLICE_X125Y132_BO5),
.O6(CLBLM_L_X80Y132_SLICE_X125Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X80Y132_SLICE_X125Y132_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X80Y132_SLICE_X125Y132_AO5),
.O6(CLBLM_L_X80Y132_SLICE_X125Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X82Y98_SLICE_X128Y98_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X82Y98_SLICE_X128Y98_AO5),
.Q(CLBLM_L_X82Y98_SLICE_X128Y98_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X82Y98_SLICE_X128Y98_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X82Y98_SLICE_X128Y98_AO6),
.Q(CLBLM_L_X82Y98_SLICE_X128Y98_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X82Y98_SLICE_X128Y98_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X82Y98_SLICE_X128Y98_AQ),
.Q(CLBLM_L_X82Y98_SLICE_X128Y98_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X82Y98_SLICE_X128Y98_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X82Y98_SLICE_X128Y98_DO5),
.O6(CLBLM_L_X82Y98_SLICE_X128Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X82Y98_SLICE_X128Y98_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X82Y98_SLICE_X128Y98_CO5),
.O6(CLBLM_L_X82Y98_SLICE_X128Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X82Y98_SLICE_X128Y98_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X82Y98_SLICE_X128Y98_BO5),
.O6(CLBLM_L_X82Y98_SLICE_X128Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ff003c3ccccc)
  ) CLBLM_L_X82Y98_SLICE_X128Y98_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X82Y98_SLICE_X128Y98_BQ),
.I2(CLBLM_L_X82Y98_SLICE_X128Y98_AQ),
.I3(CLBLL_R_X77Y104_SLICE_X118Y104_AQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLM_L_X82Y98_SLICE_X128Y98_AO5),
.O6(CLBLM_L_X82Y98_SLICE_X128Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X82Y98_SLICE_X129Y98_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X82Y98_SLICE_X129Y98_DO5),
.O6(CLBLM_L_X82Y98_SLICE_X129Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X82Y98_SLICE_X129Y98_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X82Y98_SLICE_X129Y98_CO5),
.O6(CLBLM_L_X82Y98_SLICE_X129Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X82Y98_SLICE_X129Y98_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X82Y98_SLICE_X129Y98_BO5),
.O6(CLBLM_L_X82Y98_SLICE_X129Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X82Y98_SLICE_X129Y98_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X82Y98_SLICE_X129Y98_AO5),
.O6(CLBLM_L_X82Y98_SLICE_X129Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X82Y130_SLICE_X128Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y125_SLICE_X118Y125_AQ),
.Q(CLBLM_L_X82Y130_SLICE_X128Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X82Y130_SLICE_X128Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X82Y130_SLICE_X128Y130_DO5),
.O6(CLBLM_L_X82Y130_SLICE_X128Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X82Y130_SLICE_X128Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X82Y130_SLICE_X128Y130_CO5),
.O6(CLBLM_L_X82Y130_SLICE_X128Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X82Y130_SLICE_X128Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X82Y130_SLICE_X128Y130_BO5),
.O6(CLBLM_L_X82Y130_SLICE_X128Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X82Y130_SLICE_X128Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X82Y130_SLICE_X128Y130_AO5),
.O6(CLBLM_L_X82Y130_SLICE_X128Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X82Y130_SLICE_X129Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X82Y130_SLICE_X129Y130_DO5),
.O6(CLBLM_L_X82Y130_SLICE_X129Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X82Y130_SLICE_X129Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X82Y130_SLICE_X129Y130_CO5),
.O6(CLBLM_L_X82Y130_SLICE_X129Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X82Y130_SLICE_X129Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X82Y130_SLICE_X129Y130_BO5),
.O6(CLBLM_L_X82Y130_SLICE_X129Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X82Y130_SLICE_X129Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X82Y130_SLICE_X129Y130_AO5),
.O6(CLBLM_L_X82Y130_SLICE_X129Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X53Y122_SLICE_X80Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y122_SLICE_X95Y122_AQ),
.Q(CLBLM_R_X53Y122_SLICE_X80Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X53Y122_SLICE_X80Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X53Y122_SLICE_X80Y122_DO5),
.O6(CLBLM_R_X53Y122_SLICE_X80Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X53Y122_SLICE_X80Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X53Y122_SLICE_X80Y122_CO5),
.O6(CLBLM_R_X53Y122_SLICE_X80Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X53Y122_SLICE_X80Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X53Y122_SLICE_X80Y122_BO5),
.O6(CLBLM_R_X53Y122_SLICE_X80Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X53Y122_SLICE_X80Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X53Y122_SLICE_X80Y122_AO5),
.O6(CLBLM_R_X53Y122_SLICE_X80Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X53Y122_SLICE_X81Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X53Y122_SLICE_X81Y122_DO5),
.O6(CLBLM_R_X53Y122_SLICE_X81Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X53Y122_SLICE_X81Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X53Y122_SLICE_X81Y122_CO5),
.O6(CLBLM_R_X53Y122_SLICE_X81Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X53Y122_SLICE_X81Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X53Y122_SLICE_X81Y122_BO5),
.O6(CLBLM_R_X53Y122_SLICE_X81Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X53Y122_SLICE_X81Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X53Y122_SLICE_X81Y122_AO5),
.O6(CLBLM_R_X53Y122_SLICE_X81Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y96_SLICE_X94Y96_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y96_SLICE_X94Y96_AO6),
.Q(CLBLM_R_X63Y96_SLICE_X94Y96_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y96_SLICE_X94Y96_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y96_SLICE_X94Y96_BO6),
.Q(CLBLM_R_X63Y96_SLICE_X94Y96_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y96_SLICE_X94Y96_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y96_SLICE_X94Y96_DO5),
.O6(CLBLM_R_X63Y96_SLICE_X94Y96_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y96_SLICE_X94Y96_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y96_SLICE_X94Y96_CO5),
.O6(CLBLM_R_X63Y96_SLICE_X94Y96_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8d8fad8d8d850)
  ) CLBLM_R_X63Y96_SLICE_X94Y96_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_R_X63Y96_SLICE_X94Y96_BQ),
.I2(CLBLM_R_X63Y96_SLICE_X94Y96_AQ),
.I3(CLBLM_L_X64Y97_SLICE_X97Y97_BO6),
.I4(CLBLM_R_X63Y99_SLICE_X94Y99_BO5),
.I5(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.O5(CLBLM_R_X63Y96_SLICE_X94Y96_BO5),
.O6(CLBLM_R_X63Y96_SLICE_X94Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f5ccccf0a0cccc)
  ) CLBLM_R_X63Y96_SLICE_X94Y96_ALUT (
.I0(CLBLM_R_X63Y99_SLICE_X94Y99_BO6),
.I1(CLBLM_L_X64Y97_SLICE_X96Y97_BQ),
.I2(CLBLM_R_X63Y96_SLICE_X94Y96_AQ),
.I3(CLBLM_L_X64Y97_SLICE_X97Y97_BO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.O5(CLBLM_R_X63Y96_SLICE_X94Y96_AO5),
.O6(CLBLM_R_X63Y96_SLICE_X94Y96_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y96_SLICE_X95Y96_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y96_SLICE_X95Y96_AO6),
.Q(CLBLM_R_X63Y96_SLICE_X95Y96_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y96_SLICE_X95Y96_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y96_SLICE_X95Y96_BO6),
.Q(CLBLM_R_X63Y96_SLICE_X95Y96_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y96_SLICE_X95Y96_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y96_SLICE_X95Y96_CO6),
.Q(CLBLM_R_X63Y96_SLICE_X95Y96_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y96_SLICE_X95Y96_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y96_SLICE_X95Y96_DO6),
.Q(CLBLM_R_X63Y96_SLICE_X95Y96_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aaaaf3c0aaaa)
  ) CLBLM_R_X63Y96_SLICE_X95Y96_DLUT (
.I0(CLBLM_R_X63Y96_SLICE_X95Y96_BQ),
.I1(CLBLM_R_X63Y99_SLICE_X94Y99_CO6),
.I2(CLBLM_R_X63Y96_SLICE_X95Y96_DQ),
.I3(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X64Y98_SLICE_X96Y98_AO6),
.O5(CLBLM_R_X63Y96_SLICE_X95Y96_DO5),
.O6(CLBLM_R_X63Y96_SLICE_X95Y96_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfdfc0d0cf8fc080)
  ) CLBLM_R_X63Y96_SLICE_X95Y96_CLUT (
.I0(CLBLM_L_X64Y97_SLICE_X97Y97_BO5),
.I1(CLBLM_R_X63Y96_SLICE_X95Y96_CQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_R_X63Y99_SLICE_X94Y99_CO6),
.I4(CLBLM_R_X63Y96_SLICE_X95Y96_AQ),
.I5(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.O5(CLBLM_R_X63Y96_SLICE_X95Y96_CO5),
.O6(CLBLM_R_X63Y96_SLICE_X95Y96_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffd5755aaa80200)
  ) CLBLM_R_X63Y96_SLICE_X95Y96_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X64Y98_SLICE_X96Y98_AO6),
.I2(CLBLM_R_X63Y99_SLICE_X94Y99_BO5),
.I3(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I4(CLBLM_R_X63Y96_SLICE_X95Y96_BQ),
.I5(CLBLM_L_X64Y97_SLICE_X96Y97_CQ),
.O5(CLBLM_R_X63Y96_SLICE_X95Y96_BO5),
.O6(CLBLM_R_X63Y96_SLICE_X95Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4eee4e4e444)
  ) CLBLM_R_X63Y96_SLICE_X95Y96_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X64Y97_SLICE_X96Y97_AQ),
.I2(CLBLM_R_X63Y96_SLICE_X95Y96_AQ),
.I3(CLBLM_L_X64Y97_SLICE_X97Y97_BO5),
.I4(CLBLM_R_X63Y99_SLICE_X94Y99_BO5),
.I5(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.O5(CLBLM_R_X63Y96_SLICE_X95Y96_AO5),
.O6(CLBLM_R_X63Y96_SLICE_X95Y96_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y97_SLICE_X94Y97_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y97_SLICE_X94Y97_AQ),
.Q(CLBLM_R_X63Y97_SLICE_X94Y97_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y97_SLICE_X94Y97_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y97_SLICE_X95Y97_AQ),
.Q(CLBLM_R_X63Y97_SLICE_X94Y97_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y97_SLICE_X94Y97_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y97_SLICE_X94Y97_BO6),
.Q(CLBLM_R_X63Y97_SLICE_X94Y97_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y97_SLICE_X94Y97_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y97_SLICE_X94Y97_B5Q),
.Q(CLBLM_R_X63Y97_SLICE_X94Y97_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfef0faf0fcf0f0f0)
  ) CLBLM_R_X63Y97_SLICE_X94Y97_DLUT (
.I0(CLBLM_R_X63Y97_SLICE_X95Y97_AQ),
.I1(CLBLM_L_X64Y98_SLICE_X96Y98_BQ),
.I2(CLBLM_R_X63Y97_SLICE_X95Y97_BO6),
.I3(CLBLM_R_X63Y97_SLICE_X94Y97_AO5),
.I4(CLBLM_L_X62Y99_SLICE_X93Y99_AQ),
.I5(CLBLM_R_X63Y96_SLICE_X95Y96_BQ),
.O5(CLBLM_R_X63Y97_SLICE_X94Y97_DO5),
.O6(CLBLM_R_X63Y97_SLICE_X94Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0002222c0000000)
  ) CLBLM_R_X63Y97_SLICE_X94Y97_CLUT (
.I0(CLBLM_L_X62Y97_SLICE_X93Y97_BQ),
.I1(CLBLM_R_X63Y99_SLICE_X95Y99_BQ),
.I2(CLBLM_R_X63Y98_SLICE_X94Y98_BQ),
.I3(CLBLM_L_X62Y97_SLICE_X93Y97_AQ),
.I4(CLBLM_R_X63Y99_SLICE_X95Y99_B5Q),
.I5(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.O5(CLBLM_R_X63Y97_SLICE_X94Y97_CO5),
.O6(CLBLM_R_X63Y97_SLICE_X94Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfd58a80dddd8888)
  ) CLBLM_R_X63Y97_SLICE_X94Y97_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_R_X63Y97_SLICE_X94Y97_BQ),
.I2(CLBLM_L_X64Y97_SLICE_X97Y97_BO6),
.I3(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I4(CLBLM_L_X62Y97_SLICE_X93Y97_BQ),
.I5(CLBLM_R_X63Y99_SLICE_X94Y99_A5Q),
.O5(CLBLM_R_X63Y97_SLICE_X94Y97_BO5),
.O6(CLBLM_R_X63Y97_SLICE_X94Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00200000cc00cc00)
  ) CLBLM_R_X63Y97_SLICE_X94Y97_ALUT (
.I0(CLBLM_L_X64Y97_SLICE_X97Y97_A5Q),
.I1(CLBLM_R_X63Y99_SLICE_X95Y99_B5Q),
.I2(CLBLM_L_X64Y97_SLICE_X96Y97_BQ),
.I3(CLBLM_R_X63Y99_SLICE_X95Y99_BQ),
.I4(CLBLM_R_X63Y97_SLICE_X94Y97_CQ),
.I5(1'b1),
.O5(CLBLM_R_X63Y97_SLICE_X94Y97_AO5),
.O6(CLBLM_R_X63Y97_SLICE_X94Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y97_SLICE_X95Y97_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y98_SLICE_X94Y98_AQ),
.Q(CLBLM_R_X63Y97_SLICE_X95Y97_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5050501050505050)
  ) CLBLM_R_X63Y97_SLICE_X95Y97_DLUT (
.I0(CLBLM_R_X63Y97_SLICE_X95Y97_AO6),
.I1(CLBLM_R_X63Y98_SLICE_X94Y98_AQ),
.I2(CLBLM_L_X64Y97_SLICE_X97Y97_A5Q),
.I3(CLBLM_R_X63Y99_SLICE_X95Y99_BQ),
.I4(CLBLM_R_X63Y99_SLICE_X95Y99_B5Q),
.I5(CLBLM_L_X64Y97_SLICE_X96Y97_AQ),
.O5(CLBLM_R_X63Y97_SLICE_X95Y97_DO5),
.O6(CLBLM_R_X63Y97_SLICE_X95Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5777ffff5fff)
  ) CLBLM_R_X63Y97_SLICE_X95Y97_CLUT (
.I0(CLBLM_R_X63Y99_SLICE_X95Y99_B5Q),
.I1(CLBLM_L_X60Y92_SLICE_X90Y92_BQ),
.I2(CLBLM_L_X64Y97_SLICE_X97Y97_DQ),
.I3(CLBLM_R_X63Y97_SLICE_X94Y97_B5Q),
.I4(CLBLM_R_X63Y99_SLICE_X95Y99_BQ),
.I5(CLBLM_R_X63Y97_SLICE_X94Y97_BQ),
.O5(CLBLM_R_X63Y97_SLICE_X95Y97_CO5),
.O6(CLBLM_R_X63Y97_SLICE_X95Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ec000000a000)
  ) CLBLM_R_X63Y97_SLICE_X95Y97_BLUT (
.I0(CLBLM_L_X64Y97_SLICE_X96Y97_CQ),
.I1(CLBLM_L_X64Y97_SLICE_X97Y97_CQ),
.I2(CLBLM_R_X63Y98_SLICE_X94Y98_AQ),
.I3(CLBLM_R_X63Y99_SLICE_X95Y99_BQ),
.I4(CLBLM_R_X63Y99_SLICE_X95Y99_B5Q),
.I5(CLBLM_R_X63Y97_SLICE_X94Y97_CQ),
.O5(CLBLM_R_X63Y97_SLICE_X95Y97_BO5),
.O6(CLBLM_R_X63Y97_SLICE_X95Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcca0000000a00000)
  ) CLBLM_R_X63Y97_SLICE_X95Y97_ALUT (
.I0(CLBLM_R_X63Y96_SLICE_X95Y96_AQ),
.I1(CLBLM_R_X63Y97_SLICE_X94Y97_B5Q),
.I2(CLBLM_R_X63Y97_SLICE_X95Y97_AQ),
.I3(CLBLM_R_X63Y99_SLICE_X95Y99_BQ),
.I4(CLBLM_R_X63Y99_SLICE_X95Y99_B5Q),
.I5(CLBLM_L_X64Y97_SLICE_X96Y97_DQ),
.O5(CLBLM_R_X63Y97_SLICE_X95Y97_AO5),
.O6(CLBLM_R_X63Y97_SLICE_X95Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y98_SLICE_X94Y98_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X60Y92_SLICE_X90Y92_BQ),
.Q(CLBLM_R_X63Y98_SLICE_X94Y98_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y98_SLICE_X94Y98_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y111_SLICE_X116Y111_BQ),
.Q(CLBLM_R_X63Y98_SLICE_X94Y98_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00c000c000aa0000)
  ) CLBLM_R_X63Y98_SLICE_X94Y98_DLUT (
.I0(CLBLM_L_X76Y111_SLICE_X116Y111_BQ),
.I1(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I2(CLBLM_L_X62Y98_SLICE_X93Y98_CQ),
.I3(CLBLM_R_X63Y99_SLICE_X95Y99_B5Q),
.I4(CLBLM_L_X62Y98_SLICE_X93Y98_AQ),
.I5(CLBLM_R_X63Y99_SLICE_X95Y99_BQ),
.O5(CLBLM_R_X63Y98_SLICE_X94Y98_DO5),
.O6(CLBLM_R_X63Y98_SLICE_X94Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeeeeeee4444444)
  ) CLBLM_R_X63Y98_SLICE_X94Y98_CLUT (
.I0(CLBLM_R_X63Y98_SLICE_X94Y98_AO6),
.I1(CLBLM_R_X63Y97_SLICE_X94Y97_CO6),
.I2(CLBLM_L_X62Y98_SLICE_X93Y98_BQ),
.I3(CLBLM_R_X63Y98_SLICE_X94Y98_BQ),
.I4(CLBLM_R_X63Y98_SLICE_X94Y98_BO5),
.I5(CLBLM_R_X63Y98_SLICE_X94Y98_DO6),
.O5(CLBLM_R_X63Y98_SLICE_X94Y98_CO5),
.O6(CLBLM_R_X63Y98_SLICE_X94Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2000000033003300)
  ) CLBLM_R_X63Y98_SLICE_X94Y98_BLUT (
.I0(CLBLM_L_X62Y99_SLICE_X93Y99_AQ),
.I1(CLBLM_R_X63Y99_SLICE_X95Y99_BQ),
.I2(CLBLM_L_X64Y97_SLICE_X97Y97_A5Q),
.I3(CLBLM_R_X63Y99_SLICE_X95Y99_B5Q),
.I4(CLBLM_R_X63Y96_SLICE_X94Y96_AQ),
.I5(1'b1),
.O5(CLBLM_R_X63Y98_SLICE_X94Y98_BO5),
.O6(CLBLM_R_X63Y98_SLICE_X94Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa55aa80800000)
  ) CLBLM_R_X63Y98_SLICE_X94Y98_ALUT (
.I0(CLBLM_L_X62Y99_SLICE_X93Y99_AQ),
.I1(CLBLM_R_X63Y98_SLICE_X94Y98_BQ),
.I2(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I3(CLBLM_L_X64Y97_SLICE_X97Y97_A5Q),
.I4(CLBLM_L_X76Y111_SLICE_X116Y111_BQ),
.I5(1'b1),
.O5(CLBLM_R_X63Y98_SLICE_X94Y98_AO5),
.O6(CLBLM_R_X63Y98_SLICE_X94Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y98_SLICE_X95Y98_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y98_SLICE_X95Y98_DO5),
.O6(CLBLM_R_X63Y98_SLICE_X95Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f000f000d000f0)
  ) CLBLM_R_X63Y98_SLICE_X95Y98_CLUT (
.I0(CLBLM_R_X63Y97_SLICE_X94Y97_AQ),
.I1(CLBLM_R_X63Y99_SLICE_X95Y99_B5Q),
.I2(CLBLM_R_X63Y97_SLICE_X95Y97_CO6),
.I3(CLBLM_L_X64Y97_SLICE_X97Y97_A5Q),
.I4(CLBLM_R_X63Y96_SLICE_X95Y96_DQ),
.I5(CLBLM_R_X63Y99_SLICE_X95Y99_BQ),
.O5(CLBLM_R_X63Y98_SLICE_X95Y98_CO5),
.O6(CLBLM_R_X63Y98_SLICE_X95Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffcfefffffccee)
  ) CLBLM_R_X63Y98_SLICE_X95Y98_BLUT (
.I0(CLBLM_R_X63Y99_SLICE_X95Y99_DO6),
.I1(CLBLM_R_X63Y98_SLICE_X94Y98_BO6),
.I2(CLBLM_R_X63Y99_SLICE_X95Y99_AO6),
.I3(CLBLM_L_X64Y98_SLICE_X96Y98_CO6),
.I4(CLBLM_R_X63Y97_SLICE_X94Y97_AO6),
.I5(CLBLM_L_X64Y99_SLICE_X96Y99_CQ),
.O5(CLBLM_R_X63Y98_SLICE_X95Y98_BO5),
.O6(CLBLM_R_X63Y98_SLICE_X95Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff20000fff30000)
  ) CLBLM_R_X63Y98_SLICE_X95Y98_ALUT (
.I0(CLBLM_R_X63Y97_SLICE_X94Y97_DO6),
.I1(CLBLM_R_X63Y97_SLICE_X95Y97_DO6),
.I2(CLBLM_R_X63Y98_SLICE_X94Y98_CO6),
.I3(CLBLM_R_X63Y98_SLICE_X95Y98_BO6),
.I4(CLBLM_L_X64Y103_SLICE_X97Y103_CO6),
.I5(CLBLM_R_X63Y98_SLICE_X95Y98_CO6),
.O5(CLBLM_R_X63Y98_SLICE_X95Y98_AO5),
.O6(CLBLM_R_X63Y98_SLICE_X95Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y99_SLICE_X94Y99_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y99_SLICE_X94Y99_AO5),
.Q(CLBLM_R_X63Y99_SLICE_X94Y99_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y99_SLICE_X94Y99_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y99_SLICE_X94Y99_DO5),
.Q(CLBLM_R_X63Y99_SLICE_X94Y99_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y99_SLICE_X94Y99_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y99_SLICE_X94Y99_AO6),
.Q(CLBLM_R_X63Y99_SLICE_X94Y99_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y99_SLICE_X94Y99_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y99_SLICE_X94Y99_DO6),
.Q(CLBLM_R_X63Y99_SLICE_X94Y99_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1133ff0050f0f0f0)
  ) CLBLM_R_X63Y99_SLICE_X94Y99_DLUT (
.I0(CLBLM_R_X63Y98_SLICE_X94Y98_AO5),
.I1(CLBLM_R_X63Y99_SLICE_X94Y99_D5Q),
.I2(CLBLM_R_X63Y99_SLICE_X94Y99_DQ),
.I3(CLBLM_L_X64Y97_SLICE_X97Y97_A5Q),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLM_R_X63Y99_SLICE_X94Y99_DO5),
.O6(CLBLM_R_X63Y99_SLICE_X94Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbbbbb77777777)
  ) CLBLM_R_X63Y99_SLICE_X94Y99_CLUT (
.I0(CLBLM_L_X64Y99_SLICE_X96Y99_AQ),
.I1(CLBLM_R_X63Y99_SLICE_X94Y99_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y99_SLICE_X94Y99_CO5),
.O6(CLBLM_R_X63Y99_SLICE_X94Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffcfcf0f0ffff)
  ) CLBLM_R_X63Y99_SLICE_X94Y99_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X63Y99_SLICE_X94Y99_A5Q),
.I2(CLBLM_R_X63Y99_SLICE_X94Y99_AQ),
.I3(1'b1),
.I4(CLBLM_L_X64Y99_SLICE_X96Y99_AQ),
.I5(1'b1),
.O5(CLBLM_R_X63Y99_SLICE_X94Y99_BO5),
.O6(CLBLM_R_X63Y99_SLICE_X94Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff0ff003000f0f0)
  ) CLBLM_R_X63Y99_SLICE_X94Y99_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X63Y99_SLICE_X94Y99_A5Q),
.I2(CLBLM_R_X63Y99_SLICE_X94Y99_AQ),
.I3(CLBLM_L_X64Y99_SLICE_X96Y99_AQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLM_R_X63Y99_SLICE_X94Y99_AO5),
.O6(CLBLM_R_X63Y99_SLICE_X94Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y99_SLICE_X95Y99_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y99_SLICE_X95Y99_BO5),
.Q(CLBLM_R_X63Y99_SLICE_X95Y99_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y99_SLICE_X95Y99_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y99_SLICE_X95Y99_BO6),
.Q(CLBLM_R_X63Y99_SLICE_X95Y99_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ff000000ff00)
  ) CLBLM_R_X63Y99_SLICE_X95Y99_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X63Y99_SLICE_X95Y99_BQ),
.I4(CLBLM_R_X63Y99_SLICE_X95Y99_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X63Y99_SLICE_X95Y99_DO5),
.O6(CLBLM_R_X63Y99_SLICE_X95Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8f4f8f4fcf0f0fc)
  ) CLBLM_R_X63Y99_SLICE_X95Y99_CLUT (
.I0(CLBLM_R_X63Y99_SLICE_X94Y99_D5Q),
.I1(CLBLM_L_X64Y103_SLICE_X97Y103_CO6),
.I2(CLBLM_L_X64Y102_SLICE_X97Y102_AQ),
.I3(CLBLM_R_X63Y99_SLICE_X95Y99_BQ),
.I4(CLBLM_R_X63Y99_SLICE_X94Y99_DQ),
.I5(CLBLM_R_X63Y99_SLICE_X95Y99_B5Q),
.O5(CLBLM_R_X63Y99_SLICE_X95Y99_CO5),
.O6(CLBLM_R_X63Y99_SLICE_X95Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6aca6aca5faf50a0)
  ) CLBLM_R_X63Y99_SLICE_X95Y99_BLUT (
.I0(CLBLM_R_X63Y99_SLICE_X95Y99_B5Q),
.I1(CLBLM_R_X63Y99_SLICE_X95Y99_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X64Y103_SLICE_X97Y103_CO6),
.I4(CLBLM_R_X63Y99_SLICE_X94Y99_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X63Y99_SLICE_X95Y99_BO5),
.O6(CLBLM_R_X63Y99_SLICE_X95Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f7fffff80000000)
  ) CLBLM_R_X63Y99_SLICE_X95Y99_ALUT (
.I0(CLBLM_R_X63Y99_SLICE_X95Y99_B5Q),
.I1(CLBLM_R_X63Y99_SLICE_X95Y99_BQ),
.I2(CLBLM_L_X60Y92_SLICE_X90Y92_BQ),
.I3(CLBLM_L_X64Y103_SLICE_X97Y103_CO6),
.I4(CLBLM_L_X64Y97_SLICE_X97Y97_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X63Y99_SLICE_X95Y99_AO5),
.O6(CLBLM_R_X63Y99_SLICE_X95Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y101_SLICE_X94Y101_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X60Y99_SLICE_X90Y99_CQ),
.Q(CLBLM_R_X63Y101_SLICE_X94Y101_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y101_SLICE_X94Y101_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y103_SLICE_X94Y103_AQ),
.Q(CLBLM_R_X63Y101_SLICE_X94Y101_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbfaffff00000000)
  ) CLBLM_R_X63Y101_SLICE_X94Y101_DLUT (
.I0(CLBLM_L_X62Y101_SLICE_X93Y101_DO6),
.I1(CLBLM_R_X63Y103_SLICE_X94Y103_CO6),
.I2(CLBLM_L_X62Y101_SLICE_X93Y101_CO6),
.I3(CLBLM_R_X63Y101_SLICE_X94Y101_AO5),
.I4(CLBLM_R_X63Y103_SLICE_X94Y103_DO6),
.I5(CLBLM_L_X64Y103_SLICE_X97Y103_DO6),
.O5(CLBLM_R_X63Y101_SLICE_X94Y101_DO5),
.O6(CLBLM_R_X63Y101_SLICE_X94Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ec000000a000)
  ) CLBLM_R_X63Y101_SLICE_X94Y101_CLUT (
.I0(CLBLM_R_X63Y101_SLICE_X94Y101_BQ),
.I1(CLBLM_R_X63Y101_SLICE_X94Y101_AQ),
.I2(CLBLM_R_X63Y102_SLICE_X95Y102_BQ),
.I3(CLBLM_L_X64Y101_SLICE_X96Y101_BQ),
.I4(CLBLM_L_X64Y101_SLICE_X96Y101_B5Q),
.I5(CLBLM_R_X63Y102_SLICE_X94Y102_AQ),
.O5(CLBLM_R_X63Y101_SLICE_X94Y101_CO5),
.O6(CLBLM_R_X63Y101_SLICE_X94Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000555580000000)
  ) CLBLM_R_X63Y101_SLICE_X94Y101_BLUT (
.I0(CLBLM_L_X64Y101_SLICE_X96Y101_B5Q),
.I1(CLBLM_L_X64Y103_SLICE_X97Y103_DO6),
.I2(CLBLM_L_X60Y99_SLICE_X90Y99_CQ),
.I3(CLBLM_L_X64Y101_SLICE_X96Y101_A5Q),
.I4(CLBLM_L_X64Y101_SLICE_X96Y101_BQ),
.I5(1'b1),
.O5(CLBLM_R_X63Y101_SLICE_X94Y101_BO5),
.O6(CLBLM_R_X63Y101_SLICE_X94Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000030303030)
  ) CLBLM_R_X63Y101_SLICE_X94Y101_ALUT (
.I0(CLBLM_R_X63Y102_SLICE_X95Y102_DQ),
.I1(CLBLM_L_X64Y101_SLICE_X96Y101_B5Q),
.I2(CLBLM_L_X64Y101_SLICE_X96Y101_BQ),
.I3(CLBLM_L_X64Y101_SLICE_X96Y101_A5Q),
.I4(CLBLM_L_X60Y99_SLICE_X90Y99_CQ),
.I5(1'b1),
.O5(CLBLM_R_X63Y101_SLICE_X94Y101_AO5),
.O6(CLBLM_R_X63Y101_SLICE_X94Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y101_SLICE_X95Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y101_SLICE_X95Y101_DO5),
.O6(CLBLM_R_X63Y101_SLICE_X95Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y101_SLICE_X95Y101_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y101_SLICE_X95Y101_CO5),
.O6(CLBLM_R_X63Y101_SLICE_X95Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y101_SLICE_X95Y101_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y101_SLICE_X95Y101_BO5),
.O6(CLBLM_R_X63Y101_SLICE_X95Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y101_SLICE_X95Y101_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y101_SLICE_X95Y101_AO5),
.O6(CLBLM_R_X63Y101_SLICE_X95Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y102_SLICE_X94Y102_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y102_SLICE_X94Y102_AO6),
.Q(CLBLM_R_X63Y102_SLICE_X94Y102_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y102_SLICE_X94Y102_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y102_SLICE_X94Y102_BO6),
.Q(CLBLM_R_X63Y102_SLICE_X94Y102_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fffaaaaffff)
  ) CLBLM_R_X63Y102_SLICE_X94Y102_DLUT (
.I0(CLBLM_R_X63Y102_SLICE_X95Y102_AQ),
.I1(1'b1),
.I2(CLBLM_L_X64Y105_SLICE_X96Y105_C5Q),
.I3(CLBLM_L_X64Y105_SLICE_X96Y105_CQ),
.I4(CLBLM_L_X64Y102_SLICE_X96Y102_AQ),
.I5(1'b1),
.O5(CLBLM_R_X63Y102_SLICE_X94Y102_DO5),
.O6(CLBLM_R_X63Y102_SLICE_X94Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfdfffdfffdfff)
  ) CLBLM_R_X63Y102_SLICE_X94Y102_CLUT (
.I0(CLBLM_R_X63Y102_SLICE_X95Y102_CQ),
.I1(CLBLM_L_X64Y101_SLICE_X96Y101_BQ),
.I2(CLBLM_L_X64Y101_SLICE_X96Y101_B5Q),
.I3(CLBLM_R_X63Y103_SLICE_X94Y103_AQ),
.I4(CLBLM_L_X62Y102_SLICE_X93Y102_AQ),
.I5(CLBLM_L_X60Y99_SLICE_X90Y99_CQ),
.O5(CLBLM_R_X63Y102_SLICE_X94Y102_CO5),
.O6(CLBLM_R_X63Y102_SLICE_X94Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0f0dd88f0f0)
  ) CLBLM_R_X63Y102_SLICE_X94Y102_BLUT (
.I0(CLBLM_L_X64Y102_SLICE_X96Y102_BO5),
.I1(CLBLM_R_X63Y102_SLICE_X94Y102_BQ),
.I2(CLBLM_R_X63Y102_SLICE_X94Y102_AQ),
.I3(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_R_X63Y103_SLICE_X94Y103_AO6),
.O5(CLBLM_R_X63Y102_SLICE_X94Y102_BO5),
.O6(CLBLM_R_X63Y102_SLICE_X94Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0ccaaaaaaaa)
  ) CLBLM_R_X63Y102_SLICE_X94Y102_ALUT (
.I0(CLBLM_L_X62Y102_SLICE_X93Y102_AQ),
.I1(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I2(CLBLM_R_X63Y102_SLICE_X94Y102_AQ),
.I3(CLBLM_R_X63Y102_SLICE_X95Y102_AO5),
.I4(CLBLM_L_X64Y102_SLICE_X96Y102_BO5),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_R_X63Y102_SLICE_X94Y102_AO5),
.O6(CLBLM_R_X63Y102_SLICE_X94Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y102_SLICE_X95Y102_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y102_SLICE_X95Y102_AO6),
.Q(CLBLM_R_X63Y102_SLICE_X95Y102_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y102_SLICE_X95Y102_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y102_SLICE_X95Y102_BO6),
.Q(CLBLM_R_X63Y102_SLICE_X95Y102_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y102_SLICE_X95Y102_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y102_SLICE_X95Y102_CO6),
.Q(CLBLM_R_X63Y102_SLICE_X95Y102_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y102_SLICE_X95Y102_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y102_SLICE_X95Y102_DO6),
.Q(CLBLM_R_X63Y102_SLICE_X95Y102_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaf0aa00aaf0aa)
  ) CLBLM_R_X63Y102_SLICE_X95Y102_DLUT (
.I0(CLBLM_L_X62Y102_SLICE_X92Y102_CQ),
.I1(1'b1),
.I2(CLBLM_R_X63Y102_SLICE_X95Y102_DQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_R_X63Y103_SLICE_X95Y103_BO5),
.I5(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.O5(CLBLM_R_X63Y102_SLICE_X95Y102_DO5),
.O6(CLBLM_R_X63Y102_SLICE_X95Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffacccc000acccc)
  ) CLBLM_R_X63Y102_SLICE_X95Y102_CLUT (
.I0(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I1(CLBLM_L_X64Y102_SLICE_X96Y102_CQ),
.I2(CLBLM_R_X63Y103_SLICE_X94Y103_AO5),
.I3(CLBLM_L_X64Y102_SLICE_X96Y102_BO5),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_R_X63Y102_SLICE_X95Y102_CQ),
.O5(CLBLM_R_X63Y102_SLICE_X95Y102_CO5),
.O6(CLBLM_R_X63Y102_SLICE_X95Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcecec4c4ff00ff00)
  ) CLBLM_R_X63Y102_SLICE_X95Y102_BLUT (
.I0(CLBLM_L_X64Y102_SLICE_X96Y102_A5Q),
.I1(CLBLM_R_X63Y102_SLICE_X95Y102_BQ),
.I2(CLBLM_L_X64Y102_SLICE_X96Y102_BO5),
.I3(CLBLM_R_X63Y102_SLICE_X95Y102_CQ),
.I4(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_R_X63Y102_SLICE_X95Y102_BO5),
.O6(CLBLM_R_X63Y102_SLICE_X95Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h04040404fffafffa)
  ) CLBLM_R_X63Y102_SLICE_X95Y102_ALUT (
.I0(CLBLM_L_X64Y102_SLICE_X96Y102_A5Q),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_R_X63Y102_SLICE_X95Y102_AQ),
.I3(CLBLM_L_X64Y102_SLICE_X96Y102_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y102_SLICE_X95Y102_AO5),
.O6(CLBLM_R_X63Y102_SLICE_X95Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y103_SLICE_X94Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y103_SLICE_X92Y103_B5Q),
.Q(CLBLM_R_X63Y103_SLICE_X94Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00100010ffff0010)
  ) CLBLM_R_X63Y103_SLICE_X94Y103_DLUT (
.I0(CLBLM_L_X62Y102_SLICE_X92Y102_DO6),
.I1(CLBLM_R_X63Y103_SLICE_X95Y103_CO6),
.I2(CLBLM_R_X63Y102_SLICE_X94Y102_CO6),
.I3(CLBLM_R_X63Y101_SLICE_X94Y101_CO6),
.I4(CLBLM_L_X62Y103_SLICE_X92Y103_CO6),
.I5(CLBLM_R_X63Y103_SLICE_X94Y103_BO6),
.O5(CLBLM_R_X63Y103_SLICE_X94Y103_DO5),
.O6(CLBLM_R_X63Y103_SLICE_X94Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h153f55ffcfcfffff)
  ) CLBLM_R_X63Y103_SLICE_X94Y103_CLUT (
.I0(CLBLM_L_X62Y103_SLICE_X92Y103_B5Q),
.I1(CLBLM_L_X62Y100_SLICE_X92Y100_AQ),
.I2(CLBLM_L_X62Y101_SLICE_X92Y101_AQ),
.I3(CLBLM_L_X62Y103_SLICE_X92Y103_BQ),
.I4(CLBLM_L_X62Y103_SLICE_X93Y103_CQ),
.I5(CLBLM_L_X64Y101_SLICE_X96Y101_A5Q),
.O5(CLBLM_R_X63Y103_SLICE_X94Y103_CO5),
.O6(CLBLM_R_X63Y103_SLICE_X94Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc022c00000220000)
  ) CLBLM_R_X63Y103_SLICE_X94Y103_BLUT (
.I0(CLBLM_R_X63Y103_SLICE_X95Y103_AQ),
.I1(CLBLM_L_X64Y101_SLICE_X96Y101_BQ),
.I2(CLBLM_R_X63Y103_SLICE_X94Y103_AQ),
.I3(CLBLM_L_X64Y101_SLICE_X96Y101_B5Q),
.I4(CLBLM_R_X63Y101_SLICE_X94Y101_AQ),
.I5(CLBLM_L_X62Y103_SLICE_X93Y103_DQ),
.O5(CLBLM_R_X63Y103_SLICE_X94Y103_BO5),
.O6(CLBLM_R_X63Y103_SLICE_X94Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0f0f0f0fffff)
  ) CLBLM_R_X63Y103_SLICE_X94Y103_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X63Y102_SLICE_X95Y102_AQ),
.I3(1'b1),
.I4(CLBLM_L_X64Y102_SLICE_X96Y102_AQ),
.I5(1'b1),
.O5(CLBLM_R_X63Y103_SLICE_X94Y103_AO5),
.O6(CLBLM_R_X63Y103_SLICE_X94Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y103_SLICE_X95Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y103_SLICE_X95Y103_AO6),
.Q(CLBLM_R_X63Y103_SLICE_X95Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y103_SLICE_X95Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y103_SLICE_X95Y103_DO5),
.O6(CLBLM_R_X63Y103_SLICE_X95Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00ff08ff08)
  ) CLBLM_R_X63Y103_SLICE_X95Y103_CLUT (
.I0(CLBLM_L_X62Y103_SLICE_X92Y103_B5Q),
.I1(CLBLM_L_X64Y102_SLICE_X96Y102_CQ),
.I2(CLBLM_L_X64Y101_SLICE_X96Y101_B5Q),
.I3(CLBLM_L_X64Y101_SLICE_X96Y101_A5Q),
.I4(1'b1),
.I5(CLBLM_L_X64Y101_SLICE_X96Y101_BQ),
.O5(CLBLM_R_X63Y103_SLICE_X95Y103_CO5),
.O6(CLBLM_R_X63Y103_SLICE_X95Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff00cc000000)
  ) CLBLM_R_X63Y103_SLICE_X95Y103_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X64Y102_SLICE_X96Y102_A5Q),
.I2(1'b1),
.I3(CLBLM_L_X64Y105_SLICE_X96Y105_C5Q),
.I4(CLBLM_L_X64Y105_SLICE_X96Y105_CQ),
.I5(1'b1),
.O5(CLBLM_R_X63Y103_SLICE_X95Y103_BO5),
.O6(CLBLM_R_X63Y103_SLICE_X95Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0e4aaaaaaaa)
  ) CLBLM_R_X63Y103_SLICE_X95Y103_ALUT (
.I0(CLBLM_L_X64Y105_SLICE_X96Y105_C5Q),
.I1(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I2(CLBLM_R_X63Y103_SLICE_X95Y103_AQ),
.I3(CLBLM_L_X64Y105_SLICE_X96Y105_CQ),
.I4(CLBLM_R_X63Y102_SLICE_X95Y102_AO5),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_R_X63Y103_SLICE_X95Y103_AO5),
.O6(CLBLM_R_X63Y103_SLICE_X95Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y105_SLICE_X94Y105_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y105_SLICE_X94Y105_CO5),
.Q(CLBLM_R_X63Y105_SLICE_X94Y105_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y105_SLICE_X94Y105_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y105_SLICE_X94Y105_AO6),
.Q(CLBLM_R_X63Y105_SLICE_X94Y105_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y105_SLICE_X94Y105_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y105_SLICE_X94Y105_BO6),
.Q(CLBLM_R_X63Y105_SLICE_X94Y105_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y105_SLICE_X94Y105_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y105_SLICE_X94Y105_CO6),
.Q(CLBLM_R_X63Y105_SLICE_X94Y105_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9111800080008000)
  ) CLBLM_R_X63Y105_SLICE_X94Y105_DLUT (
.I0(CLBLM_R_X63Y105_SLICE_X94Y105_C5Q),
.I1(CLBLM_R_X63Y105_SLICE_X94Y105_CQ),
.I2(CLBLM_L_X62Y107_SLICE_X93Y107_A5Q),
.I3(CLBLM_L_X62Y105_SLICE_X93Y105_BQ),
.I4(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I5(CLBLM_R_X63Y105_SLICE_X94Y105_AQ),
.O5(CLBLM_R_X63Y105_SLICE_X94Y105_DO5),
.O6(CLBLM_R_X63Y105_SLICE_X94Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h66aaccaa55f0aaf0)
  ) CLBLM_R_X63Y105_SLICE_X94Y105_CLUT (
.I0(CLBLM_R_X63Y105_SLICE_X94Y105_C5Q),
.I1(CLBLM_R_X63Y105_SLICE_X94Y105_CQ),
.I2(CLBLM_R_X63Y105_SLICE_X95Y105_C5Q),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X64Y105_SLICE_X97Y105_DO6),
.I5(1'b1),
.O5(CLBLM_R_X63Y105_SLICE_X94Y105_CO5),
.O6(CLBLM_R_X63Y105_SLICE_X94Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee4444ff00ff00)
  ) CLBLM_R_X63Y105_SLICE_X94Y105_BLUT (
.I0(CLBLM_L_X64Y106_SLICE_X97Y106_AO6),
.I1(CLBLM_R_X63Y105_SLICE_X94Y105_BQ),
.I2(1'b1),
.I3(CLBLM_R_X63Y105_SLICE_X95Y105_BQ),
.I4(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_R_X63Y105_SLICE_X94Y105_BO5),
.O6(CLBLM_R_X63Y105_SLICE_X94Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0ccf5cca0cc)
  ) CLBLM_R_X63Y105_SLICE_X94Y105_ALUT (
.I0(CLBLM_L_X64Y105_SLICE_X96Y105_AO6),
.I1(CLBLM_L_X62Y105_SLICE_X93Y105_BQ),
.I2(CLBLM_R_X63Y105_SLICE_X94Y105_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I5(CLBLM_L_X64Y106_SLICE_X96Y106_DO5),
.O5(CLBLM_R_X63Y105_SLICE_X94Y105_AO5),
.O6(CLBLM_R_X63Y105_SLICE_X94Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y105_SLICE_X95Y105_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y105_SLICE_X95Y105_AO5),
.Q(CLBLM_R_X63Y105_SLICE_X95Y105_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y105_SLICE_X95Y105_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y105_SLICE_X95Y105_CO5),
.Q(CLBLM_R_X63Y105_SLICE_X95Y105_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y105_SLICE_X95Y105_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y105_SLICE_X95Y105_AO6),
.Q(CLBLM_R_X63Y105_SLICE_X95Y105_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y105_SLICE_X95Y105_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y105_SLICE_X95Y105_BO6),
.Q(CLBLM_R_X63Y105_SLICE_X95Y105_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y105_SLICE_X95Y105_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y105_SLICE_X95Y105_CO6),
.Q(CLBLM_R_X63Y105_SLICE_X95Y105_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaaaaafaeabaeaba)
  ) CLBLM_R_X63Y105_SLICE_X95Y105_DLUT (
.I0(CLBLM_L_X64Y105_SLICE_X97Y105_BQ),
.I1(CLBLM_R_X63Y105_SLICE_X95Y105_CQ),
.I2(CLBLM_L_X64Y105_SLICE_X97Y105_DO6),
.I3(CLBLM_R_X63Y105_SLICE_X94Y105_CQ),
.I4(CLBLM_R_X63Y105_SLICE_X95Y105_C5Q),
.I5(CLBLM_R_X63Y105_SLICE_X94Y105_C5Q),
.O5(CLBLM_R_X63Y105_SLICE_X95Y105_DO5),
.O6(CLBLM_R_X63Y105_SLICE_X95Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f505f500ccccccc)
  ) CLBLM_R_X63Y105_SLICE_X95Y105_CLUT (
.I0(CLBLM_R_X63Y105_SLICE_X95Y105_C5Q),
.I1(CLBLM_R_X63Y105_SLICE_X95Y105_CQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_R_X63Y105_SLICE_X95Y105_A5Q),
.I4(CLBLM_L_X62Y107_SLICE_X93Y107_CO6),
.I5(1'b1),
.O5(CLBLM_R_X63Y105_SLICE_X95Y105_CO5),
.O6(CLBLM_R_X63Y105_SLICE_X95Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaaaaccf0aaaa)
  ) CLBLM_R_X63Y105_SLICE_X95Y105_BLUT (
.I0(CLBLM_R_X63Y107_SLICE_X95Y107_DQ),
.I1(CLBLM_R_X63Y105_SLICE_X95Y105_BQ),
.I2(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I3(CLBLM_L_X64Y106_SLICE_X96Y106_DO5),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_L_X64Y105_SLICE_X96Y105_BO6),
.O5(CLBLM_R_X63Y105_SLICE_X95Y105_BO5),
.O6(CLBLM_R_X63Y105_SLICE_X95Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff00f003a3acaca)
  ) CLBLM_R_X63Y105_SLICE_X95Y105_ALUT (
.I0(CLBLM_L_X64Y106_SLICE_X96Y106_BQ),
.I1(CLBLM_L_X62Y107_SLICE_X93Y107_CO6),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_R_X67Y103_SLICE_X100Y103_BQ),
.I4(CLBLM_R_X63Y105_SLICE_X95Y105_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X63Y105_SLICE_X95Y105_AO5),
.O6(CLBLM_R_X63Y105_SLICE_X95Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y106_SLICE_X94Y106_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y106_SLICE_X94Y106_BO6),
.Q(CLBLM_R_X63Y106_SLICE_X94Y106_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0ec00cc00cc00cc)
  ) CLBLM_R_X63Y106_SLICE_X94Y106_DLUT (
.I0(CLBLM_L_X62Y106_SLICE_X93Y106_BQ),
.I1(CLBLM_R_X63Y105_SLICE_X94Y105_BQ),
.I2(CLBLM_R_X63Y105_SLICE_X95Y105_A5Q),
.I3(CLBLM_R_X63Y106_SLICE_X94Y106_AO5),
.I4(CLBLM_L_X62Y106_SLICE_X93Y106_AO6),
.I5(CLBLM_L_X64Y106_SLICE_X96Y106_BQ),
.O5(CLBLM_R_X63Y106_SLICE_X94Y106_DO5),
.O6(CLBLM_R_X63Y106_SLICE_X94Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff07ffffff77ffff)
  ) CLBLM_R_X63Y106_SLICE_X94Y106_CLUT (
.I0(CLBLM_R_X63Y106_SLICE_X94Y106_BQ),
.I1(CLBLM_L_X60Y101_SLICE_X90Y101_BQ),
.I2(CLBLM_L_X64Y106_SLICE_X96Y106_A5Q),
.I3(CLBLM_R_X63Y105_SLICE_X94Y105_CQ),
.I4(CLBLM_R_X63Y105_SLICE_X94Y105_C5Q),
.I5(CLBLM_R_X63Y107_SLICE_X94Y107_BQ),
.O5(CLBLM_R_X63Y106_SLICE_X94Y106_CO5),
.O6(CLBLM_R_X63Y106_SLICE_X94Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00e4ffe400)
  ) CLBLM_R_X63Y106_SLICE_X94Y106_BLUT (
.I0(CLBLM_L_X64Y106_SLICE_X97Y106_C5Q),
.I1(CLBLM_R_X63Y106_SLICE_X94Y106_BQ),
.I2(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_R_X63Y105_SLICE_X94Y105_AQ),
.I5(CLBLM_L_X64Y105_SLICE_X96Y105_AO6),
.O5(CLBLM_R_X63Y106_SLICE_X94Y106_BO5),
.O6(CLBLM_R_X63Y106_SLICE_X94Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h800000007fff7fff)
  ) CLBLM_R_X63Y106_SLICE_X94Y106_ALUT (
.I0(CLBLM_R_X63Y105_SLICE_X94Y105_CQ),
.I1(CLBLM_R_X63Y105_SLICE_X94Y105_C5Q),
.I2(CLBLM_R_X63Y105_SLICE_X95Y105_A5Q),
.I3(CLBLM_L_X60Y101_SLICE_X90Y101_BQ),
.I4(CLBLM_L_X64Y105_SLICE_X97Y105_DO6),
.I5(1'b1),
.O5(CLBLM_R_X63Y106_SLICE_X94Y106_AO5),
.O6(CLBLM_R_X63Y106_SLICE_X94Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y106_SLICE_X95Y106_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y106_SLICE_X95Y106_AO6),
.Q(CLBLM_R_X63Y106_SLICE_X95Y106_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y106_SLICE_X95Y106_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y106_SLICE_X95Y106_BO6),
.Q(CLBLM_R_X63Y106_SLICE_X95Y106_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y106_SLICE_X95Y106_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y106_SLICE_X95Y106_CO6),
.Q(CLBLM_R_X63Y106_SLICE_X95Y106_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000eca00000)
  ) CLBLM_R_X63Y106_SLICE_X95Y106_DLUT (
.I0(CLBLM_R_X63Y107_SLICE_X95Y107_AQ),
.I1(CLBLM_R_X63Y106_SLICE_X95Y106_CQ),
.I2(CLBLM_L_X62Y106_SLICE_X93Y106_AQ),
.I3(CLBLM_L_X64Y106_SLICE_X96Y106_BQ),
.I4(CLBLM_R_X63Y105_SLICE_X94Y105_CQ),
.I5(CLBLM_R_X63Y105_SLICE_X94Y105_C5Q),
.O5(CLBLM_R_X63Y106_SLICE_X95Y106_DO5),
.O6(CLBLM_R_X63Y106_SLICE_X95Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hddfddd5d88a88808)
  ) CLBLM_R_X63Y106_SLICE_X95Y106_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_R_X63Y106_SLICE_X95Y106_CQ),
.I2(CLBLM_L_X64Y106_SLICE_X97Y106_C5Q),
.I3(CLBLM_L_X64Y105_SLICE_X96Y105_AO5),
.I4(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I5(CLBLM_R_X63Y107_SLICE_X94Y107_BQ),
.O5(CLBLM_R_X63Y106_SLICE_X95Y106_CO5),
.O6(CLBLM_R_X63Y106_SLICE_X95Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ddf0ccf088f0)
  ) CLBLM_R_X63Y106_SLICE_X95Y106_BLUT (
.I0(CLBLM_L_X64Y105_SLICE_X96Y105_AO6),
.I1(CLBLM_R_X63Y106_SLICE_X95Y106_BQ),
.I2(CLBLM_L_X62Y106_SLICE_X93Y106_BQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X64Y106_SLICE_X96Y106_BO6),
.I5(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.O5(CLBLM_R_X63Y106_SLICE_X95Y106_BO5),
.O6(CLBLM_R_X63Y106_SLICE_X95Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccffcc00ccf0cc)
  ) CLBLM_R_X63Y106_SLICE_X95Y106_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X63Y105_SLICE_X94Y105_BQ),
.I2(CLBLM_R_X63Y106_SLICE_X95Y106_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X64Y105_SLICE_X97Y105_DO6),
.I5(CLBLM_L_X62Y106_SLICE_X93Y106_DO6),
.O5(CLBLM_R_X63Y106_SLICE_X95Y106_AO5),
.O6(CLBLM_R_X63Y106_SLICE_X95Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y107_SLICE_X94Y107_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y107_SLICE_X94Y107_AO6),
.Q(CLBLM_R_X63Y107_SLICE_X94Y107_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y107_SLICE_X94Y107_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y107_SLICE_X94Y107_BO6),
.Q(CLBLM_R_X63Y107_SLICE_X94Y107_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5000000050000000)
  ) CLBLM_R_X63Y107_SLICE_X94Y107_DLUT (
.I0(CLBLM_R_X63Y105_SLICE_X94Y105_CQ),
.I1(1'b1),
.I2(CLBLM_L_X62Y107_SLICE_X93Y107_A5Q),
.I3(CLBLM_R_X63Y105_SLICE_X94Y105_C5Q),
.I4(CLBLM_R_X63Y107_SLICE_X95Y107_DQ),
.I5(1'b1),
.O5(CLBLM_R_X63Y107_SLICE_X94Y107_DO5),
.O6(CLBLM_R_X63Y107_SLICE_X94Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffa000cccccccc)
  ) CLBLM_R_X63Y107_SLICE_X94Y107_CLUT (
.I0(CLBLL_R_X75Y107_SLICE_X114Y107_AQ),
.I1(CLBLM_R_X63Y105_SLICE_X94Y105_DO6),
.I2(CLBLM_L_X62Y106_SLICE_X93Y106_AO6),
.I3(CLBLM_R_X63Y107_SLICE_X95Y107_CQ),
.I4(CLBLM_R_X63Y107_SLICE_X94Y107_DO6),
.I5(CLBLM_L_X62Y107_SLICE_X93Y107_CO5),
.O5(CLBLM_R_X63Y107_SLICE_X94Y107_CO5),
.O6(CLBLM_R_X63Y107_SLICE_X94Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccf0ddf088f0)
  ) CLBLM_R_X63Y107_SLICE_X94Y107_BLUT (
.I0(CLBLM_L_X64Y105_SLICE_X96Y105_AO5),
.I1(CLBLM_R_X63Y107_SLICE_X94Y107_BQ),
.I2(CLBLM_R_X63Y107_SLICE_X94Y107_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I5(CLBLM_L_X64Y106_SLICE_X96Y106_DO5),
.O5(CLBLM_R_X63Y107_SLICE_X94Y107_BO5),
.O6(CLBLM_R_X63Y107_SLICE_X94Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3c0f3c0f7c4b380)
  ) CLBLM_R_X63Y107_SLICE_X94Y107_ALUT (
.I0(CLBLM_L_X64Y105_SLICE_X96Y105_AO5),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_R_X63Y107_SLICE_X94Y107_AQ),
.I3(CLBLM_R_X63Y107_SLICE_X95Y107_BQ),
.I4(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I5(CLBLM_L_X64Y106_SLICE_X96Y106_DO6),
.O5(CLBLM_R_X63Y107_SLICE_X94Y107_AO5),
.O6(CLBLM_R_X63Y107_SLICE_X94Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y107_SLICE_X95Y107_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y107_SLICE_X95Y107_AO6),
.Q(CLBLM_R_X63Y107_SLICE_X95Y107_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y107_SLICE_X95Y107_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y107_SLICE_X95Y107_BO6),
.Q(CLBLM_R_X63Y107_SLICE_X95Y107_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y107_SLICE_X95Y107_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y107_SLICE_X95Y107_CO6),
.Q(CLBLM_R_X63Y107_SLICE_X95Y107_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y107_SLICE_X95Y107_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y107_SLICE_X95Y107_DO6),
.Q(CLBLM_R_X63Y107_SLICE_X95Y107_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0e2fffff0e20000)
  ) CLBLM_R_X63Y107_SLICE_X95Y107_DLUT (
.I0(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I1(CLBLM_L_X64Y105_SLICE_X96Y105_BO6),
.I2(CLBLM_R_X63Y107_SLICE_X95Y107_DQ),
.I3(CLBLM_L_X64Y106_SLICE_X96Y106_DO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_R_X63Y107_SLICE_X95Y107_CQ),
.O5(CLBLM_R_X63Y107_SLICE_X95Y107_DO5),
.O6(CLBLM_R_X63Y107_SLICE_X95Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffacccc0050cccc)
  ) CLBLM_R_X63Y107_SLICE_X95Y107_CLUT (
.I0(CLBLM_L_X64Y106_SLICE_X96Y106_BO5),
.I1(CLBLM_L_X64Y106_SLICE_X96Y106_CQ),
.I2(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I3(CLBLM_L_X64Y105_SLICE_X96Y105_BO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_R_X63Y107_SLICE_X95Y107_CQ),
.O5(CLBLM_R_X63Y107_SLICE_X95Y107_CO5),
.O6(CLBLM_R_X63Y107_SLICE_X95Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccdd88f0f0f0f0)
  ) CLBLM_R_X63Y107_SLICE_X95Y107_BLUT (
.I0(CLBLM_L_X64Y105_SLICE_X96Y105_AO5),
.I1(CLBLM_R_X63Y107_SLICE_X95Y107_BQ),
.I2(CLBLM_R_X63Y107_SLICE_X95Y107_AQ),
.I3(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I4(CLBLM_L_X64Y106_SLICE_X96Y106_BO5),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_R_X63Y107_SLICE_X95Y107_BO5),
.O6(CLBLM_R_X63Y107_SLICE_X95Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f7f3b3c0c4c080)
  ) CLBLM_R_X63Y107_SLICE_X95Y107_ALUT (
.I0(CLBLM_L_X64Y105_SLICE_X96Y105_AO5),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_R_X63Y107_SLICE_X95Y107_AQ),
.I3(CLBLM_L_X64Y106_SLICE_X96Y106_BO6),
.I4(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I5(CLBLM_R_X63Y106_SLICE_X94Y106_BQ),
.O5(CLBLM_R_X63Y107_SLICE_X95Y107_AO5),
.O6(CLBLM_R_X63Y107_SLICE_X95Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y122_SLICE_X94Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y122_SLICE_X94Y122_DO5),
.O6(CLBLM_R_X63Y122_SLICE_X94Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y122_SLICE_X94Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y122_SLICE_X94Y122_CO5),
.O6(CLBLM_R_X63Y122_SLICE_X94Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y122_SLICE_X94Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y122_SLICE_X94Y122_BO5),
.O6(CLBLM_R_X63Y122_SLICE_X94Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y122_SLICE_X94Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y122_SLICE_X94Y122_AO5),
.O6(CLBLM_R_X63Y122_SLICE_X94Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y122_SLICE_X95Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X64Y122_SLICE_X96Y122_AQ),
.Q(CLBLM_R_X63Y122_SLICE_X95Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y122_SLICE_X95Y122_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X76Y109_SLICE_X116Y109_AO6),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X53Y122_SLICE_X80Y122_AQ),
.Q(CLBLM_R_X63Y122_SLICE_X95Y122_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y122_SLICE_X95Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y122_SLICE_X95Y122_DO5),
.O6(CLBLM_R_X63Y122_SLICE_X95Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y122_SLICE_X95Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y122_SLICE_X95Y122_CO5),
.O6(CLBLM_R_X63Y122_SLICE_X95Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y122_SLICE_X95Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y122_SLICE_X95Y122_BO5),
.O6(CLBLM_R_X63Y122_SLICE_X95Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y122_SLICE_X95Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y122_SLICE_X95Y122_AO5),
.O6(CLBLM_R_X63Y122_SLICE_X95Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y99_SLICE_X98Y99_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y99_SLICE_X98Y99_AO6),
.Q(CLBLM_R_X65Y99_SLICE_X98Y99_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y99_SLICE_X98Y99_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y99_SLICE_X98Y99_BO6),
.Q(CLBLM_R_X65Y99_SLICE_X98Y99_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y99_SLICE_X98Y99_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y99_SLICE_X98Y99_CO6),
.Q(CLBLM_R_X65Y99_SLICE_X98Y99_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y99_SLICE_X98Y99_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y99_SLICE_X98Y99_DO5),
.O6(CLBLM_R_X65Y99_SLICE_X98Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4b00c300c300c300)
  ) CLBLM_R_X65Y99_SLICE_X98Y99_CLUT (
.I0(CLBLM_L_X64Y99_SLICE_X96Y99_BQ),
.I1(CLBLM_R_X65Y99_SLICE_X98Y99_CQ),
.I2(CLBLL_R_X79Y99_SLICE_X122Y99_AO6),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X64Y99_SLICE_X96Y99_A5Q),
.I5(CLBLM_R_X63Y99_SLICE_X94Y99_A5Q),
.O5(CLBLM_R_X65Y99_SLICE_X98Y99_CO5),
.O6(CLBLM_R_X65Y99_SLICE_X98Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he4ccccccf0f0f0f0)
  ) CLBLM_R_X65Y99_SLICE_X98Y99_BLUT (
.I0(CLBLM_L_X64Y99_SLICE_X96Y99_A5Q),
.I1(CLBLM_R_X65Y99_SLICE_X98Y99_BQ),
.I2(CLBLM_R_X65Y99_SLICE_X98Y99_CQ),
.I3(CLBLM_R_X63Y99_SLICE_X94Y99_A5Q),
.I4(CLBLM_L_X64Y99_SLICE_X96Y99_BQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_R_X65Y99_SLICE_X98Y99_BO5),
.O6(CLBLM_R_X65Y99_SLICE_X98Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaacc5acc5acc)
  ) CLBLM_R_X65Y99_SLICE_X98Y99_ALUT (
.I0(CLBLM_R_X63Y98_SLICE_X95Y98_AO6),
.I1(CLBLM_R_X65Y99_SLICE_X98Y99_BQ),
.I2(CLBLM_R_X65Y99_SLICE_X98Y99_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(1'b1),
.I5(CLBLM_R_X63Y99_SLICE_X95Y99_AO5),
.O5(CLBLM_R_X65Y99_SLICE_X98Y99_AO5),
.O6(CLBLM_R_X65Y99_SLICE_X98Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y99_SLICE_X99Y99_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y99_SLICE_X99Y99_CO5),
.Q(CLBLM_R_X65Y99_SLICE_X99Y99_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y99_SLICE_X99Y99_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y99_SLICE_X99Y99_AO6),
.Q(CLBLM_R_X65Y99_SLICE_X99Y99_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y99_SLICE_X99Y99_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y99_SLICE_X99Y99_BO6),
.Q(CLBLM_R_X65Y99_SLICE_X99Y99_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y99_SLICE_X99Y99_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y99_SLICE_X99Y99_CO6),
.Q(CLBLM_R_X65Y99_SLICE_X99Y99_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y99_SLICE_X99Y99_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y99_SLICE_X99Y99_DO6),
.Q(CLBLM_R_X65Y99_SLICE_X99Y99_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5eda1edaaaaaaaa)
  ) CLBLM_R_X65Y99_SLICE_X99Y99_DLUT (
.I0(CLBLM_R_X65Y99_SLICE_X99Y99_C5Q),
.I1(CLBLM_R_X65Y99_SLICE_X99Y99_CQ),
.I2(CLBLM_R_X65Y99_SLICE_X99Y99_DQ),
.I3(CLBLM_R_X65Y99_SLICE_X99Y99_BQ),
.I4(CLBLM_R_X65Y99_SLICE_X99Y99_AQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_R_X65Y99_SLICE_X99Y99_DO5),
.O6(CLBLM_R_X65Y99_SLICE_X99Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff005500444cc4cc)
  ) CLBLM_R_X65Y99_SLICE_X99Y99_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_R_X65Y99_SLICE_X99Y99_CQ),
.I2(CLBLM_R_X65Y99_SLICE_X99Y99_DQ),
.I3(CLBLM_R_X65Y99_SLICE_X99Y99_BQ),
.I4(CLBLM_R_X65Y99_SLICE_X99Y99_AQ),
.I5(1'b1),
.O5(CLBLM_R_X65Y99_SLICE_X99Y99_CO5),
.O6(CLBLM_R_X65Y99_SLICE_X99Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff77fff0f0f0f0)
  ) CLBLM_R_X65Y99_SLICE_X99Y99_BLUT (
.I0(CLBLM_R_X67Y100_SLICE_X100Y100_CQ),
.I1(CLBLM_R_X67Y103_SLICE_X100Y103_BQ),
.I2(CLBLM_R_X65Y99_SLICE_X99Y99_AQ),
.I3(CLBLM_R_X67Y99_SLICE_X100Y99_AQ),
.I4(CLBLM_R_X67Y99_SLICE_X100Y99_BQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_R_X65Y99_SLICE_X99Y99_BO5),
.O6(CLBLM_R_X65Y99_SLICE_X99Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaaaaff77aaaa)
  ) CLBLM_R_X65Y99_SLICE_X99Y99_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_R_X67Y100_SLICE_X100Y100_BQ),
.I2(1'b1),
.I3(CLBLM_R_X67Y99_SLICE_X100Y99_AQ),
.I4(CLBLM_R_X67Y99_SLICE_X100Y99_BQ),
.I5(CLBLM_R_X67Y100_SLICE_X100Y100_CQ),
.O5(CLBLM_R_X65Y99_SLICE_X99Y99_AO5),
.O6(CLBLM_R_X65Y99_SLICE_X99Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y100_SLICE_X98Y100_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y100_SLICE_X98Y100_AO6),
.Q(CLBLM_R_X65Y100_SLICE_X98Y100_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y100_SLICE_X98Y100_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y100_SLICE_X98Y100_BO6),
.Q(CLBLM_R_X65Y100_SLICE_X98Y100_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y100_SLICE_X98Y100_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y100_SLICE_X98Y100_DO5),
.O6(CLBLM_R_X65Y100_SLICE_X98Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y100_SLICE_X98Y100_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y100_SLICE_X98Y100_CO5),
.O6(CLBLM_R_X65Y100_SLICE_X98Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h72d8d8d8d8d8d8d8)
  ) CLBLM_R_X65Y100_SLICE_X98Y100_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_R_X65Y100_SLICE_X98Y100_BQ),
.I2(CLBLM_R_X65Y100_SLICE_X98Y100_AQ),
.I3(CLBLM_L_X64Y99_SLICE_X96Y99_A5Q),
.I4(CLBLM_R_X63Y99_SLICE_X94Y99_A5Q),
.I5(CLBLM_L_X64Y99_SLICE_X96Y99_BQ),
.O5(CLBLM_R_X65Y100_SLICE_X98Y100_BO5),
.O6(CLBLM_R_X65Y100_SLICE_X98Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h72cc72ccd8ccd8cc)
  ) CLBLM_R_X65Y100_SLICE_X98Y100_ALUT (
.I0(CLBLM_R_X63Y99_SLICE_X95Y99_AO5),
.I1(CLBLM_R_X65Y99_SLICE_X98Y99_AQ),
.I2(CLBLM_R_X65Y100_SLICE_X98Y100_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(1'b1),
.I5(CLBLM_R_X65Y99_SLICE_X98Y99_BQ),
.O5(CLBLM_R_X65Y100_SLICE_X98Y100_AO5),
.O6(CLBLM_R_X65Y100_SLICE_X98Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y100_SLICE_X99Y100_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y100_SLICE_X99Y100_AO5),
.Q(CLBLM_R_X65Y100_SLICE_X99Y100_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y100_SLICE_X99Y100_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y100_SLICE_X99Y100_AO6),
.Q(CLBLM_R_X65Y100_SLICE_X99Y100_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y100_SLICE_X99Y100_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y100_SLICE_X99Y100_BO6),
.Q(CLBLM_R_X65Y100_SLICE_X99Y100_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y100_SLICE_X99Y100_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y100_SLICE_X99Y100_CO6),
.Q(CLBLM_R_X65Y100_SLICE_X99Y100_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y100_SLICE_X99Y100_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y100_SLICE_X99Y100_DO5),
.O6(CLBLM_R_X65Y100_SLICE_X99Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hac5cff00ac5cff00)
  ) CLBLM_R_X65Y100_SLICE_X99Y100_CLUT (
.I0(CLBLM_R_X65Y101_SLICE_X99Y101_AQ),
.I1(CLBLM_R_X65Y100_SLICE_X99Y100_CQ),
.I2(CLBLM_L_X64Y99_SLICE_X96Y99_BO5),
.I3(CLBLM_R_X65Y100_SLICE_X99Y100_BQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLM_R_X65Y100_SLICE_X99Y100_CO5),
.O6(CLBLM_R_X65Y100_SLICE_X99Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf2fafafad0505050)
  ) CLBLM_R_X65Y100_SLICE_X99Y100_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X64Y99_SLICE_X96Y99_A5Q),
.I2(CLBLM_R_X65Y101_SLICE_X99Y101_AQ),
.I3(CLBLM_L_X64Y99_SLICE_X96Y99_BQ),
.I4(CLBLM_R_X63Y99_SLICE_X94Y99_A5Q),
.I5(CLBLM_R_X65Y100_SLICE_X99Y100_BQ),
.O5(CLBLM_R_X65Y100_SLICE_X99Y100_BO5),
.O6(CLBLM_R_X65Y100_SLICE_X99Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfb40fb40f47cb038)
  ) CLBLM_R_X65Y100_SLICE_X99Y100_ALUT (
.I0(CLBLM_R_X63Y99_SLICE_X95Y99_AO5),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_R_X65Y100_SLICE_X99Y100_AQ),
.I3(CLBLM_R_X65Y100_SLICE_X98Y100_BQ),
.I4(CLBLM_R_X65Y100_SLICE_X99Y100_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X65Y100_SLICE_X99Y100_AO5),
.O6(CLBLM_R_X65Y100_SLICE_X99Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y101_SLICE_X98Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y101_SLICE_X98Y101_DO5),
.O6(CLBLM_R_X65Y101_SLICE_X98Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y101_SLICE_X98Y101_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y101_SLICE_X98Y101_CO5),
.O6(CLBLM_R_X65Y101_SLICE_X98Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y101_SLICE_X98Y101_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y101_SLICE_X98Y101_BO5),
.O6(CLBLM_R_X65Y101_SLICE_X98Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y101_SLICE_X98Y101_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y101_SLICE_X98Y101_AO5),
.O6(CLBLM_R_X65Y101_SLICE_X98Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y101_SLICE_X99Y101_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y101_SLICE_X99Y101_AO5),
.Q(CLBLM_R_X65Y101_SLICE_X99Y101_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y101_SLICE_X99Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y101_SLICE_X99Y101_DO5),
.O6(CLBLM_R_X65Y101_SLICE_X99Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y101_SLICE_X99Y101_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y101_SLICE_X99Y101_CO5),
.O6(CLBLM_R_X65Y101_SLICE_X99Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y101_SLICE_X99Y101_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y101_SLICE_X99Y101_BO5),
.O6(CLBLM_R_X65Y101_SLICE_X99Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00aa003cff3c00)
  ) CLBLM_R_X65Y101_SLICE_X99Y101_ALUT (
.I0(CLBLM_R_X65Y100_SLICE_X99Y100_CQ),
.I1(CLBLM_R_X63Y99_SLICE_X95Y99_AO5),
.I2(CLBLM_R_X65Y101_SLICE_X99Y101_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_R_X65Y100_SLICE_X99Y100_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X65Y101_SLICE_X99Y101_AO5),
.O6(CLBLM_R_X65Y101_SLICE_X99Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y102_SLICE_X98Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y102_SLICE_X98Y102_DO5),
.O6(CLBLM_R_X65Y102_SLICE_X98Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y102_SLICE_X98Y102_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y102_SLICE_X98Y102_CO5),
.O6(CLBLM_R_X65Y102_SLICE_X98Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y102_SLICE_X98Y102_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y102_SLICE_X98Y102_BO5),
.O6(CLBLM_R_X65Y102_SLICE_X98Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y102_SLICE_X98Y102_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y102_SLICE_X98Y102_AO5),
.O6(CLBLM_R_X65Y102_SLICE_X98Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y102_SLICE_X99Y102_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y102_SLICE_X99Y102_AO6),
.Q(CLBLM_R_X65Y102_SLICE_X99Y102_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y102_SLICE_X99Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y102_SLICE_X99Y102_DO5),
.O6(CLBLM_R_X65Y102_SLICE_X99Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y102_SLICE_X99Y102_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y102_SLICE_X99Y102_CO5),
.O6(CLBLM_R_X65Y102_SLICE_X99Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y102_SLICE_X99Y102_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y102_SLICE_X99Y102_BO5),
.O6(CLBLM_R_X65Y102_SLICE_X99Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2020202020a02020)
  ) CLBLM_R_X65Y102_SLICE_X99Y102_ALUT (
.I0(CLBLM_L_X70Y101_SLICE_X104Y101_DO6),
.I1(CLBLM_R_X65Y103_SLICE_X99Y103_DO6),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_R_X65Y104_SLICE_X98Y104_C5Q),
.I4(CLBLM_R_X65Y104_SLICE_X99Y104_DO6),
.I5(CLBLM_R_X65Y104_SLICE_X98Y104_CQ),
.O5(CLBLM_R_X65Y102_SLICE_X99Y102_AO5),
.O6(CLBLM_R_X65Y102_SLICE_X99Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y103_SLICE_X98Y103_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y104_SLICE_X99Y104_B5Q),
.Q(CLBLM_R_X65Y103_SLICE_X98Y103_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y103_SLICE_X98Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y103_SLICE_X98Y103_AO6),
.Q(CLBLM_R_X65Y103_SLICE_X98Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y103_SLICE_X98Y103_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y103_SLICE_X98Y103_BO6),
.Q(CLBLM_R_X65Y103_SLICE_X98Y103_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888ff88ff88)
  ) CLBLM_R_X65Y103_SLICE_X98Y103_DLUT (
.I0(CLBLM_L_X64Y100_SLICE_X97Y100_AQ),
.I1(CLBLM_R_X65Y104_SLICE_X99Y104_B5Q),
.I2(1'b1),
.I3(CLBLM_R_X65Y103_SLICE_X98Y103_A5Q),
.I4(1'b1),
.I5(CLBLM_L_X64Y103_SLICE_X96Y103_AQ),
.O5(CLBLM_R_X65Y103_SLICE_X98Y103_DO5),
.O6(CLBLM_R_X65Y103_SLICE_X98Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1d1d00cc1d1d33ff)
  ) CLBLM_R_X65Y103_SLICE_X98Y103_CLUT (
.I0(CLBLM_R_X65Y103_SLICE_X99Y103_AQ),
.I1(CLBLM_R_X65Y104_SLICE_X98Y104_CQ),
.I2(CLBLM_L_X64Y103_SLICE_X97Y103_BQ),
.I3(CLBLM_L_X64Y103_SLICE_X97Y103_AQ),
.I4(CLBLM_R_X65Y104_SLICE_X98Y104_C5Q),
.I5(CLBLM_L_X64Y105_SLICE_X97Y105_AQ),
.O5(CLBLM_R_X65Y103_SLICE_X98Y103_CO5),
.O6(CLBLM_R_X65Y103_SLICE_X98Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h64ccf0f0ccccf0f0)
  ) CLBLM_R_X65Y103_SLICE_X98Y103_BLUT (
.I0(CLBLM_R_X65Y104_SLICE_X98Y104_B5Q),
.I1(CLBLM_R_X65Y103_SLICE_X98Y103_BQ),
.I2(CLBLM_R_X65Y103_SLICE_X98Y103_AQ),
.I3(CLBLM_R_X65Y104_SLICE_X98Y104_BQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_R_X65Y103_SLICE_X98Y103_A5Q),
.O5(CLBLM_R_X65Y103_SLICE_X98Y103_BO5),
.O6(CLBLM_R_X65Y103_SLICE_X98Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h52f0aaaaf0f0aaaa)
  ) CLBLM_R_X65Y103_SLICE_X98Y103_ALUT (
.I0(CLBLM_R_X65Y104_SLICE_X98Y104_B5Q),
.I1(CLBLM_R_X65Y103_SLICE_X98Y103_BQ),
.I2(CLBLM_R_X65Y103_SLICE_X98Y103_AQ),
.I3(CLBLM_R_X65Y104_SLICE_X98Y104_BQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_R_X65Y103_SLICE_X98Y103_A5Q),
.O5(CLBLM_R_X65Y103_SLICE_X98Y103_AO5),
.O6(CLBLM_R_X65Y103_SLICE_X98Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y103_SLICE_X99Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y103_SLICE_X99Y103_AO6),
.Q(CLBLM_R_X65Y103_SLICE_X99Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y103_SLICE_X99Y103_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y103_SLICE_X99Y103_BO6),
.Q(CLBLM_R_X65Y103_SLICE_X99Y103_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0f0f0f0f0f0f0f0)
  ) CLBLM_R_X65Y103_SLICE_X99Y103_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X65Y104_SLICE_X98Y104_CQ),
.I2(CLBLM_R_X65Y105_SLICE_X98Y105_B5Q),
.I3(CLBLM_R_X65Y103_SLICE_X99Y103_CO6),
.I4(CLBLM_R_X65Y103_SLICE_X99Y103_AQ),
.I5(CLBLM_R_X65Y104_SLICE_X98Y104_C5Q),
.O5(CLBLM_R_X65Y103_SLICE_X99Y103_DO5),
.O6(CLBLM_R_X65Y103_SLICE_X99Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0400000000000000)
  ) CLBLM_R_X65Y103_SLICE_X99Y103_CLUT (
.I0(CLBLM_R_X65Y103_SLICE_X99Y103_BQ),
.I1(CLBLM_R_X65Y104_SLICE_X99Y104_AQ),
.I2(CLBLM_R_X65Y104_SLICE_X99Y104_A5Q),
.I3(CLBLM_R_X65Y104_SLICE_X98Y104_B5Q),
.I4(CLBLM_R_X65Y104_SLICE_X98Y104_BQ),
.I5(CLBLM_R_X65Y103_SLICE_X98Y103_BQ),
.O5(CLBLM_R_X65Y103_SLICE_X99Y103_CO5),
.O6(CLBLM_R_X65Y103_SLICE_X99Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff800000000000)
  ) CLBLM_R_X65Y103_SLICE_X99Y103_BLUT (
.I0(CLBLM_R_X65Y104_SLICE_X98Y104_B5Q),
.I1(CLBLM_R_X65Y104_SLICE_X98Y104_BQ),
.I2(CLBLM_R_X65Y103_SLICE_X98Y103_A5Q),
.I3(CLBLM_R_X65Y103_SLICE_X98Y103_BQ),
.I4(CLBLM_R_X65Y103_SLICE_X99Y103_BQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_R_X65Y103_SLICE_X99Y103_BO5),
.O6(CLBLM_R_X65Y103_SLICE_X99Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a0f5fda020)
  ) CLBLM_R_X65Y103_SLICE_X99Y103_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_R_X65Y104_SLICE_X99Y104_DO6),
.I2(CLBLM_R_X65Y103_SLICE_X99Y103_AQ),
.I3(CLBLM_R_X65Y104_SLICE_X98Y104_C5Q),
.I4(CLBLM_R_X65Y102_SLICE_X99Y102_AQ),
.I5(CLBLM_R_X65Y104_SLICE_X98Y104_CQ),
.O5(CLBLM_R_X65Y103_SLICE_X99Y103_AO5),
.O6(CLBLM_R_X65Y103_SLICE_X99Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y104_SLICE_X98Y104_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y104_SLICE_X98Y104_BO5),
.Q(CLBLM_R_X65Y104_SLICE_X98Y104_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y104_SLICE_X98Y104_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y104_SLICE_X98Y104_CO5),
.Q(CLBLM_R_X65Y104_SLICE_X98Y104_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y104_SLICE_X98Y104_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y104_SLICE_X98Y104_BO6),
.Q(CLBLM_R_X65Y104_SLICE_X98Y104_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y104_SLICE_X98Y104_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y104_SLICE_X98Y104_CO6),
.Q(CLBLM_R_X65Y104_SLICE_X98Y104_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4ccccccccccccccc)
  ) CLBLM_R_X65Y104_SLICE_X98Y104_DLUT (
.I0(CLBLM_R_X65Y103_SLICE_X98Y103_BQ),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_R_X65Y104_SLICE_X98Y104_BQ),
.I3(CLBLM_R_X65Y103_SLICE_X98Y103_A5Q),
.I4(CLBLM_R_X65Y104_SLICE_X98Y104_B5Q),
.I5(CLBLM_R_X65Y103_SLICE_X99Y103_BQ),
.O5(CLBLM_R_X65Y104_SLICE_X98Y104_DO5),
.O6(CLBLM_R_X65Y104_SLICE_X98Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88887d88aa005af0)
  ) CLBLM_R_X65Y104_SLICE_X98Y104_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_R_X65Y104_SLICE_X98Y104_CQ),
.I2(CLBLM_R_X65Y104_SLICE_X99Y104_AQ),
.I3(CLBLM_R_X65Y104_SLICE_X98Y104_C5Q),
.I4(CLBLM_R_X65Y104_SLICE_X98Y104_DO6),
.I5(1'b1),
.O5(CLBLM_R_X65Y104_SLICE_X98Y104_CO5),
.O6(CLBLM_R_X65Y104_SLICE_X98Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3cf0f06a6acccc)
  ) CLBLM_R_X65Y104_SLICE_X98Y104_BLUT (
.I0(CLBLM_R_X65Y104_SLICE_X98Y104_B5Q),
.I1(CLBLM_R_X65Y104_SLICE_X98Y104_BQ),
.I2(CLBLM_R_X65Y103_SLICE_X98Y103_A5Q),
.I3(1'b1),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLM_R_X65Y104_SLICE_X98Y104_BO5),
.O6(CLBLM_R_X65Y104_SLICE_X98Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8080000080000000)
  ) CLBLM_R_X65Y104_SLICE_X98Y104_ALUT (
.I0(CLBLM_R_X65Y104_SLICE_X98Y104_B5Q),
.I1(CLBLM_R_X65Y104_SLICE_X98Y104_BQ),
.I2(CLBLM_R_X65Y103_SLICE_X98Y103_A5Q),
.I3(CLBLM_R_X65Y103_SLICE_X99Y103_BQ),
.I4(CLBLM_R_X65Y103_SLICE_X98Y103_BQ),
.I5(1'b1),
.O5(CLBLM_R_X65Y104_SLICE_X98Y104_AO5),
.O6(CLBLM_R_X65Y104_SLICE_X98Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y104_SLICE_X99Y104_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y104_SLICE_X99Y104_AO5),
.Q(CLBLM_R_X65Y104_SLICE_X99Y104_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y104_SLICE_X99Y104_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y105_SLICE_X98Y105_B5Q),
.Q(CLBLM_R_X65Y104_SLICE_X99Y104_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y104_SLICE_X99Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y104_SLICE_X99Y104_AO6),
.Q(CLBLM_R_X65Y104_SLICE_X99Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y104_SLICE_X99Y104_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y104_SLICE_X99Y104_BO6),
.Q(CLBLM_R_X65Y104_SLICE_X99Y104_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff000000000000)
  ) CLBLM_R_X65Y104_SLICE_X99Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X65Y104_SLICE_X99Y104_A5Q),
.I4(CLBLM_R_X65Y104_SLICE_X99Y104_AQ),
.I5(CLBLM_R_X65Y103_SLICE_X99Y103_BQ),
.O5(CLBLM_R_X65Y104_SLICE_X99Y104_DO5),
.O6(CLBLM_R_X65Y104_SLICE_X99Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0f0fafaaabb)
  ) CLBLM_R_X65Y104_SLICE_X99Y104_CLUT (
.I0(CLBLM_R_X65Y104_SLICE_X99Y104_A5Q),
.I1(CLBLM_R_X65Y104_SLICE_X98Y104_C5Q),
.I2(CLBLM_R_X65Y103_SLICE_X98Y103_CO6),
.I3(CLBLM_R_X65Y104_SLICE_X98Y104_CQ),
.I4(CLBLM_R_X65Y104_SLICE_X99Y104_AQ),
.I5(CLBLM_R_X65Y103_SLICE_X99Y103_BQ),
.O5(CLBLM_R_X65Y104_SLICE_X99Y104_CO5),
.O6(CLBLM_R_X65Y104_SLICE_X99Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf00fff00ccccff00)
  ) CLBLM_R_X65Y104_SLICE_X99Y104_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X65Y104_SLICE_X99Y104_BQ),
.I2(CLBLM_R_X65Y105_SLICE_X99Y105_C5Q),
.I3(CLBLM_L_X64Y104_SLICE_X97Y104_AQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_R_X63Y103_SLICE_X95Y103_BO5),
.O5(CLBLM_R_X65Y104_SLICE_X99Y104_BO5),
.O6(CLBLM_R_X65Y104_SLICE_X99Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5faf00a00cfc5c0c)
  ) CLBLM_R_X65Y104_SLICE_X99Y104_ALUT (
.I0(CLBLM_R_X65Y104_SLICE_X99Y104_AQ),
.I1(CLBLM_R_X65Y103_SLICE_X99Y103_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_R_X65Y104_SLICE_X98Y104_AO5),
.I4(CLBLM_R_X65Y104_SLICE_X99Y104_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X65Y104_SLICE_X99Y104_AO5),
.O6(CLBLM_R_X65Y104_SLICE_X99Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y105_SLICE_X98Y105_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y105_SLICE_X98Y105_AQ),
.Q(CLBLM_R_X65Y105_SLICE_X98Y105_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y105_SLICE_X98Y105_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y105_SLICE_X98Y105_AO5),
.Q(CLBLM_R_X65Y105_SLICE_X98Y105_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y105_SLICE_X98Y105_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y105_SLICE_X98Y105_BO6),
.Q(CLBLM_R_X65Y105_SLICE_X98Y105_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y105_SLICE_X98Y105_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y105_SLICE_X98Y105_CO6),
.Q(CLBLM_R_X65Y105_SLICE_X98Y105_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff5fff0f5f5f0f0)
  ) CLBLM_R_X65Y105_SLICE_X98Y105_DLUT (
.I0(CLBLM_L_X70Y103_SLICE_X104Y103_AQ),
.I1(1'b1),
.I2(CLBLM_R_X65Y103_SLICE_X98Y103_DO6),
.I3(CLBLM_R_X65Y105_SLICE_X98Y105_AQ),
.I4(CLBLM_R_X65Y105_SLICE_X98Y105_B5Q),
.I5(CLBLM_R_X63Y106_SLICE_X95Y106_AQ),
.O5(CLBLM_R_X65Y105_SLICE_X98Y105_DO5),
.O6(CLBLM_R_X65Y105_SLICE_X98Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hba7aba7a8a4a8a4a)
  ) CLBLM_R_X65Y105_SLICE_X98Y105_CLUT (
.I0(CLBLM_R_X65Y105_SLICE_X98Y105_BQ),
.I1(CLBLM_L_X64Y106_SLICE_X97Y106_AO6),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_R_X65Y105_SLICE_X99Y105_AQ),
.I4(1'b1),
.I5(CLBLM_R_X65Y105_SLICE_X98Y105_CQ),
.O5(CLBLM_R_X65Y105_SLICE_X98Y105_CO5),
.O6(CLBLM_R_X65Y105_SLICE_X98Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hefcf40c0cfcfc0c0)
  ) CLBLM_R_X65Y105_SLICE_X98Y105_BLUT (
.I0(CLBLM_L_X64Y106_SLICE_X97Y106_B5Q),
.I1(CLBLM_R_X65Y105_SLICE_X98Y105_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X64Y106_SLICE_X97Y106_C5Q),
.I4(CLBLM_R_X65Y105_SLICE_X99Y105_AQ),
.I5(CLBLM_L_X64Y106_SLICE_X97Y106_AQ),
.O5(CLBLM_R_X65Y105_SLICE_X98Y105_BO5),
.O6(CLBLM_R_X65Y105_SLICE_X98Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0005000500010000)
  ) CLBLM_R_X65Y105_SLICE_X98Y105_ALUT (
.I0(CLBLM_R_X65Y105_SLICE_X98Y105_B5Q),
.I1(CLBLM_R_X65Y104_SLICE_X98Y104_AO6),
.I2(CLBLM_R_X65Y105_SLICE_X98Y105_AQ),
.I3(CLBLM_R_X65Y104_SLICE_X99Y104_B5Q),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLM_R_X65Y105_SLICE_X98Y105_AO5),
.O6(CLBLM_R_X65Y105_SLICE_X98Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y105_SLICE_X99Y105_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y105_SLICE_X99Y105_CO5),
.Q(CLBLM_R_X65Y105_SLICE_X99Y105_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y105_SLICE_X99Y105_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y105_SLICE_X99Y105_DO5),
.Q(CLBLM_R_X65Y105_SLICE_X99Y105_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y105_SLICE_X99Y105_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y105_SLICE_X99Y105_AO5),
.Q(CLBLM_R_X65Y105_SLICE_X99Y105_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y105_SLICE_X99Y105_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y105_SLICE_X99Y105_CO6),
.Q(CLBLM_R_X65Y105_SLICE_X99Y105_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y105_SLICE_X99Y105_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y105_SLICE_X99Y105_DO6),
.Q(CLBLM_R_X65Y105_SLICE_X99Y105_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaae2e2b4b4fc30)
  ) CLBLM_R_X65Y105_SLICE_X99Y105_DLUT (
.I0(CLBLM_L_X64Y105_SLICE_X97Y105_CQ),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_R_X65Y105_SLICE_X99Y105_DQ),
.I3(CLBLM_R_X65Y105_SLICE_X99Y105_D5Q),
.I4(CLBLM_R_X63Y101_SLICE_X94Y101_BO5),
.I5(1'b1),
.O5(CLBLM_R_X65Y105_SLICE_X99Y105_DO5),
.O6(CLBLM_R_X65Y105_SLICE_X99Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h330033007474b8b8)
  ) CLBLM_R_X65Y105_SLICE_X99Y105_CLUT (
.I0(CLBLM_R_X65Y105_SLICE_X99Y105_C5Q),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_R_X65Y105_SLICE_X99Y105_D5Q),
.I3(CLBLM_L_X72Y118_SLICE_X108Y118_CQ),
.I4(CLBLM_R_X63Y101_SLICE_X94Y101_BO5),
.I5(1'b1),
.O5(CLBLM_R_X65Y105_SLICE_X99Y105_CO5),
.O6(CLBLM_R_X65Y105_SLICE_X99Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff00000fffe0000)
  ) CLBLM_R_X65Y105_SLICE_X99Y105_BLUT (
.I0(CLBLM_R_X65Y100_SLICE_X99Y100_A5Q),
.I1(CLBLM_R_X65Y100_SLICE_X99Y100_CQ),
.I2(CLBLM_R_X65Y104_SLICE_X99Y104_BQ),
.I3(CLBLM_R_X65Y105_SLICE_X99Y105_D5Q),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLM_R_X65Y105_SLICE_X99Y105_BO5),
.O6(CLBLM_R_X65Y105_SLICE_X99Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00cc005acc5acc)
  ) CLBLM_R_X65Y105_SLICE_X99Y105_ALUT (
.I0(CLBLM_R_X63Y106_SLICE_X94Y106_AO6),
.I1(CLBLM_R_X65Y106_SLICE_X99Y106_C5Q),
.I2(CLBLM_R_X65Y105_SLICE_X99Y105_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_R_X65Y105_SLICE_X98Y105_CQ),
.I5(1'b1),
.O5(CLBLM_R_X65Y105_SLICE_X99Y105_AO5),
.O6(CLBLM_R_X65Y105_SLICE_X99Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y106_SLICE_X98Y106_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y106_SLICE_X98Y106_AO6),
.Q(CLBLM_R_X65Y106_SLICE_X98Y106_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y106_SLICE_X98Y106_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y106_SLICE_X98Y106_BO6),
.Q(CLBLM_R_X65Y106_SLICE_X98Y106_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y106_SLICE_X98Y106_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y106_SLICE_X98Y106_CO6),
.Q(CLBLM_R_X65Y106_SLICE_X98Y106_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y106_SLICE_X98Y106_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y106_SLICE_X98Y106_DO6),
.Q(CLBLM_R_X65Y106_SLICE_X98Y106_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h20a08a0aa0a00a0a)
  ) CLBLM_R_X65Y106_SLICE_X98Y106_DLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X64Y106_SLICE_X97Y106_AQ),
.I2(CLBLM_R_X65Y106_SLICE_X98Y106_DQ),
.I3(CLBLM_L_X64Y106_SLICE_X97Y106_B5Q),
.I4(CLBLL_R_X79Y99_SLICE_X122Y99_AO6),
.I5(CLBLM_L_X64Y106_SLICE_X97Y106_C5Q),
.O5(CLBLM_R_X65Y106_SLICE_X98Y106_DO5),
.O6(CLBLM_R_X65Y106_SLICE_X98Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4ee44ee4f0f0f0f0)
  ) CLBLM_R_X65Y106_SLICE_X98Y106_CLUT (
.I0(CLBLM_R_X63Y106_SLICE_X94Y106_AO6),
.I1(CLBLM_R_X65Y106_SLICE_X98Y106_CQ),
.I2(CLBLM_R_X65Y106_SLICE_X98Y106_AQ),
.I3(CLBLM_R_X65Y106_SLICE_X98Y106_BQ),
.I4(1'b1),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_R_X65Y106_SLICE_X98Y106_CO5),
.O6(CLBLM_R_X65Y106_SLICE_X98Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hefcf40c0cfcfc0c0)
  ) CLBLM_R_X65Y106_SLICE_X98Y106_BLUT (
.I0(CLBLM_L_X64Y106_SLICE_X97Y106_AQ),
.I1(CLBLM_R_X65Y106_SLICE_X98Y106_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X64Y106_SLICE_X97Y106_B5Q),
.I4(CLBLM_R_X65Y106_SLICE_X98Y106_DQ),
.I5(CLBLM_L_X64Y106_SLICE_X97Y106_C5Q),
.O5(CLBLM_R_X65Y106_SLICE_X98Y106_BO5),
.O6(CLBLM_R_X65Y106_SLICE_X98Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc0fcc00ccf0cc)
  ) CLBLM_R_X65Y106_SLICE_X98Y106_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X65Y106_SLICE_X98Y106_BQ),
.I2(CLBLM_R_X65Y106_SLICE_X98Y106_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_R_X63Y106_SLICE_X94Y106_AO6),
.I5(CLBLM_L_X62Y106_SLICE_X93Y106_DO6),
.O5(CLBLM_R_X65Y106_SLICE_X98Y106_AO5),
.O6(CLBLM_R_X65Y106_SLICE_X98Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y106_SLICE_X99Y106_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y106_SLICE_X99Y106_CO5),
.Q(CLBLM_R_X65Y106_SLICE_X99Y106_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y106_SLICE_X99Y106_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y106_SLICE_X99Y106_AO6),
.Q(CLBLM_R_X65Y106_SLICE_X99Y106_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y106_SLICE_X99Y106_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y106_SLICE_X99Y106_BO6),
.Q(CLBLM_R_X65Y106_SLICE_X99Y106_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y106_SLICE_X99Y106_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y106_SLICE_X99Y106_CO6),
.Q(CLBLM_R_X65Y106_SLICE_X99Y106_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y106_SLICE_X99Y106_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y106_SLICE_X99Y106_DO6),
.Q(CLBLM_R_X65Y106_SLICE_X99Y106_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a2a0a2a0a0a0a0)
  ) CLBLM_R_X65Y106_SLICE_X99Y106_DLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_R_X65Y104_SLICE_X99Y104_CO6),
.I2(CLBLM_R_X65Y105_SLICE_X98Y105_DO6),
.I3(CLBLM_R_X65Y103_SLICE_X98Y103_A5Q),
.I4(1'b1),
.I5(CLBLM_R_X65Y105_SLICE_X98Y105_AO6),
.O5(CLBLM_R_X65Y106_SLICE_X99Y106_DO5),
.O6(CLBLM_R_X65Y106_SLICE_X99Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0f0c3aacccc)
  ) CLBLM_R_X65Y106_SLICE_X99Y106_CLUT (
.I0(CLBLM_R_X65Y106_SLICE_X99Y106_C5Q),
.I1(CLBLM_R_X65Y106_SLICE_X99Y106_CQ),
.I2(CLBLM_R_X65Y106_SLICE_X99Y106_BQ),
.I3(CLBLM_R_X63Y106_SLICE_X94Y106_AO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLM_R_X65Y106_SLICE_X99Y106_CO5),
.O6(CLBLM_R_X65Y106_SLICE_X99Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6cccffff6ccc0000)
  ) CLBLM_R_X65Y106_SLICE_X99Y106_BLUT (
.I0(CLBLM_L_X64Y106_SLICE_X97Y106_AQ),
.I1(CLBLM_R_X65Y106_SLICE_X99Y106_BQ),
.I2(CLBLM_L_X64Y106_SLICE_X97Y106_B5Q),
.I3(CLBLM_L_X64Y106_SLICE_X97Y106_C5Q),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_R_X65Y106_SLICE_X98Y106_CQ),
.O5(CLBLM_R_X65Y106_SLICE_X99Y106_BO5),
.O6(CLBLM_R_X65Y106_SLICE_X99Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafa0a0bfafb0a0)
  ) CLBLM_R_X65Y106_SLICE_X99Y106_ALUT (
.I0(CLBLM_R_X65Y105_SLICE_X98Y105_DO6),
.I1(CLBLM_R_X65Y103_SLICE_X98Y103_A5Q),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_R_X65Y105_SLICE_X98Y105_AO6),
.I4(CLBLM_R_X65Y106_SLICE_X99Y106_DQ),
.I5(CLBLM_R_X65Y104_SLICE_X99Y104_CO6),
.O5(CLBLM_R_X65Y106_SLICE_X99Y106_AO5),
.O6(CLBLM_R_X65Y106_SLICE_X99Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y108_SLICE_X98Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y108_SLICE_X98Y108_DO5),
.O6(CLBLM_R_X65Y108_SLICE_X98Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y108_SLICE_X98Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y108_SLICE_X98Y108_CO5),
.O6(CLBLM_R_X65Y108_SLICE_X98Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cc008000800080)
  ) CLBLM_R_X65Y108_SLICE_X98Y108_BLUT (
.I0(CLBLM_R_X65Y109_SLICE_X99Y109_CQ),
.I1(CLBLM_L_X68Y108_SLICE_X102Y108_A5Q),
.I2(CLBLM_R_X65Y109_SLICE_X98Y109_A5Q),
.I3(CLBLM_L_X68Y108_SLICE_X102Y108_AQ),
.I4(CLBLM_L_X62Y92_SLICE_X92Y92_BQ),
.I5(CLBLM_R_X65Y110_SLICE_X98Y110_AQ),
.O5(CLBLM_R_X65Y108_SLICE_X98Y108_BO5),
.O6(CLBLM_R_X65Y108_SLICE_X98Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc8880000c0000000)
  ) CLBLM_R_X65Y108_SLICE_X98Y108_ALUT (
.I0(CLBLM_R_X65Y110_SLICE_X98Y110_A5Q),
.I1(CLBLM_L_X68Y108_SLICE_X102Y108_A5Q),
.I2(CLBLM_R_X65Y111_SLICE_X98Y111_AQ),
.I3(CLBLM_R_X65Y110_SLICE_X98Y110_BQ),
.I4(CLBLM_L_X68Y108_SLICE_X102Y108_AQ),
.I5(CLBLM_R_X65Y109_SLICE_X98Y109_CQ),
.O5(CLBLM_R_X65Y108_SLICE_X98Y108_AO5),
.O6(CLBLM_R_X65Y108_SLICE_X98Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y108_SLICE_X99Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y108_SLICE_X99Y108_DO5),
.O6(CLBLM_R_X65Y108_SLICE_X99Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0020ffff0020)
  ) CLBLM_R_X65Y108_SLICE_X99Y108_CLUT (
.I0(CLBLM_R_X65Y110_SLICE_X99Y110_CQ),
.I1(CLBLM_L_X68Y108_SLICE_X102Y108_AQ),
.I2(CLBLM_R_X65Y109_SLICE_X99Y109_BQ),
.I3(CLBLM_L_X68Y108_SLICE_X102Y108_A5Q),
.I4(CLBLM_L_X68Y109_SLICE_X102Y109_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X65Y108_SLICE_X99Y108_CO5),
.O6(CLBLM_R_X65Y108_SLICE_X99Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8a800a0080800000)
  ) CLBLM_R_X65Y108_SLICE_X99Y108_BLUT (
.I0(CLBLM_L_X68Y108_SLICE_X102Y108_A5Q),
.I1(CLBLM_R_X65Y109_SLICE_X98Y109_A5Q),
.I2(CLBLM_L_X68Y108_SLICE_X102Y108_AQ),
.I3(CLBLM_R_X65Y110_SLICE_X99Y110_BQ),
.I4(CLBLM_R_X67Y109_SLICE_X101Y109_BQ),
.I5(CLBLM_R_X65Y110_SLICE_X98Y110_A5Q),
.O5(CLBLM_R_X65Y108_SLICE_X99Y108_BO5),
.O6(CLBLM_R_X65Y108_SLICE_X99Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffdfdff00fd00)
  ) CLBLM_R_X65Y108_SLICE_X99Y108_ALUT (
.I0(CLBLM_R_X65Y109_SLICE_X98Y109_DO6),
.I1(CLBLM_R_X65Y108_SLICE_X98Y108_BO6),
.I2(CLBLM_R_X65Y108_SLICE_X98Y108_AO6),
.I3(CLBLM_R_X65Y108_SLICE_X99Y108_BO6),
.I4(CLBLM_R_X65Y108_SLICE_X99Y108_CO6),
.I5(CLBLM_R_X65Y109_SLICE_X99Y109_DO5),
.O5(CLBLM_R_X65Y108_SLICE_X99Y108_AO5),
.O6(CLBLM_R_X65Y108_SLICE_X99Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y109_SLICE_X98Y109_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y110_SLICE_X99Y110_CQ),
.Q(CLBLM_R_X65Y109_SLICE_X98Y109_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y109_SLICE_X98Y109_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y109_SLICE_X98Y109_AO6),
.Q(CLBLM_R_X65Y109_SLICE_X98Y109_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y109_SLICE_X98Y109_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y109_SLICE_X98Y109_BO6),
.Q(CLBLM_R_X65Y109_SLICE_X98Y109_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y109_SLICE_X98Y109_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y109_SLICE_X98Y109_CO6),
.Q(CLBLM_R_X65Y109_SLICE_X98Y109_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff57775fff)
  ) CLBLM_R_X65Y109_SLICE_X98Y109_DLUT (
.I0(CLBLM_L_X68Y108_SLICE_X102Y108_AQ),
.I1(CLBLM_R_X65Y109_SLICE_X99Y109_A5Q),
.I2(CLBLM_R_X65Y109_SLICE_X98Y109_AQ),
.I3(CLBLM_R_X65Y110_SLICE_X99Y110_AQ),
.I4(CLBLM_R_X65Y109_SLICE_X98Y109_BQ),
.I5(CLBLM_L_X68Y108_SLICE_X102Y108_A5Q),
.O5(CLBLM_R_X65Y109_SLICE_X98Y109_DO5),
.O6(CLBLM_R_X65Y109_SLICE_X98Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffd8ffcc00d800)
  ) CLBLM_R_X65Y109_SLICE_X98Y109_CLUT (
.I0(CLBLM_R_X65Y111_SLICE_X99Y111_AO6),
.I1(CLBLM_R_X65Y109_SLICE_X98Y109_CQ),
.I2(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_R_X67Y111_SLICE_X101Y111_CO5),
.I5(CLBLM_R_X65Y109_SLICE_X98Y109_AQ),
.O5(CLBLM_R_X65Y109_SLICE_X98Y109_CO5),
.O6(CLBLM_R_X65Y109_SLICE_X98Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffacffcc00ac00)
  ) CLBLM_R_X65Y109_SLICE_X98Y109_BLUT (
.I0(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I1(CLBLM_R_X65Y109_SLICE_X98Y109_BQ),
.I2(CLBLM_R_X67Y111_SLICE_X101Y111_B5Q),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_R_X65Y111_SLICE_X99Y111_AO6),
.I5(CLBLM_R_X65Y109_SLICE_X99Y109_CQ),
.O5(CLBLM_R_X65Y109_SLICE_X98Y109_BO5),
.O6(CLBLM_R_X65Y109_SLICE_X98Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000e2ffe200)
  ) CLBLM_R_X65Y109_SLICE_X98Y109_ALUT (
.I0(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I1(CLBLM_R_X65Y111_SLICE_X99Y111_AO6),
.I2(CLBLM_R_X65Y109_SLICE_X98Y109_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_R_X65Y110_SLICE_X98Y110_AQ),
.I5(CLBLM_R_X67Y111_SLICE_X101Y111_CO6),
.O5(CLBLM_R_X65Y109_SLICE_X98Y109_AO5),
.O6(CLBLM_R_X65Y109_SLICE_X98Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y109_SLICE_X99Y109_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y109_SLICE_X98Y109_A5Q),
.Q(CLBLM_R_X65Y109_SLICE_X99Y109_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y109_SLICE_X99Y109_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y109_SLICE_X99Y109_AO6),
.Q(CLBLM_R_X65Y109_SLICE_X99Y109_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y109_SLICE_X99Y109_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y109_SLICE_X99Y109_BO6),
.Q(CLBLM_R_X65Y109_SLICE_X99Y109_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y109_SLICE_X99Y109_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y109_SLICE_X99Y109_CO6),
.Q(CLBLM_R_X65Y109_SLICE_X99Y109_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0505050537333333)
  ) CLBLM_R_X65Y109_SLICE_X99Y109_DLUT (
.I0(CLBLM_L_X68Y108_SLICE_X102Y108_AQ),
.I1(CLBLM_L_X68Y109_SLICE_X102Y109_A5Q),
.I2(CLBLM_L_X68Y108_SLICE_X102Y108_A5Q),
.I3(CLBLM_R_X65Y109_SLICE_X99Y109_AQ),
.I4(CLBLM_R_X65Y110_SLICE_X99Y110_AQ),
.I5(1'b1),
.O5(CLBLM_R_X65Y109_SLICE_X99Y109_DO5),
.O6(CLBLM_R_X65Y109_SLICE_X99Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcdffc8ffcd00c800)
  ) CLBLM_R_X65Y109_SLICE_X99Y109_CLUT (
.I0(CLBLM_R_X65Y111_SLICE_X99Y111_AO6),
.I1(CLBLM_R_X65Y109_SLICE_X99Y109_CQ),
.I2(CLBLM_R_X67Y111_SLICE_X101Y111_DO5),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I5(CLBLM_R_X65Y109_SLICE_X99Y109_BQ),
.O5(CLBLM_R_X65Y109_SLICE_X99Y109_CO5),
.O6(CLBLM_R_X65Y109_SLICE_X99Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffd8ffcc00d800)
  ) CLBLM_R_X65Y109_SLICE_X99Y109_BLUT (
.I0(CLBLM_R_X67Y111_SLICE_X101Y111_DO6),
.I1(CLBLM_R_X65Y109_SLICE_X99Y109_BQ),
.I2(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_R_X65Y111_SLICE_X99Y111_AO6),
.I5(CLBLM_R_X65Y109_SLICE_X98Y109_CQ),
.O5(CLBLM_R_X65Y109_SLICE_X99Y109_BO5),
.O6(CLBLM_R_X65Y109_SLICE_X99Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaab8ff00ff00)
  ) CLBLM_R_X65Y109_SLICE_X99Y109_ALUT (
.I0(CLBLM_R_X65Y109_SLICE_X99Y109_AQ),
.I1(CLBLM_R_X67Y111_SLICE_X101Y111_CO6),
.I2(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I3(CLBLM_R_X67Y111_SLICE_X100Y111_A5Q),
.I4(CLBLM_R_X67Y111_SLICE_X101Y111_A5Q),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_R_X65Y109_SLICE_X99Y109_AO5),
.O6(CLBLM_R_X65Y109_SLICE_X99Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y110_SLICE_X98Y110_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y110_SLICE_X99Y110_AQ),
.Q(CLBLM_R_X65Y110_SLICE_X98Y110_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y110_SLICE_X98Y110_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y110_SLICE_X98Y110_AO6),
.Q(CLBLM_R_X65Y110_SLICE_X98Y110_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y110_SLICE_X98Y110_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y110_SLICE_X98Y110_BO6),
.Q(CLBLM_R_X65Y110_SLICE_X98Y110_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y110_SLICE_X98Y110_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y110_SLICE_X98Y110_CO6),
.Q(CLBLM_R_X65Y110_SLICE_X98Y110_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y110_SLICE_X98Y110_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y110_SLICE_X98Y110_DO6),
.Q(CLBLM_R_X65Y110_SLICE_X98Y110_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0ccf0ccaacc)
  ) CLBLM_R_X65Y110_SLICE_X98Y110_DLUT (
.I0(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I1(CLBLM_R_X65Y110_SLICE_X98Y110_CQ),
.I2(CLBLM_R_X65Y110_SLICE_X98Y110_DQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_R_X65Y111_SLICE_X99Y111_AO5),
.I5(CLBLM_R_X67Y111_SLICE_X101Y111_DO6),
.O5(CLBLM_R_X65Y110_SLICE_X98Y110_DO5),
.O6(CLBLM_R_X65Y110_SLICE_X98Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaacfaaccaac0aa)
  ) CLBLM_R_X65Y110_SLICE_X98Y110_CLUT (
.I0(CLBLM_R_X65Y110_SLICE_X98Y110_BQ),
.I1(CLBLM_R_X65Y110_SLICE_X98Y110_CQ),
.I2(CLBLM_R_X67Y111_SLICE_X101Y111_CO5),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_R_X65Y111_SLICE_X99Y111_AO5),
.I5(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.O5(CLBLM_R_X65Y110_SLICE_X98Y110_CO5),
.O6(CLBLM_R_X65Y110_SLICE_X98Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcdc8cdc8ffff0000)
  ) CLBLM_R_X65Y110_SLICE_X98Y110_BLUT (
.I0(CLBLM_R_X65Y111_SLICE_X99Y111_AO5),
.I1(CLBLM_R_X65Y110_SLICE_X98Y110_BQ),
.I2(CLBLM_R_X67Y111_SLICE_X101Y111_CO6),
.I3(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I4(CLBLM_R_X65Y109_SLICE_X98Y109_BQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_R_X65Y110_SLICE_X98Y110_BO5),
.O6(CLBLM_R_X65Y110_SLICE_X98Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2e2e2ee22e2e2)
  ) CLBLM_R_X65Y110_SLICE_X98Y110_ALUT (
.I0(CLBLM_R_X67Y110_SLICE_X100Y110_BQ),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_R_X65Y110_SLICE_X98Y110_AQ),
.I3(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I4(CLBLM_R_X67Y111_SLICE_X101Y111_B5Q),
.I5(CLBLM_R_X65Y110_SLICE_X99Y110_AO6),
.O5(CLBLM_R_X65Y110_SLICE_X98Y110_AO5),
.O6(CLBLM_R_X65Y110_SLICE_X98Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y110_SLICE_X99Y110_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X76Y111_SLICE_X116Y111_AQ),
.Q(CLBLM_R_X65Y110_SLICE_X99Y110_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y110_SLICE_X99Y110_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_L_X62Y92_SLICE_X92Y92_BQ),
.Q(CLBLM_R_X65Y110_SLICE_X99Y110_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y110_SLICE_X99Y110_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y110_SLICE_X99Y110_BO6),
.Q(CLBLM_R_X65Y110_SLICE_X99Y110_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y110_SLICE_X99Y110_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y110_SLICE_X98Y110_A5Q),
.Q(CLBLM_R_X65Y110_SLICE_X99Y110_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3300000000000000)
  ) CLBLM_R_X65Y110_SLICE_X99Y110_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X68Y108_SLICE_X102Y108_AQ),
.I2(1'b1),
.I3(CLBLM_L_X68Y108_SLICE_X102Y108_A5Q),
.I4(CLBLM_R_X65Y110_SLICE_X98Y110_DQ),
.I5(CLBLM_R_X65Y110_SLICE_X99Y110_B5Q),
.O5(CLBLM_R_X65Y110_SLICE_X99Y110_DO5),
.O6(CLBLM_R_X65Y110_SLICE_X99Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffc000aaaaaaaa)
  ) CLBLM_R_X65Y110_SLICE_X99Y110_CLUT (
.I0(CLBLM_R_X67Y110_SLICE_X100Y110_DO6),
.I1(CLBLM_L_X76Y111_SLICE_X116Y111_AQ),
.I2(CLBLM_R_X65Y109_SLICE_X99Y109_DO6),
.I3(CLBLM_R_X65Y110_SLICE_X98Y110_CQ),
.I4(CLBLM_R_X65Y110_SLICE_X99Y110_DO6),
.I5(CLBLM_R_X67Y109_SLICE_X100Y109_DO6),
.O5(CLBLM_R_X65Y110_SLICE_X99Y110_CO5),
.O6(CLBLM_R_X65Y110_SLICE_X99Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0f0dd88f0f0)
  ) CLBLM_R_X65Y110_SLICE_X99Y110_BLUT (
.I0(CLBLM_R_X67Y111_SLICE_X101Y111_CO5),
.I1(CLBLM_R_X65Y110_SLICE_X99Y110_BQ),
.I2(CLBLM_R_X65Y109_SLICE_X99Y109_AQ),
.I3(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_R_X65Y110_SLICE_X99Y110_AO5),
.O5(CLBLM_R_X65Y110_SLICE_X99Y110_BO5),
.O6(CLBLM_R_X65Y110_SLICE_X99Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddddddeeeeeeee)
  ) CLBLM_R_X65Y110_SLICE_X99Y110_ALUT (
.I0(CLBLM_R_X67Y111_SLICE_X101Y111_A5Q),
.I1(CLBLM_R_X67Y111_SLICE_X100Y111_A5Q),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y110_SLICE_X99Y110_AO5),
.O6(CLBLM_R_X65Y110_SLICE_X99Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X65Y111_SLICE_X98Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X65Y111_SLICE_X98Y111_AO6),
.Q(CLBLM_R_X65Y111_SLICE_X98Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y111_SLICE_X98Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y111_SLICE_X98Y111_DO5),
.O6(CLBLM_R_X65Y111_SLICE_X98Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y111_SLICE_X98Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y111_SLICE_X98Y111_CO5),
.O6(CLBLM_R_X65Y111_SLICE_X98Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0004000f3005100)
  ) CLBLM_R_X65Y111_SLICE_X98Y111_BLUT (
.I0(CLBLM_R_X65Y110_SLICE_X99Y110_AQ),
.I1(CLBLM_L_X76Y111_SLICE_X116Y111_AQ),
.I2(CLBLM_R_X65Y111_SLICE_X98Y111_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_L_X62Y92_SLICE_X92Y92_BQ),
.I5(CLBLM_R_X65Y110_SLICE_X99Y110_B5Q),
.O5(CLBLM_R_X65Y111_SLICE_X98Y111_BO5),
.O6(CLBLM_R_X65Y111_SLICE_X98Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2a007f0000005500)
  ) CLBLM_R_X65Y111_SLICE_X98Y111_ALUT (
.I0(CLBLM_L_X60Y97_SLICE_X91Y97_AQ),
.I1(CLBLM_L_X76Y111_SLICE_X116Y111_AQ),
.I2(CLBLM_R_X65Y111_SLICE_X98Y111_AQ),
.I3(CLBLM_R_X65Y111_SLICE_X98Y111_BO6),
.I4(CLBLM_L_X62Y92_SLICE_X92Y92_BQ),
.I5(CLBLM_R_X65Y110_SLICE_X99Y110_B5Q),
.O5(CLBLM_R_X65Y111_SLICE_X98Y111_AO5),
.O6(CLBLM_R_X65Y111_SLICE_X98Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y111_SLICE_X99Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y111_SLICE_X99Y111_DO5),
.O6(CLBLM_R_X65Y111_SLICE_X99Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y111_SLICE_X99Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y111_SLICE_X99Y111_CO5),
.O6(CLBLM_R_X65Y111_SLICE_X99Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y111_SLICE_X99Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y111_SLICE_X99Y111_BO5),
.O6(CLBLM_R_X65Y111_SLICE_X99Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaff55ff55ff)
  ) CLBLM_R_X65Y111_SLICE_X99Y111_ALUT (
.I0(CLBLM_R_X67Y111_SLICE_X101Y111_A5Q),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X67Y111_SLICE_X100Y111_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y111_SLICE_X99Y111_AO5),
.O6(CLBLM_R_X65Y111_SLICE_X99Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y96_SLICE_X100Y96_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y96_SLICE_X100Y96_DO5),
.O6(CLBLM_R_X67Y96_SLICE_X100Y96_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y96_SLICE_X100Y96_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y96_SLICE_X100Y96_CO5),
.O6(CLBLM_R_X67Y96_SLICE_X100Y96_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y96_SLICE_X100Y96_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y96_SLICE_X100Y96_BO5),
.O6(CLBLM_R_X67Y96_SLICE_X100Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y96_SLICE_X100Y96_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y96_SLICE_X100Y96_AO5),
.O6(CLBLM_R_X67Y96_SLICE_X100Y96_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y96_SLICE_X101Y96_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y96_SLICE_X101Y96_AO6),
.Q(CLBLM_R_X67Y96_SLICE_X101Y96_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y96_SLICE_X101Y96_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y96_SLICE_X101Y96_BO6),
.Q(CLBLM_R_X67Y96_SLICE_X101Y96_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y96_SLICE_X101Y96_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y96_SLICE_X101Y96_CO6),
.Q(CLBLM_R_X67Y96_SLICE_X101Y96_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y96_SLICE_X101Y96_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y96_SLICE_X101Y96_DO6),
.Q(CLBLM_R_X67Y96_SLICE_X101Y96_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f5dda0a0a088)
  ) CLBLM_R_X67Y96_SLICE_X101Y96_DLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I2(CLBLM_R_X67Y96_SLICE_X101Y96_DQ),
.I3(CLBLM_R_X67Y98_SLICE_X101Y98_CO6),
.I4(CLBLM_R_X67Y98_SLICE_X100Y98_CO5),
.I5(CLBLM_R_X67Y97_SLICE_X101Y97_DQ),
.O5(CLBLM_R_X67Y96_SLICE_X101Y96_DO5),
.O6(CLBLM_R_X67Y96_SLICE_X101Y96_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8888dfd58a80)
  ) CLBLM_R_X67Y96_SLICE_X101Y96_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_R_X67Y96_SLICE_X101Y96_CQ),
.I2(CLBLM_R_X67Y98_SLICE_X100Y98_CO5),
.I3(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I4(CLBLM_L_X68Y96_SLICE_X102Y96_AQ),
.I5(CLBLM_R_X67Y98_SLICE_X101Y98_BO6),
.O5(CLBLM_R_X67Y96_SLICE_X101Y96_CO5),
.O6(CLBLM_R_X67Y96_SLICE_X101Y96_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0f0aaccf0f0)
  ) CLBLM_R_X67Y96_SLICE_X101Y96_BLUT (
.I0(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I1(CLBLM_R_X67Y96_SLICE_X101Y96_BQ),
.I2(CLBLM_R_X67Y96_SLICE_X101Y96_DQ),
.I3(CLBLM_R_X67Y98_SLICE_X100Y98_B5Q),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_R_X67Y98_SLICE_X101Y98_CO6),
.O5(CLBLM_R_X67Y96_SLICE_X101Y96_BO5),
.O6(CLBLM_R_X67Y96_SLICE_X101Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f0aaaac0f0aaaa)
  ) CLBLM_R_X67Y96_SLICE_X101Y96_ALUT (
.I0(CLBLM_R_X67Y96_SLICE_X101Y96_CQ),
.I1(CLBLM_R_X67Y98_SLICE_X101Y98_BO6),
.I2(CLBLM_R_X67Y96_SLICE_X101Y96_AQ),
.I3(CLBLM_R_X67Y98_SLICE_X100Y98_B5Q),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.O5(CLBLM_R_X67Y96_SLICE_X101Y96_AO5),
.O6(CLBLM_R_X67Y96_SLICE_X101Y96_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y97_SLICE_X100Y97_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y97_SLICE_X100Y97_AO6),
.Q(CLBLM_R_X67Y97_SLICE_X100Y97_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y97_SLICE_X100Y97_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y97_SLICE_X100Y97_DO5),
.O6(CLBLM_R_X67Y97_SLICE_X100Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y97_SLICE_X100Y97_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y97_SLICE_X100Y97_CO5),
.O6(CLBLM_R_X67Y97_SLICE_X100Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y97_SLICE_X100Y97_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y97_SLICE_X100Y97_BO5),
.O6(CLBLM_R_X67Y97_SLICE_X100Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aaaaf0ccaaaa)
  ) CLBLM_R_X67Y97_SLICE_X100Y97_ALUT (
.I0(CLBLM_R_X67Y98_SLICE_X101Y98_DQ),
.I1(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I2(CLBLM_R_X67Y97_SLICE_X100Y97_AQ),
.I3(CLBLM_R_X67Y98_SLICE_X101Y98_CO5),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_R_X67Y98_SLICE_X100Y98_CO6),
.O5(CLBLM_R_X67Y97_SLICE_X100Y97_AO5),
.O6(CLBLM_R_X67Y97_SLICE_X100Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y97_SLICE_X101Y97_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y97_SLICE_X101Y97_AO6),
.Q(CLBLM_R_X67Y97_SLICE_X101Y97_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y97_SLICE_X101Y97_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y97_SLICE_X101Y97_BO6),
.Q(CLBLM_R_X67Y97_SLICE_X101Y97_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y97_SLICE_X101Y97_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y97_SLICE_X101Y97_CO6),
.Q(CLBLM_R_X67Y97_SLICE_X101Y97_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y97_SLICE_X101Y97_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y97_SLICE_X101Y97_DO6),
.Q(CLBLM_R_X67Y97_SLICE_X101Y97_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4e4e4eee444)
  ) CLBLM_R_X67Y97_SLICE_X101Y97_DLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_R_X67Y97_SLICE_X101Y97_CQ),
.I2(CLBLM_R_X67Y97_SLICE_X101Y97_DQ),
.I3(CLBLM_R_X67Y98_SLICE_X100Y98_CO6),
.I4(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I5(CLBLM_R_X67Y98_SLICE_X101Y98_CO6),
.O5(CLBLM_R_X67Y97_SLICE_X101Y97_DO5),
.O6(CLBLM_R_X67Y97_SLICE_X101Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00caffca00)
  ) CLBLM_R_X67Y97_SLICE_X101Y97_CLUT (
.I0(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I1(CLBLM_R_X67Y97_SLICE_X101Y97_CQ),
.I2(CLBLM_R_X67Y98_SLICE_X101Y98_AO5),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_R_X67Y97_SLICE_X101Y97_AQ),
.I5(CLBLM_R_X67Y98_SLICE_X101Y98_CO6),
.O5(CLBLM_R_X67Y97_SLICE_X101Y97_CO5),
.O6(CLBLM_R_X67Y97_SLICE_X101Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfdfcf8fc0d0c080)
  ) CLBLM_R_X67Y97_SLICE_X101Y97_BLUT (
.I0(CLBLM_R_X67Y98_SLICE_X101Y98_AO6),
.I1(CLBLM_R_X67Y97_SLICE_X101Y97_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_R_X67Y98_SLICE_X101Y98_CO5),
.I4(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I5(CLBLM_R_X67Y96_SLICE_X101Y96_BQ),
.O5(CLBLM_R_X67Y97_SLICE_X101Y97_BO5),
.O6(CLBLM_R_X67Y97_SLICE_X101Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0afa0bfb08f80)
  ) CLBLM_R_X67Y97_SLICE_X101Y97_ALUT (
.I0(CLBLM_R_X67Y97_SLICE_X101Y97_AQ),
.I1(CLBLM_R_X67Y98_SLICE_X101Y98_AO6),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_R_X67Y96_SLICE_X101Y96_AQ),
.I4(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I5(CLBLM_R_X67Y98_SLICE_X101Y98_CO6),
.O5(CLBLM_R_X67Y97_SLICE_X101Y97_AO5),
.O6(CLBLM_R_X67Y97_SLICE_X101Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y98_SLICE_X100Y98_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y98_SLICE_X100Y98_AO5),
.Q(CLBLM_R_X67Y98_SLICE_X100Y98_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y98_SLICE_X100Y98_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y98_SLICE_X100Y98_BO5),
.Q(CLBLM_R_X67Y98_SLICE_X100Y98_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y98_SLICE_X100Y98_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y98_SLICE_X100Y98_AO6),
.Q(CLBLM_R_X67Y98_SLICE_X100Y98_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y98_SLICE_X100Y98_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y98_SLICE_X100Y98_BO6),
.Q(CLBLM_R_X67Y98_SLICE_X100Y98_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y98_SLICE_X100Y98_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y98_SLICE_X100Y98_DO5),
.O6(CLBLM_R_X67Y98_SLICE_X100Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfcfcf3f3f3f3f)
  ) CLBLM_R_X67Y98_SLICE_X100Y98_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X67Y98_SLICE_X100Y98_AQ),
.I2(CLBLM_R_X67Y98_SLICE_X100Y98_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y98_SLICE_X100Y98_CO5),
.O6(CLBLM_R_X67Y98_SLICE_X100Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3cf0f04040cccc)
  ) CLBLM_R_X67Y98_SLICE_X100Y98_BLUT (
.I0(CLBLM_R_X67Y98_SLICE_X100Y98_B5Q),
.I1(CLBLM_R_X67Y98_SLICE_X100Y98_BQ),
.I2(CLBLM_R_X67Y98_SLICE_X100Y98_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLM_R_X67Y98_SLICE_X100Y98_BO5),
.O6(CLBLM_R_X67Y98_SLICE_X100Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h050500006666aaaa)
  ) CLBLM_R_X67Y98_SLICE_X100Y98_ALUT (
.I0(CLBLM_R_X67Y98_SLICE_X100Y98_B5Q),
.I1(CLBLM_R_X67Y98_SLICE_X100Y98_A5Q),
.I2(CLBLM_R_X67Y98_SLICE_X100Y98_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLM_R_X67Y98_SLICE_X100Y98_AO5),
.O6(CLBLM_R_X67Y98_SLICE_X100Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y98_SLICE_X101Y98_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y98_SLICE_X101Y98_DO6),
.Q(CLBLM_R_X67Y98_SLICE_X101Y98_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f7f3b3c0c4c080)
  ) CLBLM_R_X67Y98_SLICE_X101Y98_DLUT (
.I0(CLBLM_R_X67Y98_SLICE_X101Y98_CO5),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_R_X67Y98_SLICE_X101Y98_DQ),
.I3(CLBLM_R_X67Y98_SLICE_X101Y98_AO5),
.I4(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I5(CLBLM_R_X67Y97_SLICE_X101Y97_BQ),
.O5(CLBLM_R_X67Y98_SLICE_X101Y98_DO5),
.O6(CLBLM_R_X67Y98_SLICE_X101Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddddddd77777777)
  ) CLBLM_R_X67Y98_SLICE_X101Y98_CLUT (
.I0(CLBLM_L_X68Y101_SLICE_X102Y101_BQ),
.I1(CLBLM_R_X67Y98_SLICE_X100Y98_A5Q),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y98_SLICE_X101Y98_CO5),
.O6(CLBLM_R_X67Y98_SLICE_X101Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5555ffffaaaa)
  ) CLBLM_R_X67Y98_SLICE_X101Y98_BLUT (
.I0(CLBLM_R_X67Y98_SLICE_X100Y98_A5Q),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X68Y101_SLICE_X102Y101_BQ),
.I5(1'b1),
.O5(CLBLM_R_X67Y98_SLICE_X101Y98_BO5),
.O6(CLBLM_R_X67Y98_SLICE_X101Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffaaaaaaffff)
  ) CLBLM_R_X67Y98_SLICE_X101Y98_ALUT (
.I0(CLBLM_R_X67Y98_SLICE_X100Y98_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X67Y98_SLICE_X100Y98_B5Q),
.I4(CLBLM_R_X67Y98_SLICE_X100Y98_AQ),
.I5(1'b1),
.O5(CLBLM_R_X67Y98_SLICE_X101Y98_AO5),
.O6(CLBLM_R_X67Y98_SLICE_X101Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y99_SLICE_X100Y99_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y99_SLICE_X100Y99_AO6),
.Q(CLBLM_R_X67Y99_SLICE_X100Y99_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y99_SLICE_X100Y99_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y99_SLICE_X100Y99_BO6),
.Q(CLBLM_R_X67Y99_SLICE_X100Y99_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888888833330000)
  ) CLBLM_R_X67Y99_SLICE_X100Y99_DLUT (
.I0(CLBLM_R_X67Y101_SLICE_X100Y101_DO6),
.I1(CLBLM_R_X67Y99_SLICE_X100Y99_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X67Y101_SLICE_X101Y101_DO6),
.I5(CLBLM_R_X67Y100_SLICE_X100Y100_CQ),
.O5(CLBLM_R_X67Y99_SLICE_X100Y99_DO5),
.O6(CLBLM_R_X67Y99_SLICE_X100Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3ffffdfdfdfdf)
  ) CLBLM_R_X67Y99_SLICE_X100Y99_CLUT (
.I0(CLBLM_R_X67Y100_SLICE_X100Y100_BQ),
.I1(CLBLM_R_X67Y99_SLICE_X100Y99_AQ),
.I2(CLBLM_R_X67Y99_SLICE_X100Y99_BQ),
.I3(1'b1),
.I4(CLBLM_R_X67Y103_SLICE_X100Y103_BQ),
.I5(CLBLM_R_X67Y100_SLICE_X100Y100_CQ),
.O5(CLBLM_R_X67Y99_SLICE_X100Y99_CO5),
.O6(CLBLM_R_X67Y99_SLICE_X100Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6666f0f02222f0f0)
  ) CLBLM_R_X67Y99_SLICE_X100Y99_BLUT (
.I0(CLBLM_R_X67Y99_SLICE_X100Y99_DO6),
.I1(CLBLM_R_X67Y99_SLICE_X100Y99_BQ),
.I2(CLBLM_R_X67Y99_SLICE_X100Y99_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_R_X67Y99_SLICE_X100Y99_CO6),
.O5(CLBLM_R_X67Y99_SLICE_X100Y99_BO5),
.O6(CLBLM_R_X67Y99_SLICE_X100Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c5aff000c0aff00)
  ) CLBLM_R_X67Y99_SLICE_X100Y99_ALUT (
.I0(CLBLM_R_X67Y101_SLICE_X101Y101_DO6),
.I1(CLBLM_R_X67Y101_SLICE_X100Y101_DO6),
.I2(CLBLM_R_X67Y99_SLICE_X100Y99_AQ),
.I3(CLBLM_R_X67Y100_SLICE_X100Y100_CQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_R_X67Y99_SLICE_X100Y99_CO6),
.O5(CLBLM_R_X67Y99_SLICE_X100Y99_AO5),
.O6(CLBLM_R_X67Y99_SLICE_X100Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y99_SLICE_X101Y99_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y99_SLICE_X101Y99_DO5),
.O6(CLBLM_R_X67Y99_SLICE_X101Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y99_SLICE_X101Y99_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y99_SLICE_X101Y99_CO5),
.O6(CLBLM_R_X67Y99_SLICE_X101Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y99_SLICE_X101Y99_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y99_SLICE_X101Y99_BO5),
.O6(CLBLM_R_X67Y99_SLICE_X101Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y99_SLICE_X101Y99_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y99_SLICE_X101Y99_AO5),
.O6(CLBLM_R_X67Y99_SLICE_X101Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y100_SLICE_X100Y100_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X63Y105_SLICE_X95Y105_AQ),
.Q(CLBLM_R_X67Y100_SLICE_X100Y100_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y100_SLICE_X100Y100_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y100_SLICE_X100Y100_AO6),
.Q(CLBLM_R_X67Y100_SLICE_X100Y100_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y100_SLICE_X100Y100_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y100_SLICE_X100Y100_BO6),
.Q(CLBLM_R_X67Y100_SLICE_X100Y100_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y100_SLICE_X100Y100_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y100_SLICE_X100Y100_CO6),
.Q(CLBLM_R_X67Y100_SLICE_X100Y100_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y100_SLICE_X100Y100_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y100_SLICE_X100Y100_DO5),
.O6(CLBLM_R_X67Y100_SLICE_X100Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3632ffff36320000)
  ) CLBLM_R_X67Y100_SLICE_X100Y100_CLUT (
.I0(CLBLM_R_X67Y101_SLICE_X100Y101_DO6),
.I1(CLBLM_R_X67Y100_SLICE_X100Y100_CQ),
.I2(CLBLM_R_X67Y101_SLICE_X101Y101_DO6),
.I3(CLBLM_R_X67Y99_SLICE_X100Y99_CO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_R_X67Y101_SLICE_X101Y101_BQ),
.O5(CLBLM_R_X67Y100_SLICE_X100Y100_CO5),
.O6(CLBLM_R_X67Y100_SLICE_X100Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5d5d5d5d0a080a08)
  ) CLBLM_R_X67Y100_SLICE_X100Y100_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_R_X67Y100_SLICE_X100Y100_BQ),
.I2(CLBLL_R_X77Y104_SLICE_X119Y104_A5Q),
.I3(CLBLM_R_X63Y105_SLICE_X95Y105_AQ),
.I4(1'b1),
.I5(CLBLM_R_X67Y100_SLICE_X100Y100_A5Q),
.O5(CLBLM_R_X67Y100_SLICE_X100Y100_BO5),
.O6(CLBLM_R_X67Y100_SLICE_X100Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0acc0acc38cc38cc)
  ) CLBLM_R_X67Y100_SLICE_X100Y100_ALUT (
.I0(CLBLM_R_X67Y99_SLICE_X100Y99_CO6),
.I1(CLBLM_R_X67Y100_SLICE_X100Y100_BQ),
.I2(CLBLM_R_X67Y100_SLICE_X100Y100_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(1'b1),
.I5(CLBLM_R_X67Y103_SLICE_X100Y103_BQ),
.O5(CLBLM_R_X67Y100_SLICE_X100Y100_AO5),
.O6(CLBLM_R_X67Y100_SLICE_X100Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y100_SLICE_X101Y100_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y100_SLICE_X101Y100_DO5),
.O6(CLBLM_R_X67Y100_SLICE_X101Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y100_SLICE_X101Y100_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y100_SLICE_X101Y100_CO5),
.O6(CLBLM_R_X67Y100_SLICE_X101Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y100_SLICE_X101Y100_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y100_SLICE_X101Y100_BO5),
.O6(CLBLM_R_X67Y100_SLICE_X101Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y100_SLICE_X101Y100_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y100_SLICE_X101Y100_AO5),
.O6(CLBLM_R_X67Y100_SLICE_X101Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y101_SLICE_X100Y101_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y101_SLICE_X100Y101_AO6),
.Q(CLBLM_R_X67Y101_SLICE_X100Y101_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y101_SLICE_X100Y101_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y101_SLICE_X100Y101_CO6),
.Q(CLBLM_R_X67Y101_SLICE_X100Y101_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X67Y101_SLICE_X100Y101_DLUT (
.I0(CLBLM_R_X67Y100_SLICE_X100Y100_AQ),
.I1(CLBLM_R_X67Y101_SLICE_X100Y101_CQ),
.I2(CLBLM_R_X67Y103_SLICE_X100Y103_BQ),
.I3(CLBLM_R_X67Y101_SLICE_X101Y101_AQ),
.I4(CLBLM_R_X67Y101_SLICE_X100Y101_AQ),
.I5(CLBLM_R_X67Y101_SLICE_X101Y101_BQ),
.O5(CLBLM_R_X67Y101_SLICE_X100Y101_DO5),
.O6(CLBLM_R_X67Y101_SLICE_X100Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777dd5522228800)
  ) CLBLM_R_X67Y101_SLICE_X100Y101_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_R_X67Y101_SLICE_X100Y101_CQ),
.I2(1'b1),
.I3(CLBLM_R_X67Y99_SLICE_X100Y99_CO6),
.I4(CLBLM_R_X67Y101_SLICE_X100Y101_BO5),
.I5(CLBLM_R_X67Y101_SLICE_X100Y101_AQ),
.O5(CLBLM_R_X67Y101_SLICE_X100Y101_CO5),
.O6(CLBLM_R_X67Y101_SLICE_X100Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc303c00081018000)
  ) CLBLM_R_X67Y101_SLICE_X100Y101_BLUT (
.I0(CLBLM_R_X67Y101_SLICE_X100Y101_AQ),
.I1(CLBLM_R_X67Y101_SLICE_X101Y101_AQ),
.I2(CLBLM_R_X67Y100_SLICE_X100Y100_AQ),
.I3(CLBLM_R_X67Y103_SLICE_X100Y103_BQ),
.I4(CLBLM_R_X67Y100_SLICE_X100Y100_BQ),
.I5(1'b1),
.O5(CLBLM_R_X67Y101_SLICE_X100Y101_BO5),
.O6(CLBLM_R_X67Y101_SLICE_X100Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3ff30cc03f330c00)
  ) CLBLM_R_X67Y101_SLICE_X100Y101_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_R_X67Y101_SLICE_X100Y101_AQ),
.I3(CLBLM_R_X67Y101_SLICE_X100Y101_BO6),
.I4(CLBLM_R_X67Y101_SLICE_X101Y101_AQ),
.I5(CLBLM_R_X67Y99_SLICE_X100Y99_CO6),
.O5(CLBLM_R_X67Y101_SLICE_X100Y101_AO5),
.O6(CLBLM_R_X67Y101_SLICE_X100Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y101_SLICE_X101Y101_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y101_SLICE_X101Y101_AO6),
.Q(CLBLM_R_X67Y101_SLICE_X101Y101_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y101_SLICE_X101Y101_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y101_SLICE_X101Y101_BO6),
.Q(CLBLM_R_X67Y101_SLICE_X101Y101_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000010000)
  ) CLBLM_R_X67Y101_SLICE_X101Y101_DLUT (
.I0(CLBLM_R_X67Y100_SLICE_X100Y100_AQ),
.I1(CLBLM_R_X67Y101_SLICE_X100Y101_AQ),
.I2(CLBLM_R_X67Y101_SLICE_X101Y101_BQ),
.I3(CLBLM_R_X67Y101_SLICE_X100Y101_CQ),
.I4(CLBLM_R_X67Y100_SLICE_X100Y100_BQ),
.I5(CLBLM_R_X67Y101_SLICE_X101Y101_AQ),
.O5(CLBLM_R_X67Y101_SLICE_X101Y101_DO5),
.O6(CLBLM_R_X67Y101_SLICE_X101Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000800000050000)
  ) CLBLM_R_X67Y101_SLICE_X101Y101_CLUT (
.I0(CLBLM_R_X67Y100_SLICE_X100Y100_AQ),
.I1(CLBLM_R_X67Y103_SLICE_X100Y103_BQ),
.I2(CLBLM_R_X67Y101_SLICE_X100Y101_AQ),
.I3(CLBLM_R_X67Y101_SLICE_X100Y101_CQ),
.I4(CLBLM_R_X67Y100_SLICE_X100Y100_BQ),
.I5(CLBLM_R_X67Y101_SLICE_X101Y101_AQ),
.O5(CLBLM_R_X67Y101_SLICE_X101Y101_CO5),
.O6(CLBLM_R_X67Y101_SLICE_X101Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff88ff33008800)
  ) CLBLM_R_X67Y101_SLICE_X101Y101_BLUT (
.I0(CLBLM_R_X67Y99_SLICE_X100Y99_CO6),
.I1(CLBLM_R_X67Y101_SLICE_X101Y101_BQ),
.I2(1'b1),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_R_X67Y101_SLICE_X101Y101_CO6),
.I5(CLBLM_R_X67Y101_SLICE_X100Y101_CQ),
.O5(CLBLM_R_X67Y101_SLICE_X101Y101_BO5),
.O6(CLBLM_R_X67Y101_SLICE_X101Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h20cff0f02ac0f0f0)
  ) CLBLM_R_X67Y101_SLICE_X101Y101_ALUT (
.I0(CLBLM_R_X67Y99_SLICE_X100Y99_CO6),
.I1(CLBLM_R_X67Y103_SLICE_X100Y103_BQ),
.I2(CLBLM_R_X67Y100_SLICE_X100Y100_AQ),
.I3(CLBLM_R_X67Y101_SLICE_X101Y101_AQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_R_X67Y100_SLICE_X100Y100_BQ),
.O5(CLBLM_R_X67Y101_SLICE_X101Y101_AO5),
.O6(CLBLM_R_X67Y101_SLICE_X101Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y103_SLICE_X100Y103_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y103_SLICE_X100Y103_AO5),
.Q(CLBLM_R_X67Y103_SLICE_X100Y103_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y103_SLICE_X100Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X77Y104_SLICE_X119Y104_A5Q),
.Q(CLBLM_R_X67Y103_SLICE_X100Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y103_SLICE_X100Y103_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y103_SLICE_X100Y103_BO6),
.Q(CLBLM_R_X67Y103_SLICE_X100Y103_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y103_SLICE_X100Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y103_SLICE_X100Y103_DO5),
.O6(CLBLM_R_X67Y103_SLICE_X100Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y103_SLICE_X100Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y103_SLICE_X100Y103_CO5),
.O6(CLBLM_R_X67Y103_SLICE_X100Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5050dad85050dad8)
  ) CLBLM_R_X67Y103_SLICE_X100Y103_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_R_X67Y103_SLICE_X100Y103_BQ),
.I2(CLBLM_R_X67Y103_SLICE_X100Y103_AQ),
.I3(CLBLL_R_X77Y104_SLICE_X119Y104_A5Q),
.I4(CLBLM_R_X63Y105_SLICE_X95Y105_AQ),
.I5(1'b1),
.O5(CLBLM_R_X67Y103_SLICE_X100Y103_BO5),
.O6(CLBLM_R_X67Y103_SLICE_X100Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccc0c074b874b8)
  ) CLBLM_R_X67Y103_SLICE_X100Y103_ALUT (
.I0(CLBLM_R_X67Y103_SLICE_X100Y103_B5Q),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_L_X68Y103_SLICE_X102Y103_B5Q),
.I3(CLBLM_L_X68Y99_SLICE_X102Y99_AO5),
.I4(CLBLM_L_X68Y103_SLICE_X102Y103_DQ),
.I5(1'b1),
.O5(CLBLM_R_X67Y103_SLICE_X100Y103_AO5),
.O6(CLBLM_R_X67Y103_SLICE_X100Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y103_SLICE_X101Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y103_SLICE_X101Y103_AO6),
.Q(CLBLM_R_X67Y103_SLICE_X101Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y103_SLICE_X101Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y103_SLICE_X101Y103_DO5),
.O6(CLBLM_R_X67Y103_SLICE_X101Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y103_SLICE_X101Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y103_SLICE_X101Y103_CO5),
.O6(CLBLM_R_X67Y103_SLICE_X101Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y103_SLICE_X101Y103_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y103_SLICE_X101Y103_BO5),
.O6(CLBLM_R_X67Y103_SLICE_X101Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4ee4e4e4e4e4e4e4)
  ) CLBLM_R_X67Y103_SLICE_X101Y103_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X68Y102_SLICE_X102Y102_CQ),
.I2(CLBLM_R_X67Y103_SLICE_X101Y103_AQ),
.I3(CLBLM_L_X68Y101_SLICE_X102Y101_BQ),
.I4(CLBLM_R_X67Y98_SLICE_X100Y98_B5Q),
.I5(CLBLM_R_X67Y98_SLICE_X100Y98_A5Q),
.O5(CLBLM_R_X67Y103_SLICE_X101Y103_AO5),
.O6(CLBLM_R_X67Y103_SLICE_X101Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0505050500330033)
  ) CLBLM_R_X67Y105_SLICE_X100Y105_DLUT (
.I0(CLBLM_L_X72Y105_SLICE_X109Y105_B5Q),
.I1(CLBLM_R_X65Y105_SLICE_X98Y105_CQ),
.I2(CLBLM_L_X72Y104_SLICE_X108Y104_CQ),
.I3(CLBLM_R_X65Y106_SLICE_X99Y106_C5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y105_SLICE_X100Y105_DO5),
.O6(CLBLM_R_X67Y105_SLICE_X100Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0505050500330033)
  ) CLBLM_R_X67Y105_SLICE_X100Y105_CLUT (
.I0(CLBLL_R_X71Y109_SLICE_X106Y109_AQ),
.I1(CLBLM_R_X65Y100_SLICE_X99Y100_CQ),
.I2(CLBLL_R_X71Y108_SLICE_X106Y108_D5Q),
.I3(CLBLM_R_X65Y100_SLICE_X99Y100_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y105_SLICE_X100Y105_CO5),
.O6(CLBLM_R_X67Y105_SLICE_X100Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000a0b0f0002000b)
  ) CLBLM_R_X67Y105_SLICE_X100Y105_BLUT (
.I0(CLBLM_R_X67Y105_SLICE_X100Y105_DO6),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_R_X67Y103_SLICE_X100Y103_AO6),
.I3(CLBLM_R_X67Y108_SLICE_X100Y108_BO6),
.I4(CLBLM_R_X65Y105_SLICE_X99Y105_AO6),
.I5(CLBLM_R_X67Y105_SLICE_X100Y105_CO6),
.O5(CLBLM_R_X67Y105_SLICE_X100Y105_BO5),
.O6(CLBLM_R_X67Y105_SLICE_X100Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff00fffdff00)
  ) CLBLM_R_X67Y105_SLICE_X100Y105_ALUT (
.I0(CLBLM_R_X67Y105_SLICE_X100Y105_DO6),
.I1(CLBLM_L_X68Y103_SLICE_X102Y103_B5Q),
.I2(CLBLM_L_X68Y103_SLICE_X102Y103_DQ),
.I3(CLBLM_L_X68Y105_SLICE_X102Y105_AO6),
.I4(CLBLM_R_X65Y101_SLICE_X99Y101_AO6),
.I5(CLBLM_R_X67Y108_SLICE_X100Y108_BO6),
.O5(CLBLM_R_X67Y105_SLICE_X100Y105_AO5),
.O6(CLBLM_R_X67Y105_SLICE_X100Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000011112120)
  ) CLBLM_R_X67Y105_SLICE_X101Y105_DLUT (
.I0(CLBLM_R_X65Y105_SLICE_X99Y105_BO6),
.I1(CLBLM_R_X67Y105_SLICE_X100Y105_AO6),
.I2(CLBLM_R_X67Y105_SLICE_X100Y105_CO5),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_R_X67Y103_SLICE_X100Y103_AO6),
.I5(CLBLM_R_X67Y105_SLICE_X101Y105_BO6),
.O5(CLBLM_R_X67Y105_SLICE_X101Y105_DO5),
.O6(CLBLM_R_X67Y105_SLICE_X101Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f00000f1f0000)
  ) CLBLM_R_X67Y105_SLICE_X101Y105_CLUT (
.I0(CLBLM_L_X68Y103_SLICE_X102Y103_B5Q),
.I1(CLBLM_L_X72Y104_SLICE_X108Y104_CQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_L_X68Y103_SLICE_X102Y103_DQ),
.I4(CLBLM_R_X67Y108_SLICE_X100Y108_BO5),
.I5(CLBLM_L_X72Y105_SLICE_X109Y105_B5Q),
.O5(CLBLM_R_X67Y105_SLICE_X101Y105_CO5),
.O6(CLBLM_R_X67Y105_SLICE_X101Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaffaaffaaffa8)
  ) CLBLM_R_X67Y105_SLICE_X101Y105_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_L_X72Y104_SLICE_X108Y104_CQ),
.I2(CLBLM_L_X72Y105_SLICE_X109Y105_B5Q),
.I3(CLBLM_R_X67Y108_SLICE_X100Y108_BO6),
.I4(CLBLL_R_X71Y109_SLICE_X106Y109_AQ),
.I5(CLBLL_R_X71Y108_SLICE_X106Y108_D5Q),
.O5(CLBLM_R_X67Y105_SLICE_X101Y105_BO5),
.O6(CLBLM_R_X67Y105_SLICE_X101Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0eff04ff04ff04)
  ) CLBLM_R_X67Y105_SLICE_X101Y105_ALUT (
.I0(CLBLM_L_X68Y105_SLICE_X102Y105_AO5),
.I1(CLBLM_R_X67Y105_SLICE_X100Y105_BO6),
.I2(CLBLM_R_X65Y105_SLICE_X99Y105_BO5),
.I3(CLBLM_R_X67Y105_SLICE_X101Y105_DO6),
.I4(CLBLM_R_X67Y105_SLICE_X100Y105_DO5),
.I5(CLBLM_R_X67Y105_SLICE_X101Y105_CO6),
.O5(CLBLM_R_X67Y105_SLICE_X101Y105_AO5),
.O6(CLBLM_R_X67Y105_SLICE_X101Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y108_SLICE_X100Y108_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y108_SLICE_X100Y108_CO5),
.Q(CLBLM_R_X67Y108_SLICE_X100Y108_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y108_SLICE_X100Y108_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y108_SLICE_X100Y108_AO5),
.Q(CLBLM_R_X67Y108_SLICE_X100Y108_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y108_SLICE_X100Y108_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y108_SLICE_X100Y108_CO6),
.Q(CLBLM_R_X67Y108_SLICE_X100Y108_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y108_SLICE_X100Y108_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y108_SLICE_X100Y108_DO6),
.Q(CLBLM_R_X67Y108_SLICE_X100Y108_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d87272ffff0000)
  ) CLBLM_R_X67Y108_SLICE_X100Y108_DLUT (
.I0(CLBLM_R_X67Y111_SLICE_X100Y111_CO5),
.I1(CLBLM_R_X67Y108_SLICE_X100Y108_AQ),
.I2(CLBLM_R_X67Y108_SLICE_X100Y108_DQ),
.I3(1'b1),
.I4(CLBLM_R_X67Y109_SLICE_X100Y109_CQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_R_X67Y108_SLICE_X100Y108_DO5),
.O6(CLBLM_R_X67Y108_SLICE_X100Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcff0c00cacc3acc)
  ) CLBLM_R_X67Y108_SLICE_X100Y108_CLUT (
.I0(CLBLM_R_X67Y108_SLICE_X100Y108_C5Q),
.I1(CLBLM_R_X67Y108_SLICE_X100Y108_CQ),
.I2(CLBLM_R_X67Y108_SLICE_X101Y108_AO6),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_R_X67Y108_SLICE_X101Y108_BQ),
.I5(1'b1),
.O5(CLBLM_R_X67Y108_SLICE_X100Y108_CO5),
.O6(CLBLM_R_X67Y108_SLICE_X100Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa888855555557)
  ) CLBLM_R_X67Y108_SLICE_X100Y108_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_R_X67Y108_SLICE_X100Y108_DQ),
.I2(CLBLL_R_X71Y109_SLICE_X106Y109_AQ),
.I3(CLBLL_R_X71Y108_SLICE_X106Y108_D5Q),
.I4(CLBLM_R_X67Y108_SLICE_X100Y108_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X67Y108_SLICE_X100Y108_BO5),
.O6(CLBLM_R_X67Y108_SLICE_X100Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0c0c0c5faf50a0)
  ) CLBLM_R_X67Y108_SLICE_X100Y108_ALUT (
.I0(CLBLM_R_X67Y108_SLICE_X101Y108_AO6),
.I1(CLBLM_L_X72Y105_SLICE_X108Y105_AQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_R_X67Y108_SLICE_X100Y108_AQ),
.I4(CLBLM_R_X67Y108_SLICE_X100Y108_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X67Y108_SLICE_X100Y108_AO5),
.O6(CLBLM_R_X67Y108_SLICE_X100Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y108_SLICE_X101Y108_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y108_SLICE_X101Y108_BO6),
.Q(CLBLM_R_X67Y108_SLICE_X101Y108_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y108_SLICE_X101Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y108_SLICE_X101Y108_DO5),
.O6(CLBLM_R_X67Y108_SLICE_X101Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y108_SLICE_X101Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y108_SLICE_X101Y108_CO5),
.O6(CLBLM_R_X67Y108_SLICE_X101Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cccaaaaccccaaaa)
  ) CLBLM_R_X67Y108_SLICE_X101Y108_BLUT (
.I0(CLBLM_R_X67Y109_SLICE_X100Y109_BQ),
.I1(CLBLM_R_X67Y108_SLICE_X101Y108_BQ),
.I2(CLBLM_R_X67Y111_SLICE_X101Y111_B5Q),
.I3(CLBLM_R_X67Y111_SLICE_X101Y111_A5Q),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_R_X67Y111_SLICE_X100Y111_A5Q),
.O5(CLBLM_R_X67Y108_SLICE_X101Y108_BO5),
.O6(CLBLM_R_X67Y108_SLICE_X101Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h800000007f7fffff)
  ) CLBLM_R_X67Y108_SLICE_X101Y108_ALUT (
.I0(CLBLM_L_X68Y109_SLICE_X102Y109_A5Q),
.I1(CLBLM_L_X68Y108_SLICE_X102Y108_A5Q),
.I2(CLBLM_L_X68Y108_SLICE_X102Y108_AQ),
.I3(CLBLM_L_X70Y106_SLICE_X105Y106_DO6),
.I4(CLBLM_L_X62Y92_SLICE_X92Y92_BQ),
.I5(1'b1),
.O5(CLBLM_R_X67Y108_SLICE_X101Y108_AO5),
.O6(CLBLM_R_X67Y108_SLICE_X101Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y109_SLICE_X100Y109_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y109_SLICE_X100Y109_AO6),
.Q(CLBLM_R_X67Y109_SLICE_X100Y109_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y109_SLICE_X100Y109_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y109_SLICE_X100Y109_BO6),
.Q(CLBLM_R_X67Y109_SLICE_X100Y109_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y109_SLICE_X100Y109_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y109_SLICE_X100Y109_CO6),
.Q(CLBLM_R_X67Y109_SLICE_X100Y109_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h66666666a0000000)
  ) CLBLM_R_X67Y109_SLICE_X100Y109_DLUT (
.I0(CLBLM_R_X65Y111_SLICE_X98Y111_AQ),
.I1(CLBLM_L_X68Y109_SLICE_X102Y109_A5Q),
.I2(CLBLM_L_X76Y111_SLICE_X116Y111_AQ),
.I3(CLBLM_L_X60Y97_SLICE_X91Y97_AQ),
.I4(CLBLM_R_X65Y110_SLICE_X99Y110_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X67Y109_SLICE_X100Y109_DO5),
.O6(CLBLM_R_X67Y109_SLICE_X100Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heccc4cccffff0000)
  ) CLBLM_R_X67Y109_SLICE_X100Y109_CLUT (
.I0(CLBLM_R_X67Y111_SLICE_X101Y111_B5Q),
.I1(CLBLM_R_X67Y109_SLICE_X100Y109_CQ),
.I2(CLBLM_R_X67Y111_SLICE_X101Y111_A5Q),
.I3(CLBLM_R_X67Y111_SLICE_X100Y111_A5Q),
.I4(CLBLM_R_X67Y108_SLICE_X100Y108_AQ),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_R_X67Y109_SLICE_X100Y109_CO5),
.O6(CLBLM_R_X67Y109_SLICE_X100Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5accccf0f0f0f0)
  ) CLBLM_R_X67Y109_SLICE_X100Y109_BLUT (
.I0(CLBLM_R_X67Y111_SLICE_X100Y111_AQ),
.I1(CLBLM_R_X67Y109_SLICE_X100Y109_BQ),
.I2(CLBLM_R_X67Y109_SLICE_X100Y109_AQ),
.I3(1'b1),
.I4(CLBLM_R_X67Y108_SLICE_X101Y108_AO6),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_R_X67Y109_SLICE_X100Y109_BO5),
.O6(CLBLM_R_X67Y109_SLICE_X100Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000ff0aaaaaaaa)
  ) CLBLM_R_X67Y109_SLICE_X100Y109_ALUT (
.I0(CLBLM_R_X67Y111_SLICE_X100Y111_AQ),
.I1(1'b1),
.I2(CLBLM_R_X67Y109_SLICE_X100Y109_AQ),
.I3(CLBLM_L_X68Y109_SLICE_X102Y109_CO6),
.I4(CLBLM_R_X67Y108_SLICE_X101Y108_AO6),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_R_X67Y109_SLICE_X100Y109_AO5),
.O6(CLBLM_R_X67Y109_SLICE_X100Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y109_SLICE_X101Y109_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y109_SLICE_X101Y109_AO6),
.Q(CLBLM_R_X67Y109_SLICE_X101Y109_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y109_SLICE_X101Y109_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y109_SLICE_X101Y109_BO6),
.Q(CLBLM_R_X67Y109_SLICE_X101Y109_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hddfdddffddffddff)
  ) CLBLM_R_X67Y109_SLICE_X101Y109_DLUT (
.I0(CLBLM_L_X68Y108_SLICE_X102Y108_AQ),
.I1(CLBLM_L_X68Y108_SLICE_X102Y108_A5Q),
.I2(CLBLM_R_X67Y109_SLICE_X100Y109_DO6),
.I3(CLBLM_R_X67Y109_SLICE_X101Y109_CO6),
.I4(CLBLM_L_X76Y111_SLICE_X116Y111_AQ),
.I5(CLBLM_R_X67Y110_SLICE_X101Y110_BQ),
.O5(CLBLM_R_X67Y109_SLICE_X101Y109_DO5),
.O6(CLBLM_R_X67Y109_SLICE_X101Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888f000f8880000)
  ) CLBLM_R_X67Y109_SLICE_X101Y109_CLUT (
.I0(CLBLM_R_X65Y110_SLICE_X99Y110_CQ),
.I1(CLBLM_R_X67Y110_SLICE_X101Y110_CQ),
.I2(CLBLM_R_X67Y110_SLICE_X100Y110_CQ),
.I3(CLBLM_L_X60Y97_SLICE_X91Y97_AQ),
.I4(CLBLM_L_X68Y109_SLICE_X102Y109_A5Q),
.I5(CLBLM_R_X65Y111_SLICE_X98Y111_AQ),
.O5(CLBLM_R_X67Y109_SLICE_X101Y109_CO5),
.O6(CLBLM_R_X67Y109_SLICE_X101Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfdfcf8fc0d0c080)
  ) CLBLM_R_X67Y109_SLICE_X101Y109_BLUT (
.I0(CLBLM_R_X65Y110_SLICE_X99Y110_AO5),
.I1(CLBLM_R_X67Y109_SLICE_X101Y109_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_R_X67Y111_SLICE_X101Y111_DO5),
.I4(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I5(CLBLM_R_X67Y110_SLICE_X101Y110_CQ),
.O5(CLBLM_R_X67Y109_SLICE_X101Y109_BO5),
.O6(CLBLM_R_X67Y109_SLICE_X101Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4e4eee444e4)
  ) CLBLM_R_X67Y109_SLICE_X101Y109_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_R_X67Y109_SLICE_X101Y109_BQ),
.I2(CLBLM_R_X67Y109_SLICE_X101Y109_AQ),
.I3(CLBLM_R_X67Y111_SLICE_X101Y111_B5Q),
.I4(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I5(CLBLM_R_X65Y110_SLICE_X99Y110_AO5),
.O5(CLBLM_R_X67Y109_SLICE_X101Y109_AO5),
.O6(CLBLM_R_X67Y109_SLICE_X101Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y110_SLICE_X100Y110_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y110_SLICE_X100Y110_AO6),
.Q(CLBLM_R_X67Y110_SLICE_X100Y110_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y110_SLICE_X100Y110_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y110_SLICE_X100Y110_BO6),
.Q(CLBLM_R_X67Y110_SLICE_X100Y110_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y110_SLICE_X100Y110_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y110_SLICE_X100Y110_CO6),
.Q(CLBLM_R_X67Y110_SLICE_X100Y110_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9180110080800000)
  ) CLBLM_R_X67Y110_SLICE_X100Y110_DLUT (
.I0(CLBLM_L_X68Y108_SLICE_X102Y108_AQ),
.I1(CLBLM_L_X68Y108_SLICE_X102Y108_A5Q),
.I2(CLBLM_R_X67Y110_SLICE_X100Y110_AQ),
.I3(CLBLM_R_X67Y110_SLICE_X100Y110_BQ),
.I4(CLBLM_R_X65Y110_SLICE_X99Y110_B5Q),
.I5(CLBLM_L_X60Y97_SLICE_X91Y97_AQ),
.O5(CLBLM_R_X67Y110_SLICE_X100Y110_DO5),
.O6(CLBLM_R_X67Y110_SLICE_X100Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8888dfd58a80)
  ) CLBLM_R_X67Y110_SLICE_X100Y110_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_R_X67Y110_SLICE_X100Y110_CQ),
.I2(CLBLM_R_X65Y111_SLICE_X99Y111_AO5),
.I3(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I4(CLBLM_R_X65Y110_SLICE_X98Y110_DQ),
.I5(CLBLM_R_X67Y111_SLICE_X101Y111_DO5),
.O5(CLBLM_R_X67Y110_SLICE_X100Y110_CO5),
.O6(CLBLM_R_X67Y110_SLICE_X100Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8d8fad8d8d850)
  ) CLBLM_R_X67Y110_SLICE_X100Y110_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_R_X67Y110_SLICE_X100Y110_BQ),
.I2(CLBLM_R_X67Y110_SLICE_X100Y110_AQ),
.I3(CLBLM_R_X67Y111_SLICE_X101Y111_DO5),
.I4(CLBLM_R_X65Y110_SLICE_X99Y110_AO6),
.I5(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.O5(CLBLM_R_X67Y110_SLICE_X100Y110_BO5),
.O6(CLBLM_R_X67Y110_SLICE_X100Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3c0f7c4f3c0b380)
  ) CLBLM_R_X67Y110_SLICE_X100Y110_ALUT (
.I0(CLBLM_R_X67Y111_SLICE_X101Y111_DO6),
.I1(RIOB33_X105Y51_IOB_X1Y51_I),
.I2(CLBLM_R_X67Y110_SLICE_X100Y110_AQ),
.I3(CLBLM_R_X67Y110_SLICE_X101Y110_BQ),
.I4(CLBLM_R_X65Y110_SLICE_X99Y110_AO6),
.I5(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.O5(CLBLM_R_X67Y110_SLICE_X100Y110_AO5),
.O6(CLBLM_R_X67Y110_SLICE_X100Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y110_SLICE_X101Y110_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y110_SLICE_X101Y110_AO6),
.Q(CLBLM_R_X67Y110_SLICE_X101Y110_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y110_SLICE_X101Y110_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y110_SLICE_X101Y110_BO6),
.Q(CLBLM_R_X67Y110_SLICE_X101Y110_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y110_SLICE_X101Y110_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y110_SLICE_X101Y110_CO6),
.Q(CLBLM_R_X67Y110_SLICE_X101Y110_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y110_SLICE_X101Y110_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y110_SLICE_X101Y110_DO6),
.Q(CLBLM_R_X67Y110_SLICE_X101Y110_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8d8d8ff00ff00)
  ) CLBLM_R_X67Y110_SLICE_X101Y110_DLUT (
.I0(CLBLM_R_X67Y111_SLICE_X100Y111_CO5),
.I1(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I2(CLBLM_R_X67Y110_SLICE_X101Y110_DQ),
.I3(CLBLM_R_X67Y110_SLICE_X100Y110_CQ),
.I4(1'b1),
.I5(RIOB33_X105Y51_IOB_X1Y51_I),
.O5(CLBLM_R_X67Y110_SLICE_X101Y110_DO5),
.O6(CLBLM_R_X67Y110_SLICE_X101Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddfddd5888a8880)
  ) CLBLM_R_X67Y110_SLICE_X101Y110_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_R_X67Y110_SLICE_X101Y110_CQ),
.I2(CLBLM_R_X67Y111_SLICE_X101Y111_DO6),
.I3(CLBLM_R_X65Y110_SLICE_X99Y110_AO5),
.I4(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I5(CLBLM_R_X65Y110_SLICE_X99Y110_BQ),
.O5(CLBLM_R_X67Y110_SLICE_X101Y110_CO5),
.O6(CLBLM_R_X67Y110_SLICE_X101Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8d8fad8d8d850)
  ) CLBLM_R_X67Y110_SLICE_X101Y110_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_R_X67Y110_SLICE_X101Y110_BQ),
.I2(CLBLM_R_X67Y110_SLICE_X101Y110_AQ),
.I3(CLBLM_R_X67Y111_SLICE_X101Y111_CO5),
.I4(CLBLM_R_X65Y110_SLICE_X99Y110_AO6),
.I5(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.O5(CLBLM_R_X67Y110_SLICE_X101Y110_BO5),
.O6(CLBLM_R_X67Y110_SLICE_X101Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000e2ffe200)
  ) CLBLM_R_X67Y110_SLICE_X101Y110_ALUT (
.I0(CLBLL_R_X79Y96_SLICE_X122Y96_AO6),
.I1(CLBLM_R_X65Y110_SLICE_X99Y110_AO6),
.I2(CLBLM_R_X67Y110_SLICE_X101Y110_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_R_X67Y109_SLICE_X101Y109_AQ),
.I5(CLBLM_R_X67Y111_SLICE_X101Y111_CO6),
.O5(CLBLM_R_X67Y110_SLICE_X101Y110_AO5),
.O6(CLBLM_R_X67Y110_SLICE_X101Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y111_SLICE_X100Y111_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y111_SLICE_X100Y111_CO6),
.Q(CLBLM_R_X67Y111_SLICE_X100Y111_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y111_SLICE_X100Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y111_SLICE_X100Y111_AO6),
.Q(CLBLM_R_X67Y111_SLICE_X100Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y111_SLICE_X100Y111_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y111_SLICE_X100Y111_BO6),
.Q(CLBLM_R_X67Y111_SLICE_X100Y111_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y111_SLICE_X100Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y111_SLICE_X100Y111_DO5),
.O6(CLBLM_R_X67Y111_SLICE_X100Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6ec46ec4c000c000)
  ) CLBLM_R_X67Y111_SLICE_X100Y111_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_R_X67Y111_SLICE_X101Y111_A5Q),
.I2(CLBLM_R_X67Y111_SLICE_X101Y111_B5Q),
.I3(CLBLM_R_X67Y111_SLICE_X100Y111_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y111_SLICE_X100Y111_CO5),
.O6(CLBLM_R_X67Y111_SLICE_X100Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0888a22288882222)
  ) CLBLM_R_X67Y111_SLICE_X100Y111_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_R_X67Y111_SLICE_X100Y111_BQ),
.I2(CLBLM_R_X67Y111_SLICE_X101Y111_B5Q),
.I3(CLBLM_R_X67Y111_SLICE_X101Y111_A5Q),
.I4(CLBLL_R_X79Y99_SLICE_X122Y99_AO6),
.I5(CLBLM_R_X67Y111_SLICE_X100Y111_A5Q),
.O5(CLBLM_R_X67Y111_SLICE_X100Y111_BO5),
.O6(CLBLM_R_X67Y111_SLICE_X100Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8f0ccccf0f0cccc)
  ) CLBLM_R_X67Y111_SLICE_X100Y111_ALUT (
.I0(CLBLM_R_X67Y111_SLICE_X101Y111_B5Q),
.I1(CLBLM_R_X67Y111_SLICE_X100Y111_BQ),
.I2(CLBLM_R_X67Y111_SLICE_X100Y111_AQ),
.I3(CLBLM_R_X67Y111_SLICE_X101Y111_A5Q),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_R_X67Y111_SLICE_X100Y111_A5Q),
.O5(CLBLM_R_X67Y111_SLICE_X100Y111_AO5),
.O6(CLBLM_R_X67Y111_SLICE_X100Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y111_SLICE_X101Y111_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y111_SLICE_X101Y111_AO5),
.Q(CLBLM_R_X67Y111_SLICE_X101Y111_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y111_SLICE_X101Y111_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y111_SLICE_X101Y111_BO5),
.Q(CLBLM_R_X67Y111_SLICE_X101Y111_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y111_SLICE_X101Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y111_SLICE_X101Y111_AO6),
.Q(CLBLM_R_X67Y111_SLICE_X101Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y111_SLICE_X101Y111_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y111_SLICE_X101Y111_BO6),
.Q(CLBLM_R_X67Y111_SLICE_X101Y111_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fff0f0fff0fff)
  ) CLBLM_R_X67Y111_SLICE_X101Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X67Y111_SLICE_X101Y111_BQ),
.I3(CLBLM_R_X67Y111_SLICE_X101Y111_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y111_SLICE_X101Y111_DO5),
.O6(CLBLM_R_X67Y111_SLICE_X101Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffafaf0f0ffff)
  ) CLBLM_R_X67Y111_SLICE_X101Y111_CLUT (
.I0(CLBLM_R_X67Y111_SLICE_X101Y111_B5Q),
.I1(1'b1),
.I2(CLBLM_R_X67Y111_SLICE_X101Y111_BQ),
.I3(1'b1),
.I4(CLBLM_R_X67Y111_SLICE_X101Y111_AQ),
.I5(1'b1),
.O5(CLBLM_R_X67Y111_SLICE_X101Y111_CO5),
.O6(CLBLM_R_X67Y111_SLICE_X101Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a6a6a6a0c8c0c8c)
  ) CLBLM_R_X67Y111_SLICE_X101Y111_BLUT (
.I0(CLBLM_R_X67Y111_SLICE_X101Y111_AQ),
.I1(CLBLM_R_X67Y111_SLICE_X101Y111_BQ),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_R_X67Y111_SLICE_X101Y111_B5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y111_SLICE_X101Y111_BO5),
.O6(CLBLM_R_X67Y111_SLICE_X101Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h005000503fc03fc0)
  ) CLBLM_R_X67Y111_SLICE_X101Y111_ALUT (
.I0(CLBLM_R_X67Y111_SLICE_X101Y111_AQ),
.I1(CLBLM_R_X67Y111_SLICE_X101Y111_A5Q),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_R_X67Y111_SLICE_X101Y111_B5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y111_SLICE_X101Y111_AO5),
.O6(CLBLM_R_X67Y111_SLICE_X101Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y115_SLICE_X100Y115_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y115_SLICE_X100Y115_AO5),
.Q(CLBLM_R_X67Y115_SLICE_X100Y115_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y115_SLICE_X100Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y115_SLICE_X100Y115_AO6),
.Q(CLBLM_R_X67Y115_SLICE_X100Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y115_SLICE_X100Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y115_SLICE_X100Y115_DO5),
.O6(CLBLM_R_X67Y115_SLICE_X100Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y115_SLICE_X100Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y115_SLICE_X100Y115_CO5),
.O6(CLBLM_R_X67Y115_SLICE_X100Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y115_SLICE_X100Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y115_SLICE_X100Y115_BO5),
.O6(CLBLM_R_X67Y115_SLICE_X100Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00fff000f0)
  ) CLBLM_R_X67Y115_SLICE_X100Y115_ALUT (
.I0(RIOB33_X105Y53_IOB_X1Y54_I),
.I1(1'b1),
.I2(CLBLM_R_X67Y115_SLICE_X100Y115_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(RIOB33_X105Y53_IOB_X1Y53_I),
.I5(1'b1),
.O5(CLBLM_R_X67Y115_SLICE_X100Y115_AO5),
.O6(CLBLM_R_X67Y115_SLICE_X100Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y115_SLICE_X101Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y115_SLICE_X101Y115_DO5),
.O6(CLBLM_R_X67Y115_SLICE_X101Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y115_SLICE_X101Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y115_SLICE_X101Y115_CO5),
.O6(CLBLM_R_X67Y115_SLICE_X101Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y115_SLICE_X101Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y115_SLICE_X101Y115_BO5),
.O6(CLBLM_R_X67Y115_SLICE_X101Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y115_SLICE_X101Y115_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y115_SLICE_X101Y115_AO5),
.O6(CLBLM_R_X67Y115_SLICE_X101Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y116_SLICE_X100Y116_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y116_SLICE_X100Y116_BO5),
.Q(CLBLM_R_X67Y116_SLICE_X100Y116_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y116_SLICE_X100Y116_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y116_SLICE_X100Y116_CO5),
.Q(CLBLM_R_X67Y116_SLICE_X100Y116_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y116_SLICE_X100Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y116_SLICE_X100Y116_AO6),
.Q(CLBLM_R_X67Y116_SLICE_X100Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y116_SLICE_X100Y116_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y116_SLICE_X100Y116_BO6),
.Q(CLBLM_R_X67Y116_SLICE_X100Y116_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y116_SLICE_X100Y116_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y116_SLICE_X100Y116_CO6),
.Q(CLBLM_R_X67Y116_SLICE_X100Y116_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f180f5a0f18f)
  ) CLBLM_R_X67Y116_SLICE_X100Y116_DLUT (
.I0(CLBLM_R_X67Y116_SLICE_X101Y116_AQ),
.I1(CLBLM_R_X67Y116_SLICE_X101Y116_A5Q),
.I2(CLBLM_R_X67Y115_SLICE_X100Y115_AQ),
.I3(CLBLM_R_X67Y115_SLICE_X100Y115_A5Q),
.I4(CLBLM_R_X67Y116_SLICE_X100Y116_B5Q),
.I5(CLBLM_R_X67Y116_SLICE_X101Y116_BQ),
.O5(CLBLM_R_X67Y116_SLICE_X100Y116_DO5),
.O6(CLBLM_R_X67Y116_SLICE_X100Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500e4e4e4e4)
  ) CLBLM_R_X67Y116_SLICE_X100Y116_CLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_R_X67Y116_SLICE_X100Y116_AQ),
.I2(CLBLM_R_X67Y116_SLICE_X100Y116_BQ),
.I3(CLBLM_R_X67Y116_SLICE_X101Y116_BQ),
.I4(CLBLM_R_X67Y116_SLICE_X100Y116_DO6),
.I5(1'b1),
.O5(CLBLM_R_X67Y116_SLICE_X100Y116_CO5),
.O6(CLBLM_R_X67Y116_SLICE_X100Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55a0a0eee4eee4)
  ) CLBLM_R_X67Y116_SLICE_X100Y116_BLUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_R_X67Y116_SLICE_X100Y116_BQ),
.I2(CLBLM_R_X67Y115_SLICE_X100Y115_A5Q),
.I3(CLBLM_R_X67Y115_SLICE_X100Y115_AQ),
.I4(CLBLM_R_X67Y116_SLICE_X101Y116_AQ),
.I5(1'b1),
.O5(CLBLM_R_X67Y116_SLICE_X100Y116_BO5),
.O6(CLBLM_R_X67Y116_SLICE_X100Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a3a0a0a0a3a0a)
  ) CLBLM_R_X67Y116_SLICE_X100Y116_ALUT (
.I0(CLBLM_R_X67Y118_SLICE_X100Y118_A5Q),
.I1(CLBLM_R_X67Y116_SLICE_X101Y116_BO6),
.I2(RIOB33_X105Y51_IOB_X1Y51_I),
.I3(CLBLM_R_X67Y116_SLICE_X101Y116_BQ),
.I4(CLBLM_R_X67Y116_SLICE_X100Y116_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X67Y116_SLICE_X100Y116_AO5),
.O6(CLBLM_R_X67Y116_SLICE_X100Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y116_SLICE_X101Y116_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y116_SLICE_X101Y116_AO5),
.Q(CLBLM_R_X67Y116_SLICE_X101Y116_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y116_SLICE_X101Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y116_SLICE_X101Y116_AO6),
.Q(CLBLM_R_X67Y116_SLICE_X101Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y116_SLICE_X101Y116_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y116_SLICE_X100Y116_B5Q),
.Q(CLBLM_R_X67Y116_SLICE_X101Y116_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y116_SLICE_X101Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y116_SLICE_X101Y116_DO5),
.O6(CLBLM_R_X67Y116_SLICE_X101Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y116_SLICE_X101Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y116_SLICE_X101Y116_CO5),
.O6(CLBLM_R_X67Y116_SLICE_X101Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0cfcfc0c0)
  ) CLBLM_R_X67Y116_SLICE_X101Y116_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X67Y115_SLICE_X100Y115_AQ),
.I2(CLBLM_R_X67Y116_SLICE_X101Y116_AQ),
.I3(1'b1),
.I4(CLBLM_R_X67Y115_SLICE_X100Y115_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X67Y116_SLICE_X101Y116_BO5),
.O6(CLBLM_R_X67Y116_SLICE_X101Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddfd88a8fdaadd80)
  ) CLBLM_R_X67Y116_SLICE_X101Y116_ALUT (
.I0(RIOB33_X105Y51_IOB_X1Y51_I),
.I1(CLBLM_R_X67Y115_SLICE_X100Y115_AQ),
.I2(CLBLM_R_X67Y116_SLICE_X101Y116_AQ),
.I3(CLBLM_R_X67Y115_SLICE_X100Y115_A5Q),
.I4(CLBLM_R_X67Y116_SLICE_X101Y116_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X67Y116_SLICE_X101Y116_AO5),
.O6(CLBLM_R_X67Y116_SLICE_X101Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y118_SLICE_X100Y118_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y118_SLICE_X100Y118_AO5),
.Q(CLBLM_R_X67Y118_SLICE_X100Y118_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y118_SLICE_X100Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y118_SLICE_X100Y118_AO6),
.Q(CLBLM_R_X67Y118_SLICE_X100Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y118_SLICE_X100Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y118_SLICE_X100Y118_DO5),
.O6(CLBLM_R_X67Y118_SLICE_X100Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y118_SLICE_X100Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y118_SLICE_X100Y118_CO5),
.O6(CLBLM_R_X67Y118_SLICE_X100Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y118_SLICE_X100Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y118_SLICE_X100Y118_BO5),
.O6(CLBLM_R_X67Y118_SLICE_X100Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h54aa54aafdf0a8f0)
  ) CLBLM_R_X67Y118_SLICE_X100Y118_ALUT (
.I0(CLBLM_R_X67Y118_SLICE_X101Y118_A5Q),
.I1(CLBLM_R_X67Y116_SLICE_X100Y116_CQ),
.I2(CLBLM_R_X67Y118_SLICE_X100Y118_AQ),
.I3(RIOB33_X105Y51_IOB_X1Y51_I),
.I4(CLBLM_R_X67Y118_SLICE_X100Y118_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X67Y118_SLICE_X100Y118_AO5),
.O6(CLBLM_R_X67Y118_SLICE_X100Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y118_SLICE_X101Y118_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y118_SLICE_X101Y118_AO5),
.Q(CLBLM_R_X67Y118_SLICE_X101Y118_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y118_SLICE_X101Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y118_SLICE_X101Y118_AO6),
.Q(CLBLM_R_X67Y118_SLICE_X101Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X67Y118_SLICE_X101Y118_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X67Y118_SLICE_X101Y118_AQ),
.Q(CLBLM_R_X67Y118_SLICE_X101Y118_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y118_SLICE_X101Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y118_SLICE_X101Y118_DO5),
.O6(CLBLM_R_X67Y118_SLICE_X101Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y118_SLICE_X101Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y118_SLICE_X101Y118_CO5),
.O6(CLBLM_R_X67Y118_SLICE_X101Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y118_SLICE_X101Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y118_SLICE_X101Y118_BO5),
.O6(CLBLM_R_X67Y118_SLICE_X101Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ff003030cccc)
  ) CLBLM_R_X67Y118_SLICE_X101Y118_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X67Y118_SLICE_X101Y118_BQ),
.I2(CLBLM_R_X67Y118_SLICE_X101Y118_AQ),
.I3(CLBLM_R_X67Y116_SLICE_X100Y116_CQ),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(1'b1),
.O5(CLBLM_R_X67Y118_SLICE_X101Y118_AO5),
.O6(CLBLM_R_X67Y118_SLICE_X101Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y67_SLICE_X162Y67_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X103Y69_SLICE_X162Y69_AQ),
.Q(CLBLM_R_X103Y67_SLICE_X162Y67_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y67_SLICE_X162Y67_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X103Y67_SLICE_X163Y67_AQ),
.Q(CLBLM_R_X103Y67_SLICE_X162Y67_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y67_SLICE_X162Y67_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X103Y67_SLICE_X162Y67_BQ),
.Q(CLBLM_R_X103Y67_SLICE_X162Y67_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y67_SLICE_X162Y67_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y67_SLICE_X162Y67_DO5),
.O6(CLBLM_R_X103Y67_SLICE_X162Y67_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y67_SLICE_X162Y67_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y67_SLICE_X162Y67_CO5),
.O6(CLBLM_R_X103Y67_SLICE_X162Y67_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y67_SLICE_X162Y67_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y67_SLICE_X162Y67_BO5),
.O6(CLBLM_R_X103Y67_SLICE_X162Y67_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffcfc)
  ) CLBLM_R_X103Y67_SLICE_X162Y67_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X103Y67_SLICE_X162Y67_BQ),
.I2(CLBLM_R_X103Y67_SLICE_X162Y67_CQ),
.I3(1'b1),
.I4(CLBLM_R_X103Y67_SLICE_X162Y67_AQ),
.I5(CLBLM_R_X103Y67_SLICE_X163Y67_BQ),
.O5(CLBLM_R_X103Y67_SLICE_X162Y67_AO5),
.O6(CLBLM_R_X103Y67_SLICE_X162Y67_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y67_SLICE_X163Y67_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X103Y67_SLICE_X162Y67_AQ),
.Q(CLBLM_R_X103Y67_SLICE_X163Y67_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y67_SLICE_X163Y67_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X103Y67_SLICE_X162Y67_CQ),
.Q(CLBLM_R_X103Y67_SLICE_X163Y67_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y67_SLICE_X163Y67_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X103Y67_SLICE_X163Y67_BQ),
.Q(CLBLM_R_X103Y67_SLICE_X163Y67_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y67_SLICE_X163Y67_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y67_SLICE_X163Y67_DO5),
.O6(CLBLM_R_X103Y67_SLICE_X163Y67_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y67_SLICE_X163Y67_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y67_SLICE_X163Y67_CO5),
.O6(CLBLM_R_X103Y67_SLICE_X163Y67_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y67_SLICE_X163Y67_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y67_SLICE_X163Y67_BO5),
.O6(CLBLM_R_X103Y67_SLICE_X163Y67_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y67_SLICE_X163Y67_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y67_SLICE_X163Y67_AO5),
.O6(CLBLM_R_X103Y67_SLICE_X163Y67_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y69_SLICE_X162Y69_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X103Y69_SLICE_X163Y69_AQ),
.Q(CLBLM_R_X103Y69_SLICE_X162Y69_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y69_SLICE_X162Y69_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X103Y69_SLICE_X162Y69_AO6),
.Q(CLBLM_R_X103Y69_SLICE_X162Y69_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y69_SLICE_X162Y69_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y69_SLICE_X162Y69_DO5),
.O6(CLBLM_R_X103Y69_SLICE_X162Y69_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y69_SLICE_X162Y69_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y69_SLICE_X162Y69_CO5),
.O6(CLBLM_R_X103Y69_SLICE_X162Y69_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X103Y69_SLICE_X162Y69_BLUT (
.I0(CLBLM_R_X103Y67_SLICE_X163Y67_AQ),
.I1(CLBLM_R_X103Y67_SLICE_X162Y67_AO6),
.I2(CLBLM_R_X103Y69_SLICE_X162Y69_AQ),
.I3(CLBLM_R_X103Y69_SLICE_X163Y69_AQ),
.I4(CLBLM_R_X103Y67_SLICE_X163Y67_CQ),
.I5(CLBLM_R_X103Y69_SLICE_X162Y69_A5Q),
.O5(CLBLM_R_X103Y69_SLICE_X162Y69_BO5),
.O6(CLBLM_R_X103Y69_SLICE_X162Y69_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33f0f0ffccf0f0)
  ) CLBLM_R_X103Y69_SLICE_X162Y69_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X103Y67_SLICE_X162Y67_CQ),
.I2(CLBLL_R_X83Y94_SLICE_X130Y94_AQ),
.I3(CLBLM_R_X103Y69_SLICE_X162Y69_BO6),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(CLBLM_R_X103Y69_SLICE_X162Y69_A5Q),
.O5(CLBLM_R_X103Y69_SLICE_X162Y69_AO5),
.O6(CLBLM_R_X103Y69_SLICE_X162Y69_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y69_SLICE_X163Y69_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X103Y67_SLICE_X163Y67_CQ),
.Q(CLBLM_R_X103Y69_SLICE_X163Y69_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y69_SLICE_X163Y69_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y69_SLICE_X163Y69_DO5),
.O6(CLBLM_R_X103Y69_SLICE_X163Y69_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y69_SLICE_X163Y69_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y69_SLICE_X163Y69_CO5),
.O6(CLBLM_R_X103Y69_SLICE_X163Y69_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y69_SLICE_X163Y69_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y69_SLICE_X163Y69_BO5),
.O6(CLBLM_R_X103Y69_SLICE_X163Y69_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y69_SLICE_X163Y69_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y69_SLICE_X163Y69_AO5),
.O6(CLBLM_R_X103Y69_SLICE_X163Y69_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y75_SLICE_X162Y75_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X103Y75_SLICE_X163Y75_AQ),
.Q(CLBLM_R_X103Y75_SLICE_X162Y75_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y75_SLICE_X162Y75_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X103Y75_SLICE_X162Y75_AQ),
.Q(CLBLM_R_X103Y75_SLICE_X162Y75_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y75_SLICE_X162Y75_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X103Y75_SLICE_X162Y75_BQ),
.Q(CLBLM_R_X103Y75_SLICE_X162Y75_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y75_SLICE_X162Y75_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y75_SLICE_X162Y75_DO5),
.O6(CLBLM_R_X103Y75_SLICE_X162Y75_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y75_SLICE_X162Y75_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y75_SLICE_X162Y75_CO5),
.O6(CLBLM_R_X103Y75_SLICE_X162Y75_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y75_SLICE_X162Y75_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y75_SLICE_X162Y75_BO5),
.O6(CLBLM_R_X103Y75_SLICE_X162Y75_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffff0)
  ) CLBLM_R_X103Y75_SLICE_X162Y75_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X103Y75_SLICE_X162Y75_AQ),
.I3(CLBLM_R_X103Y75_SLICE_X163Y75_BQ),
.I4(CLBLM_R_X103Y76_SLICE_X162Y76_AQ),
.I5(CLBLM_R_X103Y75_SLICE_X162Y75_CQ),
.O5(CLBLM_R_X103Y75_SLICE_X162Y75_AO5),
.O6(CLBLM_R_X103Y75_SLICE_X162Y75_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y75_SLICE_X163Y75_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X103Y76_SLICE_X162Y76_AQ),
.Q(CLBLM_R_X103Y75_SLICE_X163Y75_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y75_SLICE_X163Y75_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X103Y75_SLICE_X162Y75_CQ),
.Q(CLBLM_R_X103Y75_SLICE_X163Y75_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y75_SLICE_X163Y75_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y75_SLICE_X163Y75_DO5),
.O6(CLBLM_R_X103Y75_SLICE_X163Y75_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y75_SLICE_X163Y75_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y75_SLICE_X163Y75_CO5),
.O6(CLBLM_R_X103Y75_SLICE_X163Y75_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y75_SLICE_X163Y75_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y75_SLICE_X163Y75_BO5),
.O6(CLBLM_R_X103Y75_SLICE_X163Y75_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y75_SLICE_X163Y75_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y75_SLICE_X163Y75_AO5),
.O6(CLBLM_R_X103Y75_SLICE_X163Y75_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y76_SLICE_X162Y76_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLL_R_X79Y104_SLICE_X122Y104_AQ),
.Q(CLBLM_R_X103Y76_SLICE_X162Y76_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y76_SLICE_X162Y76_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X103Y76_SLICE_X163Y76_AQ),
.Q(CLBLM_R_X103Y76_SLICE_X162Y76_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y76_SLICE_X162Y76_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y76_SLICE_X162Y76_DO5),
.O6(CLBLM_R_X103Y76_SLICE_X162Y76_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y76_SLICE_X162Y76_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y76_SLICE_X162Y76_CO5),
.O6(CLBLM_R_X103Y76_SLICE_X162Y76_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y76_SLICE_X162Y76_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y76_SLICE_X162Y76_BO5),
.O6(CLBLM_R_X103Y76_SLICE_X162Y76_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h9999999999999998)
  ) CLBLM_R_X103Y76_SLICE_X162Y76_ALUT (
.I0(CLBLM_R_X103Y75_SLICE_X162Y75_BQ),
.I1(CLBLM_R_X103Y76_SLICE_X162Y76_BQ),
.I2(CLBLL_R_X79Y104_SLICE_X122Y104_AQ),
.I3(CLBLM_R_X103Y75_SLICE_X163Y75_AQ),
.I4(CLBLM_R_X103Y75_SLICE_X162Y75_AO6),
.I5(CLBLM_R_X103Y76_SLICE_X163Y76_AQ),
.O5(CLBLM_R_X103Y76_SLICE_X162Y76_AO5),
.O6(CLBLM_R_X103Y76_SLICE_X162Y76_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y76_SLICE_X163Y76_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.D(CLBLM_R_X103Y75_SLICE_X163Y75_BQ),
.Q(CLBLM_R_X103Y76_SLICE_X163Y76_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y76_SLICE_X163Y76_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y76_SLICE_X163Y76_DO5),
.O6(CLBLM_R_X103Y76_SLICE_X163Y76_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y76_SLICE_X163Y76_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y76_SLICE_X163Y76_CO5),
.O6(CLBLM_R_X103Y76_SLICE_X163Y76_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y76_SLICE_X163Y76_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y76_SLICE_X163Y76_BO5),
.O6(CLBLM_R_X103Y76_SLICE_X163Y76_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y76_SLICE_X163Y76_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y76_SLICE_X163Y76_AO5),
.O6(CLBLM_R_X103Y76_SLICE_X163Y76_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(RIOB33_X105Y77_IOB_X1Y78_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y51_IOB_X0Y51_OBUF (
.I(CLBLM_L_X62Y101_SLICE_X92Y101_AQ),
.O(LIOB33_X0Y51_IOB_X0Y51_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y51_IOB_X0Y52_OBUF (
.I(CLBLM_L_X68Y95_SLICE_X102Y95_A5Q),
.O(LIOB33_X0Y51_IOB_X0Y52_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y53_IOB_X0Y53_OBUF (
.I(CLBLM_L_X62Y90_SLICE_X92Y90_AQ),
.O(LIOB33_X0Y53_IOB_X0Y53_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y53_IOB_X0Y54_OBUF (
.I(CLBLM_L_X62Y92_SLICE_X92Y92_AQ),
.O(LIOB33_X0Y53_IOB_X0Y54_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y55_IOB_X0Y55_OBUF (
.I(CLBLM_L_X60Y97_SLICE_X91Y97_AQ),
.O(LIOB33_X0Y55_IOB_X0Y55_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y55_IOB_X0Y56_OBUF (
.I(CLBLM_L_X62Y92_SLICE_X92Y92_BQ),
.O(LIOB33_X0Y55_IOB_X0Y56_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y57_IOB_X0Y57_OBUF (
.I(CLBLM_L_X62Y95_SLICE_X92Y95_AQ),
.O(LIOB33_X0Y57_IOB_X0Y57_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y57_IOB_X0Y58_OBUF (
.I(CLBLM_L_X72Y107_SLICE_X108Y107_BQ),
.O(LIOB33_X0Y57_IOB_X0Y58_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y59_IOB_X0Y59_OBUF (
.I(CLBLM_L_X60Y101_SLICE_X90Y101_AQ),
.O(LIOB33_X0Y59_IOB_X0Y59_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y59_IOB_X0Y60_OBUF (
.I(CLBLM_L_X72Y106_SLICE_X108Y106_A5Q),
.O(LIOB33_X0Y59_IOB_X0Y60_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y61_IOB_X0Y61_OBUF (
.I(CLBLM_R_X65Y109_SLICE_X98Y109_A5Q),
.O(LIOB33_X0Y61_IOB_X0Y61_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y61_IOB_X0Y62_OBUF (
.I(CLBLM_R_X65Y110_SLICE_X99Y110_B5Q),
.O(LIOB33_X0Y61_IOB_X0Y62_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y63_IOB_X0Y63_OBUF (
.I(CLBLL_R_X73Y102_SLICE_X111Y102_A5Q),
.O(LIOB33_X0Y63_IOB_X0Y63_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y63_IOB_X0Y64_OBUF (
.I(CLBLL_R_X73Y103_SLICE_X111Y103_A5Q),
.O(LIOB33_X0Y63_IOB_X0Y64_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y65_IOB_X0Y65_OBUF (
.I(CLBLM_L_X72Y107_SLICE_X109Y107_BQ),
.O(LIOB33_X0Y65_IOB_X0Y65_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y65_IOB_X0Y66_OBUF (
.I(CLBLM_R_X65Y110_SLICE_X98Y110_A5Q),
.O(LIOB33_X0Y65_IOB_X0Y66_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y67_IOB_X0Y67_OBUF (
.I(CLBLM_L_X72Y103_SLICE_X109Y103_AQ),
.O(LIOB33_X0Y67_IOB_X0Y67_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y67_IOB_X0Y68_OBUF (
.I(CLBLL_R_X71Y134_SLICE_X106Y134_AQ),
.O(LIOB33_X0Y67_IOB_X0Y68_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y69_IOB_X0Y69_OBUF (
.I(CLBLM_L_X60Y92_SLICE_X90Y92_AQ),
.O(LIOB33_X0Y69_IOB_X0Y69_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y69_IOB_X0Y70_OBUF (
.I(CLBLL_R_X75Y127_SLICE_X115Y127_AQ),
.O(LIOB33_X0Y69_IOB_X0Y70_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y71_IOB_X0Y71_OBUF (
.I(CLBLM_L_X60Y94_SLICE_X90Y94_AQ),
.O(LIOB33_X0Y71_IOB_X0Y71_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y71_IOB_X0Y72_OBUF (
.I(CLBLM_L_X60Y104_SLICE_X90Y104_AQ),
.O(LIOB33_X0Y71_IOB_X0Y72_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y73_IOB_X0Y73_OBUF (
.I(CLBLM_L_X62Y105_SLICE_X93Y105_A5Q),
.O(LIOB33_X0Y73_IOB_X0Y73_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y73_IOB_X0Y74_OBUF (
.I(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.O(LIOB33_X0Y73_IOB_X0Y74_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y75_IOB_X0Y75_OBUF (
.I(CLBLM_L_X60Y101_SLICE_X90Y101_BQ),
.O(LIOB33_X0Y75_IOB_X0Y75_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y75_IOB_X0Y76_OBUF (
.I(CLBLM_L_X60Y99_SLICE_X90Y99_AQ),
.O(LIOB33_X0Y75_IOB_X0Y76_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y77_IOB_X0Y77_OBUF (
.I(CLBLM_L_X60Y97_SLICE_X90Y97_BQ),
.O(LIOB33_X0Y77_IOB_X0Y77_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y77_IOB_X0Y78_OBUF (
.I(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.O(LIOB33_X0Y77_IOB_X0Y78_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y79_IOB_X0Y79_OBUF (
.I(CLBLM_L_X64Y106_SLICE_X96Y106_A5Q),
.O(LIOB33_X0Y79_IOB_X0Y79_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y79_IOB_X0Y80_OBUF (
.I(CLBLM_L_X60Y92_SLICE_X90Y92_BQ),
.O(LIOB33_X0Y79_IOB_X0Y80_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y81_IOB_X0Y81_OBUF (
.I(CLBLM_L_X60Y99_SLICE_X90Y99_BQ),
.O(LIOB33_X0Y81_IOB_X0Y81_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y81_IOB_X0Y82_OBUF (
.I(CLBLM_L_X62Y107_SLICE_X93Y107_A5Q),
.O(LIOB33_X0Y81_IOB_X0Y82_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y83_IOB_X0Y83_OBUF (
.I(CLBLM_L_X70Y99_SLICE_X104Y99_AQ),
.O(LIOB33_X0Y83_IOB_X0Y83_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y83_IOB_X0Y84_OBUF (
.I(CLBLM_L_X60Y99_SLICE_X90Y99_CQ),
.O(LIOB33_X0Y83_IOB_X0Y84_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y85_IOB_X0Y85_OBUF (
.I(CLBLM_L_X60Y94_SLICE_X90Y94_BQ),
.O(LIOB33_X0Y85_IOB_X0Y85_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y85_IOB_X0Y86_OBUF (
.I(CLBLM_L_X70Y100_SLICE_X105Y100_CQ),
.O(LIOB33_X0Y85_IOB_X0Y86_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y87_IOB_X0Y87_OBUF (
.I(CLBLM_R_X63Y97_SLICE_X94Y97_B5Q),
.O(LIOB33_X0Y87_IOB_X0Y87_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y87_IOB_X0Y88_OBUF (
.I(CLBLM_L_X60Y94_SLICE_X90Y94_CQ),
.O(LIOB33_X0Y87_IOB_X0Y88_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y89_IOB_X0Y89_OBUF (
.I(CLBLM_R_X63Y98_SLICE_X94Y98_BQ),
.O(LIOB33_X0Y89_IOB_X0Y89_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y89_IOB_X0Y90_OBUF (
.I(CLBLM_R_X63Y103_SLICE_X94Y103_AQ),
.O(LIOB33_X0Y89_IOB_X0Y90_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y91_IOB_X0Y91_OBUF (
.I(CLBLM_L_X60Y99_SLICE_X90Y99_DQ),
.O(LIOB33_X0Y91_IOB_X0Y91_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y91_IOB_X0Y92_OBUF (
.I(CLBLM_L_X62Y95_SLICE_X92Y95_CQ),
.O(LIOB33_X0Y91_IOB_X0Y92_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y93_IOB_X0Y93_OBUF (
.I(CLBLM_L_X62Y95_SLICE_X92Y95_BQ),
.O(LIOB33_X0Y93_IOB_X0Y93_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y93_IOB_X0Y94_OBUF (
.I(CLBLM_L_X62Y106_SLICE_X92Y106_AQ),
.O(LIOB33_X0Y93_IOB_X0Y94_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y95_IOB_X0Y95_OBUF (
.I(CLBLM_L_X70Y101_SLICE_X104Y101_AQ),
.O(LIOB33_X0Y95_IOB_X0Y95_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y95_IOB_X0Y96_OBUF (
.I(CLBLM_R_X63Y97_SLICE_X95Y97_AQ),
.O(LIOB33_X0Y95_IOB_X0Y96_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y97_IOB_X0Y97_OBUF (
.I(CLBLM_L_X62Y103_SLICE_X92Y103_A5Q),
.O(LIOB33_X0Y97_IOB_X0Y97_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y97_IOB_X0Y98_OBUF (
.I(CLBLM_L_X68Y97_SLICE_X103Y97_AQ),
.O(LIOB33_X0Y97_IOB_X0Y98_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y101_OBUF (
.I(RIOB33_X105Y57_IOB_X1Y58_I),
.O(LIOB33_X0Y101_IOB_X0Y101_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y102_OBUF (
.I(RIOB33_X105Y59_IOB_X1Y59_I),
.O(LIOB33_X0Y101_IOB_X0Y102_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y103_OBUF (
.I(RIOB33_X105Y55_IOB_X1Y56_I),
.O(LIOB33_X0Y103_IOB_X0Y103_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y104_OBUF (
.I(RIOB33_X105Y53_IOB_X1Y53_I),
.O(LIOB33_X0Y103_IOB_X0Y104_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y105_OBUF (
.I(RIOB33_X105Y53_IOB_X1Y54_I),
.O(LIOB33_X0Y105_IOB_X0Y105_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y106_OBUF (
.I(RIOB33_X105Y59_IOB_X1Y60_I),
.O(LIOB33_X0Y105_IOB_X0Y106_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y107_OBUF (
.I(RIOB33_X105Y55_IOB_X1Y55_I),
.O(LIOB33_X0Y107_IOB_X0Y107_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y108_OBUF (
.I(CLBLM_L_X70Y110_SLICE_X104Y110_CQ),
.O(LIOB33_X0Y107_IOB_X0Y108_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y109_OBUF (
.I(CLBLL_R_X75Y133_SLICE_X114Y133_AQ),
.O(LIOB33_X0Y109_IOB_X0Y109_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y110_OBUF (
.I(CLBLL_R_X77Y129_SLICE_X118Y129_AQ),
.O(LIOB33_X0Y109_IOB_X0Y110_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y111_OBUF (
.I(CLBLM_R_X65Y106_SLICE_X99Y106_DQ),
.O(LIOB33_X0Y111_IOB_X0Y111_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y112_OBUF (
.I(CLBLM_L_X64Y99_SLICE_X97Y99_B5Q),
.O(LIOB33_X0Y111_IOB_X0Y112_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y113_OBUF (
.I(CLBLM_R_X63Y122_SLICE_X95Y122_CQ),
.O(LIOB33_X0Y113_IOB_X0Y113_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y114_OBUF (
.I(CLBLL_R_X71Y124_SLICE_X106Y124_AQ),
.O(LIOB33_X0Y113_IOB_X0Y114_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y115_OBUF (
.I(CLBLM_R_X67Y118_SLICE_X100Y118_A5Q),
.O(LIOB33_X0Y115_IOB_X0Y115_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y116_OBUF (
.I(CLBLM_L_X76Y118_SLICE_X117Y118_CQ),
.O(LIOB33_X0Y115_IOB_X0Y116_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y117_OBUF (
.I(CLBLM_L_X76Y125_SLICE_X116Y125_AQ),
.O(LIOB33_X0Y117_IOB_X0Y117_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y118_OBUF (
.I(CLBLM_R_X67Y116_SLICE_X100Y116_AQ),
.O(LIOB33_X0Y117_IOB_X0Y118_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y119_OBUF (
.I(CLBLM_R_X63Y106_SLICE_X95Y106_AQ),
.O(LIOB33_X0Y119_IOB_X0Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y120_OBUF (
.I(CLBLL_R_X71Y119_SLICE_X106Y119_AQ),
.O(LIOB33_X0Y119_IOB_X0Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y121_OBUF (
.I(CLBLL_R_X73Y123_SLICE_X110Y123_AQ),
.O(LIOB33_X0Y121_IOB_X0Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y122_OBUF (
.I(RIOB33_X105Y51_IOB_X1Y52_I),
.O(LIOB33_X0Y121_IOB_X0Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y123_OBUF (
.I(CLBLM_R_X67Y108_SLICE_X100Y108_AO6),
.O(LIOB33_X0Y123_IOB_X0Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y124_OBUF (
.I(CLBLL_L_X34Y123_SLICE_X50Y123_AO6),
.O(LIOB33_X0Y123_IOB_X0Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y125_OBUF (
.I(1'b1),
.O(LIOB33_X0Y125_IOB_X0Y125_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y126_OBUF (
.I(CLBLL_L_X2Y131_SLICE_X0Y131_AO6),
.O(LIOB33_X0Y125_IOB_X0Y126_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y127_OBUF (
.I(CLBLL_L_X34Y126_SLICE_X50Y126_AO6),
.O(LIOB33_X0Y127_IOB_X0Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y128_OBUF (
.I(CLBLL_R_X73Y131_SLICE_X110Y131_AQ),
.O(LIOB33_X0Y127_IOB_X0Y128_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y129_OBUF (
.I(CLBLL_L_X34Y128_SLICE_X50Y128_AO6),
.O(LIOB33_X0Y129_IOB_X0Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y130_OBUF (
.I(1'b1),
.O(LIOB33_X0Y129_IOB_X0Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y131_OBUF (
.I(CLBLM_L_X62Y107_SLICE_X92Y107_AO5),
.O(LIOB33_X0Y131_IOB_X0Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y132_OBUF (
.I(CLBLM_L_X70Y134_SLICE_X104Y134_CO5),
.O(LIOB33_X0Y131_IOB_X0Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y133_OBUF (
.I(CLBLM_R_X63Y105_SLICE_X95Y105_A5Q),
.O(LIOB33_X0Y133_IOB_X0Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y134_OBUF (
.I(CLBLM_L_X70Y135_SLICE_X104Y135_CO6),
.O(LIOB33_X0Y133_IOB_X0Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y135_OBUF (
.I(1'b1),
.O(LIOB33_X0Y135_IOB_X0Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y136_OBUF (
.I(1'b1),
.O(LIOB33_X0Y135_IOB_X0Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y137_OBUF (
.I(1'b1),
.O(LIOB33_X0Y137_IOB_X0Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y138_OBUF (
.I(1'b1),
.O(LIOB33_X0Y137_IOB_X0Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y139_OBUF (
.I(1'b1),
.O(LIOB33_X0Y139_IOB_X0Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y140_OBUF (
.I(1'b1),
.O(LIOB33_X0Y139_IOB_X0Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y141_OBUF (
.I(1'b1),
.O(LIOB33_X0Y141_IOB_X0Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y142_OBUF (
.I(1'b1),
.O(LIOB33_X0Y141_IOB_X0Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y143_IOB_X0Y143_OBUF (
.I(1'b1),
.O(LIOB33_X0Y143_IOB_X0Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y145_OBUF (
.I(CLBLL_R_X71Y130_SLICE_X106Y130_DO6),
.O(LIOB33_X0Y145_IOB_X0Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y146_OBUF (
.I(CLBLM_L_X72Y123_SLICE_X108Y123_BO6),
.O(LIOB33_X0Y145_IOB_X0Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y147_OBUF (
.I(CLBLL_R_X71Y124_SLICE_X106Y124_BO6),
.O(LIOB33_X0Y147_IOB_X0Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y148_OBUF (
.I(CLBLL_R_X73Y134_SLICE_X110Y134_AO5),
.O(LIOB33_X0Y147_IOB_X0Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y151_OBUF (
.I(CLBLM_L_X72Y128_SLICE_X109Y128_AO6),
.O(LIOB33_X0Y151_IOB_X0Y151_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y152_OBUF (
.I(CLBLM_L_X64Y105_SLICE_X97Y105_DO6),
.O(LIOB33_X0Y151_IOB_X0Y152_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y153_IOB_X0Y153_OBUF (
.I(CLBLM_R_X65Y106_SLICE_X99Y106_DQ),
.O(LIOB33_X0Y153_IOB_X0Y153_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y153_IOB_X0Y154_OBUF (
.I(CLBLM_R_X67Y118_SLICE_X100Y118_A5Q),
.O(LIOB33_X0Y153_IOB_X0Y154_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y155_IOB_X0Y155_OBUF (
.I(CLBLM_L_X76Y118_SLICE_X117Y118_CQ),
.O(LIOB33_X0Y155_IOB_X0Y155_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y155_IOB_X0Y156_OBUF (
.I(CLBLM_L_X64Y99_SLICE_X97Y99_B5Q),
.O(LIOB33_X0Y155_IOB_X0Y156_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y157_IOB_X0Y157_OBUF (
.I(CLBLM_R_X63Y122_SLICE_X95Y122_CQ),
.O(LIOB33_X0Y157_IOB_X0Y157_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y157_IOB_X0Y158_OBUF (
.I(CLBLM_L_X76Y125_SLICE_X116Y125_AQ),
.O(LIOB33_X0Y157_IOB_X0Y158_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y159_IOB_X0Y159_OBUF (
.I(CLBLM_R_X67Y116_SLICE_X100Y116_AQ),
.O(LIOB33_X0Y159_IOB_X0Y159_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y159_IOB_X0Y160_OBUF (
.I(CLBLL_R_X71Y119_SLICE_X106Y119_AQ),
.O(LIOB33_X0Y159_IOB_X0Y160_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y161_IOB_X0Y161_OBUF (
.I(CLBLM_L_X70Y110_SLICE_X104Y110_CQ),
.O(LIOB33_X0Y161_IOB_X0Y161_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y161_IOB_X0Y162_OBUF (
.I(CLBLL_R_X71Y124_SLICE_X106Y124_AQ),
.O(LIOB33_X0Y161_IOB_X0Y162_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y163_IOB_X0Y163_OBUF (
.I(CLBLM_R_X63Y106_SLICE_X95Y106_AQ),
.O(LIOB33_X0Y163_IOB_X0Y163_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y163_IOB_X0Y164_OBUF (
.I(CLBLL_R_X73Y123_SLICE_X110Y123_AQ),
.O(LIOB33_X0Y163_IOB_X0Y164_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y165_IOB_X0Y165_OBUF (
.I(CLBLL_L_X34Y123_SLICE_X50Y123_AO6),
.O(LIOB33_X0Y165_IOB_X0Y165_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y165_IOB_X0Y166_OBUF (
.I(CLBLL_L_X2Y131_SLICE_X0Y131_AO6),
.O(LIOB33_X0Y165_IOB_X0Y166_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y167_IOB_X0Y167_OBUF (
.I(CLBLL_L_X34Y126_SLICE_X50Y126_AO6),
.O(LIOB33_X0Y167_IOB_X0Y167_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y167_IOB_X0Y168_OBUF (
.I(CLBLL_L_X34Y128_SLICE_X50Y128_AO6),
.O(LIOB33_X0Y167_IOB_X0Y168_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y169_IOB_X0Y169_OBUF (
.I(CLBLL_R_X73Y131_SLICE_X110Y131_AQ),
.O(LIOB33_X0Y169_IOB_X0Y169_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y169_IOB_X0Y170_OBUF (
.I(CLBLM_L_X74Y120_SLICE_X112Y120_AO6),
.O(LIOB33_X0Y169_IOB_X0Y170_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y171_IOB_X0Y171_OBUF (
.I(1'b1),
.O(LIOB33_X0Y171_IOB_X0Y171_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y171_IOB_X0Y172_OBUF (
.I(1'b1),
.O(LIOB33_X0Y171_IOB_X0Y172_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y173_IOB_X0Y173_OBUF (
.I(CLBLM_L_X68Y107_SLICE_X102Y107_BO6),
.O(LIOB33_X0Y173_IOB_X0Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y173_IOB_X0Y174_OBUF (
.I(CLBLM_L_X62Y107_SLICE_X92Y107_AO5),
.O(LIOB33_X0Y173_IOB_X0Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y175_IOB_X0Y175_OBUF (
.I(CLBLM_R_X63Y105_SLICE_X95Y105_A5Q),
.O(LIOB33_X0Y175_IOB_X0Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y175_IOB_X0Y176_OBUF (
.I(CLBLM_L_X70Y135_SLICE_X104Y135_CO6),
.O(LIOB33_X0Y175_IOB_X0Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y177_OBUF (
.I(CLBLM_L_X70Y134_SLICE_X104Y134_CO5),
.O(LIOB33_X0Y177_IOB_X0Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y178_OBUF (
.I(CLBLM_L_X72Y122_SLICE_X108Y122_AO6),
.O(LIOB33_X0Y177_IOB_X0Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y179_OBUF (
.I(1'b1),
.O(LIOB33_X0Y179_IOB_X0Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y180_OBUF (
.I(1'b1),
.O(LIOB33_X0Y179_IOB_X0Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y181_OBUF (
.I(CLBLM_L_X64Y106_SLICE_X97Y106_AO6),
.O(LIOB33_X0Y181_IOB_X0Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y182_OBUF (
.I(CLBLM_L_X70Y126_SLICE_X104Y126_DO6),
.O(LIOB33_X0Y181_IOB_X0Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y183_OBUF (
.I(CLBLM_L_X70Y125_SLICE_X104Y125_DO6),
.O(LIOB33_X0Y183_IOB_X0Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y184_OBUF (
.I(CLBLL_R_X73Y134_SLICE_X110Y134_AO5),
.O(LIOB33_X0Y183_IOB_X0Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y185_OBUF (
.I(1'b1),
.O(LIOB33_X0Y185_IOB_X0Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y186_OBUF (
.I(1'b1),
.O(LIOB33_X0Y185_IOB_X0Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y187_OBUF (
.I(1'b1),
.O(LIOB33_X0Y187_IOB_X0Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y188_OBUF (
.I(CLBLL_R_X77Y124_SLICE_X118Y124_AO6),
.O(LIOB33_X0Y187_IOB_X0Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y189_OBUF (
.I(1'b1),
.O(LIOB33_X0Y189_IOB_X0Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y190_OBUF (
.I(1'b1),
.O(LIOB33_X0Y189_IOB_X0Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y191_OBUF (
.I(1'b1),
.O(LIOB33_X0Y191_IOB_X0Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y192_OBUF (
.I(1'b1),
.O(LIOB33_X0Y191_IOB_X0Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y193_OBUF (
.I(1'b1),
.O(LIOB33_X0Y193_IOB_X0Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y194_OBUF (
.I(1'b1),
.O(LIOB33_X0Y193_IOB_X0Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y195_OBUF (
.I(1'b1),
.O(LIOB33_X0Y195_IOB_X0Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y196_OBUF (
.I(CLBLM_L_X64Y105_SLICE_X97Y105_DO6),
.O(LIOB33_X0Y195_IOB_X0Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y197_OBUF (
.I(1'b1),
.O(LIOB33_X0Y197_IOB_X0Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y198_OBUF (
.I(1'b1),
.O(LIOB33_X0Y197_IOB_X0Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y50_IOB_X0Y50_OBUF (
.I(CLBLM_L_X60Y97_SLICE_X90Y97_DQ),
.O(LIOB33_SING_X0Y50_IOB_X0Y50_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y99_IOB_X0Y99_OBUF (
.I(RIOB33_X105Y61_IOB_X1Y62_I),
.O(LIOB33_SING_X0Y99_IOB_X0Y99_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y100_IOB_X0Y100_OBUF (
.I(RIOB33_X105Y57_IOB_X1Y57_I),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y149_IOB_X0Y149_OBUF (
.I(CLBLM_R_X67Y105_SLICE_X101Y105_AO6),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y150_IOB_X0Y150_OBUF (
.I(CLBLM_L_X74Y129_SLICE_X113Y129_BO6),
.O(LIOB33_SING_X0Y150_IOB_X0Y150_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y199_IOB_X0Y199_OBUF (
.I(1'b1),
.O(LIOB33_SING_X0Y199_IOB_X0Y199_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y51_IOB_X1Y51_IBUF (
.I(RIOB33_X105Y51_IOB_X1Y51_IPAD),
.O(RIOB33_X105Y51_IOB_X1Y51_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y51_IOB_X1Y52_IBUF (
.I(RIOB33_X105Y51_IOB_X1Y52_IPAD),
.O(RIOB33_X105Y51_IOB_X1Y52_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y53_IOB_X1Y53_IBUF (
.I(RIOB33_X105Y53_IOB_X1Y53_IPAD),
.O(RIOB33_X105Y53_IOB_X1Y53_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y53_IOB_X1Y54_IBUF (
.I(RIOB33_X105Y53_IOB_X1Y54_IPAD),
.O(RIOB33_X105Y53_IOB_X1Y54_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y55_IOB_X1Y55_IBUF (
.I(RIOB33_X105Y55_IOB_X1Y55_IPAD),
.O(RIOB33_X105Y55_IOB_X1Y55_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y55_IOB_X1Y56_IBUF (
.I(RIOB33_X105Y55_IOB_X1Y56_IPAD),
.O(RIOB33_X105Y55_IOB_X1Y56_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y57_IOB_X1Y57_IBUF (
.I(RIOB33_X105Y57_IOB_X1Y57_IPAD),
.O(RIOB33_X105Y57_IOB_X1Y57_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y57_IOB_X1Y58_IBUF (
.I(RIOB33_X105Y57_IOB_X1Y58_IPAD),
.O(RIOB33_X105Y57_IOB_X1Y58_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y59_IOB_X1Y59_IBUF (
.I(RIOB33_X105Y59_IOB_X1Y59_IPAD),
.O(RIOB33_X105Y59_IOB_X1Y59_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y59_IOB_X1Y60_IBUF (
.I(RIOB33_X105Y59_IOB_X1Y60_IPAD),
.O(RIOB33_X105Y59_IOB_X1Y60_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y61_IOB_X1Y61_IBUF (
.I(RIOB33_X105Y61_IOB_X1Y61_IPAD),
.O(RIOB33_X105Y61_IOB_X1Y61_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y61_IOB_X1Y62_IBUF (
.I(RIOB33_X105Y61_IOB_X1Y62_IPAD),
.O(RIOB33_X105Y61_IOB_X1Y62_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y63_IOB_X1Y63_OBUF (
.I(CLBLM_R_X103Y67_SLICE_X162Y67_AQ),
.O(RIOB33_X105Y63_IOB_X1Y63_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y63_IOB_X1Y64_OBUF (
.I(CLBLM_R_X103Y67_SLICE_X163Y67_AQ),
.O(RIOB33_X105Y63_IOB_X1Y64_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y65_IOB_X1Y65_OBUF (
.I(CLBLM_R_X103Y67_SLICE_X162Y67_BQ),
.O(RIOB33_X105Y65_IOB_X1Y65_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y65_IOB_X1Y66_OBUF (
.I(CLBLM_R_X103Y67_SLICE_X162Y67_CQ),
.O(RIOB33_X105Y65_IOB_X1Y66_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y67_IOB_X1Y67_OBUF (
.I(CLBLM_R_X103Y67_SLICE_X163Y67_BQ),
.O(RIOB33_X105Y67_IOB_X1Y67_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y67_IOB_X1Y68_OBUF (
.I(CLBLM_R_X103Y67_SLICE_X163Y67_CQ),
.O(RIOB33_X105Y67_IOB_X1Y68_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y69_IOB_X1Y69_OBUF (
.I(CLBLM_R_X103Y69_SLICE_X163Y69_AQ),
.O(RIOB33_X105Y69_IOB_X1Y69_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y69_IOB_X1Y70_OBUF (
.I(CLBLM_L_X82Y98_SLICE_X128Y98_AQ),
.O(RIOB33_X105Y69_IOB_X1Y70_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y71_IOB_X1Y71_OBUF (
.I(CLBLM_R_X103Y75_SLICE_X162Y75_BQ),
.O(RIOB33_X105Y71_IOB_X1Y71_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y71_IOB_X1Y72_OBUF (
.I(CLBLM_R_X103Y76_SLICE_X162Y76_AQ),
.O(RIOB33_X105Y71_IOB_X1Y72_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y73_IOB_X1Y73_OBUF (
.I(CLBLM_R_X103Y75_SLICE_X163Y75_AQ),
.O(RIOB33_X105Y73_IOB_X1Y73_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y73_IOB_X1Y74_OBUF (
.I(CLBLM_R_X103Y75_SLICE_X162Y75_AQ),
.O(RIOB33_X105Y73_IOB_X1Y74_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y75_IOB_X1Y75_OBUF (
.I(CLBLM_R_X103Y75_SLICE_X162Y75_CQ),
.O(RIOB33_X105Y75_IOB_X1Y75_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y75_IOB_X1Y76_OBUF (
.I(CLBLM_R_X103Y75_SLICE_X163Y75_BQ),
.O(RIOB33_X105Y75_IOB_X1Y76_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y77_IOB_X1Y77_OBUF (
.I(CLBLM_R_X103Y76_SLICE_X163Y76_AQ),
.O(RIOB33_X105Y77_IOB_X1Y77_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y77_IOB_X1Y78_IBUF (
.I(RIOB33_X105Y77_IOB_X1Y78_IPAD),
.O(RIOB33_X105Y77_IOB_X1Y78_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y79_IOB_X1Y79_OBUF (
.I(CLBLL_R_X83Y94_SLICE_X130Y94_A5Q),
.O(RIOB33_X105Y79_IOB_X1Y79_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y79_IOB_X1Y80_OBUF (
.I(1'b0),
.O(RIOB33_X105Y79_IOB_X1Y80_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y81_IOB_X1Y81_OBUF (
.I(CLBLL_R_X71Y110_SLICE_X106Y110_A5Q),
.O(RIOB33_X105Y81_IOB_X1Y81_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y81_IOB_X1Y82_OBUF (
.I(CLBLL_R_X77Y104_SLICE_X119Y104_A5Q),
.O(RIOB33_X105Y81_IOB_X1Y82_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y83_IOB_X1Y83_OBUF (
.I(CLBLM_R_X63Y105_SLICE_X95Y105_AQ),
.O(RIOB33_X105Y83_IOB_X1Y83_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y83_IOB_X1Y84_OBUF (
.I(CLBLM_L_X72Y118_SLICE_X108Y118_D5Q),
.O(RIOB33_X105Y83_IOB_X1Y84_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y85_IOB_X1Y85_OBUF (
.I(CLBLL_R_X71Y98_SLICE_X106Y98_AQ),
.O(RIOB33_X105Y85_IOB_X1Y85_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y85_IOB_X1Y86_OBUF (
.I(CLBLM_L_X64Y99_SLICE_X97Y99_A5Q),
.O(RIOB33_X105Y85_IOB_X1Y86_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y87_IOB_X1Y87_OBUF (
.I(CLBLM_L_X64Y97_SLICE_X97Y97_AQ),
.O(RIOB33_X105Y87_IOB_X1Y87_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y87_IOB_X1Y88_OBUF (
.I(CLBLM_L_X68Y105_SLICE_X102Y105_AQ),
.O(RIOB33_X105Y87_IOB_X1Y88_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y89_IOB_X1Y89_OBUF (
.I(CLBLM_L_X64Y101_SLICE_X96Y101_AQ),
.O(RIOB33_X105Y89_IOB_X1Y89_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y89_IOB_X1Y90_OBUF (
.I(CLBLM_L_X72Y119_SLICE_X108Y119_C5Q),
.O(RIOB33_X105Y89_IOB_X1Y90_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y91_IOB_X1Y91_OBUF (
.I(CLBLM_L_X68Y98_SLICE_X103Y98_AQ),
.O(RIOB33_X105Y91_IOB_X1Y91_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y101_IOB_X1Y101_OBUF (
.I(CLBLM_L_X72Y109_SLICE_X109Y109_DQ),
.O(RIOB33_X105Y101_IOB_X1Y101_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y101_IOB_X1Y102_OBUF (
.I(CLBLL_R_X73Y131_SLICE_X111Y131_AQ),
.O(RIOB33_X105Y101_IOB_X1Y102_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y103_IOB_X1Y103_OBUF (
.I(CLBLL_R_X77Y128_SLICE_X119Y128_DQ),
.O(RIOB33_X105Y103_IOB_X1Y103_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y103_IOB_X1Y104_OBUF (
.I(CLBLM_L_X72Y106_SLICE_X108Y106_AQ),
.O(RIOB33_X105Y103_IOB_X1Y104_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y105_IOB_X1Y105_OBUF (
.I(CLBLM_R_X65Y111_SLICE_X98Y111_AQ),
.O(RIOB33_X105Y105_IOB_X1Y105_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y105_IOB_X1Y106_OBUF (
.I(CLBLL_R_X75Y103_SLICE_X115Y103_AQ),
.O(RIOB33_X105Y105_IOB_X1Y106_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y107_IOB_X1Y107_OBUF (
.I(CLBLM_R_X103Y69_SLICE_X162Y69_AQ),
.O(RIOB33_X105Y107_IOB_X1Y107_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y107_IOB_X1Y108_OBUF (
.I(CLBLL_R_X77Y113_SLICE_X118Y113_AQ),
.O(RIOB33_X105Y107_IOB_X1Y108_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y109_IOB_X1Y109_OBUF (
.I(CLBLL_R_X79Y104_SLICE_X122Y104_AQ),
.O(RIOB33_X105Y109_IOB_X1Y109_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y109_IOB_X1Y110_OBUF (
.I(CLBLM_L_X72Y111_SLICE_X108Y111_C5Q),
.O(RIOB33_X105Y109_IOB_X1Y110_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y111_IOB_X1Y111_OBUF (
.I(CLBLM_L_X62Y107_SLICE_X93Y107_BQ),
.O(RIOB33_X105Y111_IOB_X1Y111_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y111_IOB_X1Y112_OBUF (
.I(CLBLL_R_X71Y100_SLICE_X106Y100_BQ),
.O(RIOB33_X105Y111_IOB_X1Y112_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y113_IOB_X1Y113_OBUF (
.I(CLBLM_L_X62Y99_SLICE_X93Y99_AQ),
.O(RIOB33_X105Y113_IOB_X1Y113_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y113_IOB_X1Y114_OBUF (
.I(1'b0),
.O(RIOB33_X105Y113_IOB_X1Y114_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y115_IOB_X1Y115_OBUF (
.I(CLBLM_L_X62Y100_SLICE_X92Y100_AQ),
.O(RIOB33_X105Y115_IOB_X1Y115_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y115_IOB_X1Y116_OBUF (
.I(CLBLM_L_X68Y95_SLICE_X102Y95_AQ),
.O(RIOB33_X105Y115_IOB_X1Y116_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y117_IOB_X1Y117_OBUF (
.I(CLBLL_R_X73Y118_SLICE_X111Y118_AQ),
.O(RIOB33_X105Y117_IOB_X1Y117_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y117_IOB_X1Y118_OBUF (
.I(CLBLM_L_X70Y136_SLICE_X105Y136_A5Q),
.O(RIOB33_X105Y117_IOB_X1Y118_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y119_IOB_X1Y119_OBUF (
.I(CLBLM_L_X76Y128_SLICE_X116Y128_CQ),
.O(RIOB33_X105Y119_IOB_X1Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y119_IOB_X1Y120_OBUF (
.I(CLBLM_L_X62Y106_SLICE_X93Y106_AQ),
.O(RIOB33_X105Y119_IOB_X1Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y121_IOB_X1Y121_OBUF (
.I(CLBLM_L_X70Y100_SLICE_X104Y100_A5Q),
.O(RIOB33_X105Y121_IOB_X1Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y121_IOB_X1Y122_OBUF (
.I(CLBLM_R_X63Y98_SLICE_X94Y98_AQ),
.O(RIOB33_X105Y121_IOB_X1Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y123_IOB_X1Y123_OBUF (
.I(CLBLM_R_X63Y101_SLICE_X94Y101_AQ),
.O(RIOB33_X105Y123_IOB_X1Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y123_IOB_X1Y124_OBUF (
.I(CLBLM_L_X68Y99_SLICE_X102Y99_AQ),
.O(RIOB33_X105Y123_IOB_X1Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y125_IOB_X1Y125_OBUF (
.I(CLBLM_L_X74Y129_SLICE_X112Y129_BQ),
.O(RIOB33_X105Y125_IOB_X1Y125_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y125_IOB_X1Y126_OBUF (
.I(CLBLM_L_X76Y127_SLICE_X116Y127_AQ),
.O(RIOB33_X105Y125_IOB_X1Y126_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y127_IOB_X1Y127_OBUF (
.I(CLBLM_L_X72Y107_SLICE_X108Y107_A5Q),
.O(RIOB33_X105Y127_IOB_X1Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y127_IOB_X1Y128_OBUF (
.I(CLBLM_R_X65Y110_SLICE_X99Y110_CQ),
.O(RIOB33_X105Y127_IOB_X1Y128_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y129_IOB_X1Y129_OBUF (
.I(CLBLM_L_X78Y106_SLICE_X120Y106_AQ),
.O(RIOB33_X105Y129_IOB_X1Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y129_IOB_X1Y130_OBUF (
.I(CLBLL_R_X73Y103_SLICE_X110Y103_B5Q),
.O(RIOB33_X105Y129_IOB_X1Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y131_IOB_X1Y131_OBUF (
.I(CLBLM_L_X76Y111_SLICE_X116Y111_AQ),
.O(RIOB33_X105Y131_IOB_X1Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y131_IOB_X1Y132_OBUF (
.I(CLBLL_R_X79Y104_SLICE_X122Y104_A5Q),
.O(RIOB33_X105Y131_IOB_X1Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y133_IOB_X1Y133_OBUF (
.I(CLBLL_R_X83Y130_SLICE_X130Y130_AQ),
.O(RIOB33_X105Y133_IOB_X1Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y133_IOB_X1Y134_OBUF (
.I(CLBLL_R_X83Y130_SLICE_X130Y130_BQ),
.O(RIOB33_X105Y133_IOB_X1Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y135_IOB_X1Y135_OBUF (
.I(CLBLL_R_X83Y130_SLICE_X130Y130_CQ),
.O(RIOB33_X105Y135_IOB_X1Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y135_IOB_X1Y136_OBUF (
.I(CLBLL_R_X83Y130_SLICE_X130Y130_DQ),
.O(RIOB33_X105Y135_IOB_X1Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y137_IOB_X1Y137_OBUF (
.I(CLBLL_R_X77Y125_SLICE_X118Y125_AQ),
.O(RIOB33_X105Y137_IOB_X1Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y137_IOB_X1Y138_OBUF (
.I(CLBLM_L_X82Y130_SLICE_X128Y130_AQ),
.O(RIOB33_X105Y137_IOB_X1Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y139_IOB_X1Y139_OBUF (
.I(CLBLL_R_X83Y132_SLICE_X130Y132_AQ),
.O(RIOB33_X105Y139_IOB_X1Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y139_IOB_X1Y140_OBUF (
.I(CLBLM_L_X72Y107_SLICE_X109Y107_A5Q),
.O(RIOB33_X105Y139_IOB_X1Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y141_IOB_X1Y141_OBUF (
.I(CLBLM_R_X65Y110_SLICE_X99Y110_AQ),
.O(RIOB33_X105Y141_IOB_X1Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y141_IOB_X1Y142_OBUF (
.I(CLBLL_R_X73Y103_SLICE_X110Y103_A5Q),
.O(RIOB33_X105Y141_IOB_X1Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y143_IOB_X1Y143_OBUF (
.I(CLBLM_L_X62Y106_SLICE_X92Y106_BQ),
.O(RIOB33_X105Y143_IOB_X1Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y143_IOB_X1Y144_OBUF (
.I(CLBLM_L_X70Y101_SLICE_X105Y101_AQ),
.O(RIOB33_X105Y143_IOB_X1Y144_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y145_IOB_X1Y145_OBUF (
.I(CLBLL_R_X75Y107_SLICE_X114Y107_AQ),
.O(RIOB33_X105Y145_IOB_X1Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y145_IOB_X1Y146_OBUF (
.I(CLBLM_R_X63Y97_SLICE_X94Y97_AQ),
.O(RIOB33_X105Y145_IOB_X1Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y147_IOB_X1Y147_OBUF (
.I(CLBLL_R_X77Y108_SLICE_X118Y108_AQ),
.O(RIOB33_X105Y147_IOB_X1Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y147_IOB_X1Y148_OBUF (
.I(CLBLM_L_X62Y103_SLICE_X92Y103_B5Q),
.O(RIOB33_X105Y147_IOB_X1Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y151_OBUF (
.I(1'b1),
.O(RIOB33_X105Y151_IOB_X1Y151_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y152_OBUF (
.I(1'b1),
.O(RIOB33_X105Y151_IOB_X1Y152_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y153_OBUF (
.I(1'b1),
.O(RIOB33_X105Y153_IOB_X1Y153_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y154_OBUF (
.I(1'b1),
.O(RIOB33_X105Y153_IOB_X1Y154_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y155_OBUF (
.I(1'b1),
.O(RIOB33_X105Y155_IOB_X1Y155_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y156_OBUF (
.I(1'b1),
.O(RIOB33_X105Y155_IOB_X1Y156_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y157_OBUF (
.I(1'b1),
.O(RIOB33_X105Y157_IOB_X1Y157_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y158_OBUF (
.I(1'b1),
.O(RIOB33_X105Y157_IOB_X1Y158_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y159_OBUF (
.I(1'b1),
.O(RIOB33_X105Y159_IOB_X1Y159_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y160_OBUF (
.I(CLBLM_L_X74Y120_SLICE_X112Y120_AO6),
.O(RIOB33_X105Y159_IOB_X1Y160_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y161_OBUF (
.I(1'b1),
.O(RIOB33_X105Y161_IOB_X1Y161_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y162_OBUF (
.I(1'b1),
.O(RIOB33_X105Y161_IOB_X1Y162_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y163_OBUF (
.I(1'b0),
.O(RIOB33_X105Y163_IOB_X1Y163_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y164_OBUF (
.I(CLBLL_R_X77Y124_SLICE_X118Y124_AO6),
.O(RIOB33_X105Y163_IOB_X1Y164_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y165_OBUF (
.I(CLBLM_L_X70Y111_SLICE_X105Y111_DO6),
.O(RIOB33_X105Y165_IOB_X1Y165_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y166_OBUF (
.I(1'b1),
.O(RIOB33_X105Y165_IOB_X1Y166_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y167_OBUF (
.I(1'b1),
.O(RIOB33_X105Y167_IOB_X1Y167_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y168_OBUF (
.I(1'b1),
.O(RIOB33_X105Y167_IOB_X1Y168_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y169_OBUF (
.I(1'b1),
.O(RIOB33_X105Y169_IOB_X1Y169_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y170_OBUF (
.I(1'b1),
.O(RIOB33_X105Y169_IOB_X1Y170_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y171_OBUF (
.I(1'b1),
.O(RIOB33_X105Y171_IOB_X1Y171_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y172_OBUF (
.I(1'b1),
.O(RIOB33_X105Y171_IOB_X1Y172_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y173_OBUF (
.I(1'b1),
.O(RIOB33_X105Y173_IOB_X1Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y174_OBUF (
.I(CLBLM_L_X70Y111_SLICE_X105Y111_DO6),
.O(RIOB33_X105Y173_IOB_X1Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y175_OBUF (
.I(1'b1),
.O(RIOB33_X105Y175_IOB_X1Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y176_OBUF (
.I(CLBLL_R_X73Y119_SLICE_X110Y119_AQ),
.O(RIOB33_X105Y175_IOB_X1Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y177_OBUF (
.I(CLBLM_L_X72Y119_SLICE_X109Y119_BQ),
.O(RIOB33_X105Y177_IOB_X1Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y178_OBUF (
.I(CLBLL_R_X73Y119_SLICE_X110Y119_BQ),
.O(RIOB33_X105Y177_IOB_X1Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y179_OBUF (
.I(CLBLM_L_X72Y119_SLICE_X108Y119_CQ),
.O(RIOB33_X105Y179_IOB_X1Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y180_OBUF (
.I(CLBLM_R_X67Y118_SLICE_X101Y118_AQ),
.O(RIOB33_X105Y179_IOB_X1Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y181_OBUF (
.I(CLBLL_R_X75Y133_SLICE_X114Y133_BQ),
.O(RIOB33_X105Y181_IOB_X1Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y182_OBUF (
.I(CLBLL_R_X77Y128_SLICE_X119Y128_BQ),
.O(RIOB33_X105Y181_IOB_X1Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y183_OBUF (
.I(1'b0),
.O(RIOB33_X105Y183_IOB_X1Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y184_OBUF (
.I(1'b0),
.O(RIOB33_X105Y183_IOB_X1Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y185_OBUF (
.I(CLBLL_R_X71Y117_SLICE_X106Y117_A5Q),
.O(RIOB33_X105Y185_IOB_X1Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y186_OBUF (
.I(1'b0),
.O(RIOB33_X105Y185_IOB_X1Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y187_OBUF (
.I(CLBLL_R_X73Y108_SLICE_X110Y108_AQ),
.O(RIOB33_X105Y187_IOB_X1Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y188_OBUF (
.I(CLBLL_R_X71Y117_SLICE_X106Y117_B5Q),
.O(RIOB33_X105Y187_IOB_X1Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y189_OBUF (
.I(1'b0),
.O(RIOB33_X105Y189_IOB_X1Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y190_OBUF (
.I(CLBLM_L_X76Y128_SLICE_X116Y128_C5Q),
.O(RIOB33_X105Y189_IOB_X1Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y191_OBUF (
.I(CLBLM_L_X68Y109_SLICE_X102Y109_AQ),
.O(RIOB33_X105Y191_IOB_X1Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y192_OBUF (
.I(CLBLM_L_X72Y118_SLICE_X109Y118_A5Q),
.O(RIOB33_X105Y191_IOB_X1Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y193_OBUF (
.I(1'b0),
.O(RIOB33_X105Y193_IOB_X1Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y194_OBUF (
.I(CLBLM_L_X76Y129_SLICE_X116Y129_CQ),
.O(RIOB33_X105Y193_IOB_X1Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y195_OBUF (
.I(CLBLL_R_X73Y104_SLICE_X110Y104_AQ),
.O(RIOB33_X105Y195_IOB_X1Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y196_OBUF (
.I(1'b0),
.O(RIOB33_X105Y195_IOB_X1Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y197_OBUF (
.I(CLBLL_R_X79Y135_SLICE_X122Y135_AQ),
.O(RIOB33_X105Y197_IOB_X1Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y198_OBUF (
.I(CLBLM_L_X80Y132_SLICE_X124Y132_AQ),
.O(RIOB33_X105Y197_IOB_X1Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y50_IOB_X1Y50_IBUF (
.I(RIOB33_SING_X105Y50_IOB_X1Y50_IPAD),
.O(RIOB33_SING_X105Y50_IOB_X1Y50_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y100_IOB_X1Y100_OBUF (
.I(CLBLM_L_X78Y104_SLICE_X120Y104_A5Q),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y149_IOB_X1Y149_OBUF (
.I(CLBLM_L_X76Y111_SLICE_X116Y111_BQ),
.O(RIOB33_SING_X105Y149_IOB_X1Y149_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y150_IOB_X1Y150_OBUF (
.I(1'b1),
.O(RIOB33_SING_X105Y150_IOB_X1Y150_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y199_IOB_X1Y199_OBUF (
.I(CLBLM_L_X74Y109_SLICE_X113Y109_AQ),
.O(RIOB33_SING_X105Y199_IOB_X1Y199_OPAD)
  );
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A = CLBLL_L_X2Y131_SLICE_X0Y131_AO6;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B = CLBLL_L_X2Y131_SLICE_X0Y131_BO6;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C = CLBLL_L_X2Y131_SLICE_X0Y131_CO6;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D = CLBLL_L_X2Y131_SLICE_X0Y131_DO6;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A = CLBLL_L_X2Y131_SLICE_X1Y131_AO6;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B = CLBLL_L_X2Y131_SLICE_X1Y131_BO6;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C = CLBLL_L_X2Y131_SLICE_X1Y131_CO6;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D = CLBLL_L_X2Y131_SLICE_X1Y131_DO6;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_A = CLBLL_L_X34Y123_SLICE_X50Y123_AO6;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_B = CLBLL_L_X34Y123_SLICE_X50Y123_BO6;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_C = CLBLL_L_X34Y123_SLICE_X50Y123_CO6;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_D = CLBLL_L_X34Y123_SLICE_X50Y123_DO6;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_A = CLBLL_L_X34Y123_SLICE_X51Y123_AO6;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_B = CLBLL_L_X34Y123_SLICE_X51Y123_BO6;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_C = CLBLL_L_X34Y123_SLICE_X51Y123_CO6;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_D = CLBLL_L_X34Y123_SLICE_X51Y123_DO6;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_A = CLBLL_L_X34Y126_SLICE_X50Y126_AO6;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_B = CLBLL_L_X34Y126_SLICE_X50Y126_BO6;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_C = CLBLL_L_X34Y126_SLICE_X50Y126_CO6;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_D = CLBLL_L_X34Y126_SLICE_X50Y126_DO6;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_A = CLBLL_L_X34Y126_SLICE_X51Y126_AO6;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_B = CLBLL_L_X34Y126_SLICE_X51Y126_BO6;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_C = CLBLL_L_X34Y126_SLICE_X51Y126_CO6;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_D = CLBLL_L_X34Y126_SLICE_X51Y126_DO6;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_A = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_B = CLBLL_L_X34Y128_SLICE_X50Y128_BO6;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_C = CLBLL_L_X34Y128_SLICE_X50Y128_CO6;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_D = CLBLL_L_X34Y128_SLICE_X50Y128_DO6;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_A = CLBLL_L_X34Y128_SLICE_X51Y128_AO6;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_B = CLBLL_L_X34Y128_SLICE_X51Y128_BO6;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_C = CLBLL_L_X34Y128_SLICE_X51Y128_CO6;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_D = CLBLL_L_X34Y128_SLICE_X51Y128_DO6;
  assign CLBLL_R_X71Y98_SLICE_X106Y98_A = CLBLL_R_X71Y98_SLICE_X106Y98_AO6;
  assign CLBLL_R_X71Y98_SLICE_X106Y98_B = CLBLL_R_X71Y98_SLICE_X106Y98_BO6;
  assign CLBLL_R_X71Y98_SLICE_X106Y98_C = CLBLL_R_X71Y98_SLICE_X106Y98_CO6;
  assign CLBLL_R_X71Y98_SLICE_X106Y98_D = CLBLL_R_X71Y98_SLICE_X106Y98_DO6;
  assign CLBLL_R_X71Y98_SLICE_X106Y98_AMUX = CLBLL_R_X71Y98_SLICE_X106Y98_A5Q;
  assign CLBLL_R_X71Y98_SLICE_X107Y98_A = CLBLL_R_X71Y98_SLICE_X107Y98_AO6;
  assign CLBLL_R_X71Y98_SLICE_X107Y98_B = CLBLL_R_X71Y98_SLICE_X107Y98_BO6;
  assign CLBLL_R_X71Y98_SLICE_X107Y98_C = CLBLL_R_X71Y98_SLICE_X107Y98_CO6;
  assign CLBLL_R_X71Y98_SLICE_X107Y98_D = CLBLL_R_X71Y98_SLICE_X107Y98_DO6;
  assign CLBLL_R_X71Y100_SLICE_X106Y100_A = CLBLL_R_X71Y100_SLICE_X106Y100_AO6;
  assign CLBLL_R_X71Y100_SLICE_X106Y100_B = CLBLL_R_X71Y100_SLICE_X106Y100_BO6;
  assign CLBLL_R_X71Y100_SLICE_X106Y100_C = CLBLL_R_X71Y100_SLICE_X106Y100_CO6;
  assign CLBLL_R_X71Y100_SLICE_X106Y100_D = CLBLL_R_X71Y100_SLICE_X106Y100_DO6;
  assign CLBLL_R_X71Y100_SLICE_X106Y100_AMUX = CLBLL_R_X71Y100_SLICE_X106Y100_AO5;
  assign CLBLL_R_X71Y100_SLICE_X107Y100_A = CLBLL_R_X71Y100_SLICE_X107Y100_AO6;
  assign CLBLL_R_X71Y100_SLICE_X107Y100_B = CLBLL_R_X71Y100_SLICE_X107Y100_BO6;
  assign CLBLL_R_X71Y100_SLICE_X107Y100_C = CLBLL_R_X71Y100_SLICE_X107Y100_CO6;
  assign CLBLL_R_X71Y100_SLICE_X107Y100_D = CLBLL_R_X71Y100_SLICE_X107Y100_DO6;
  assign CLBLL_R_X71Y101_SLICE_X106Y101_A = CLBLL_R_X71Y101_SLICE_X106Y101_AO6;
  assign CLBLL_R_X71Y101_SLICE_X106Y101_B = CLBLL_R_X71Y101_SLICE_X106Y101_BO6;
  assign CLBLL_R_X71Y101_SLICE_X106Y101_C = CLBLL_R_X71Y101_SLICE_X106Y101_CO6;
  assign CLBLL_R_X71Y101_SLICE_X106Y101_D = CLBLL_R_X71Y101_SLICE_X106Y101_DO6;
  assign CLBLL_R_X71Y101_SLICE_X107Y101_A = CLBLL_R_X71Y101_SLICE_X107Y101_AO6;
  assign CLBLL_R_X71Y101_SLICE_X107Y101_B = CLBLL_R_X71Y101_SLICE_X107Y101_BO6;
  assign CLBLL_R_X71Y101_SLICE_X107Y101_C = CLBLL_R_X71Y101_SLICE_X107Y101_CO6;
  assign CLBLL_R_X71Y101_SLICE_X107Y101_D = CLBLL_R_X71Y101_SLICE_X107Y101_DO6;
  assign CLBLL_R_X71Y102_SLICE_X106Y102_A = CLBLL_R_X71Y102_SLICE_X106Y102_AO6;
  assign CLBLL_R_X71Y102_SLICE_X106Y102_B = CLBLL_R_X71Y102_SLICE_X106Y102_BO6;
  assign CLBLL_R_X71Y102_SLICE_X106Y102_C = CLBLL_R_X71Y102_SLICE_X106Y102_CO6;
  assign CLBLL_R_X71Y102_SLICE_X106Y102_D = CLBLL_R_X71Y102_SLICE_X106Y102_DO6;
  assign CLBLL_R_X71Y102_SLICE_X107Y102_A = CLBLL_R_X71Y102_SLICE_X107Y102_AO6;
  assign CLBLL_R_X71Y102_SLICE_X107Y102_B = CLBLL_R_X71Y102_SLICE_X107Y102_BO6;
  assign CLBLL_R_X71Y102_SLICE_X107Y102_C = CLBLL_R_X71Y102_SLICE_X107Y102_CO6;
  assign CLBLL_R_X71Y102_SLICE_X107Y102_D = CLBLL_R_X71Y102_SLICE_X107Y102_DO6;
  assign CLBLL_R_X71Y103_SLICE_X106Y103_A = CLBLL_R_X71Y103_SLICE_X106Y103_AO6;
  assign CLBLL_R_X71Y103_SLICE_X106Y103_B = CLBLL_R_X71Y103_SLICE_X106Y103_BO6;
  assign CLBLL_R_X71Y103_SLICE_X106Y103_C = CLBLL_R_X71Y103_SLICE_X106Y103_CO6;
  assign CLBLL_R_X71Y103_SLICE_X106Y103_D = CLBLL_R_X71Y103_SLICE_X106Y103_DO6;
  assign CLBLL_R_X71Y103_SLICE_X106Y103_BMUX = CLBLL_R_X71Y103_SLICE_X106Y103_BO5;
  assign CLBLL_R_X71Y103_SLICE_X107Y103_A = CLBLL_R_X71Y103_SLICE_X107Y103_AO6;
  assign CLBLL_R_X71Y103_SLICE_X107Y103_B = CLBLL_R_X71Y103_SLICE_X107Y103_BO6;
  assign CLBLL_R_X71Y103_SLICE_X107Y103_C = CLBLL_R_X71Y103_SLICE_X107Y103_CO6;
  assign CLBLL_R_X71Y103_SLICE_X107Y103_D = CLBLL_R_X71Y103_SLICE_X107Y103_DO6;
  assign CLBLL_R_X71Y107_SLICE_X106Y107_A = CLBLL_R_X71Y107_SLICE_X106Y107_AO6;
  assign CLBLL_R_X71Y107_SLICE_X106Y107_B = CLBLL_R_X71Y107_SLICE_X106Y107_BO6;
  assign CLBLL_R_X71Y107_SLICE_X106Y107_C = CLBLL_R_X71Y107_SLICE_X106Y107_CO6;
  assign CLBLL_R_X71Y107_SLICE_X106Y107_D = CLBLL_R_X71Y107_SLICE_X106Y107_DO6;
  assign CLBLL_R_X71Y107_SLICE_X106Y107_BMUX = CLBLL_R_X71Y107_SLICE_X106Y107_BO5;
  assign CLBLL_R_X71Y107_SLICE_X106Y107_CMUX = CLBLL_R_X71Y107_SLICE_X106Y107_C5Q;
  assign CLBLL_R_X71Y107_SLICE_X107Y107_A = CLBLL_R_X71Y107_SLICE_X107Y107_AO6;
  assign CLBLL_R_X71Y107_SLICE_X107Y107_B = CLBLL_R_X71Y107_SLICE_X107Y107_BO6;
  assign CLBLL_R_X71Y107_SLICE_X107Y107_C = CLBLL_R_X71Y107_SLICE_X107Y107_CO6;
  assign CLBLL_R_X71Y107_SLICE_X107Y107_D = CLBLL_R_X71Y107_SLICE_X107Y107_DO6;
  assign CLBLL_R_X71Y107_SLICE_X107Y107_CMUX = CLBLL_R_X71Y107_SLICE_X107Y107_C5Q;
  assign CLBLL_R_X71Y108_SLICE_X106Y108_A = CLBLL_R_X71Y108_SLICE_X106Y108_AO6;
  assign CLBLL_R_X71Y108_SLICE_X106Y108_B = CLBLL_R_X71Y108_SLICE_X106Y108_BO6;
  assign CLBLL_R_X71Y108_SLICE_X106Y108_C = CLBLL_R_X71Y108_SLICE_X106Y108_CO6;
  assign CLBLL_R_X71Y108_SLICE_X106Y108_D = CLBLL_R_X71Y108_SLICE_X106Y108_DO6;
  assign CLBLL_R_X71Y108_SLICE_X106Y108_DMUX = CLBLL_R_X71Y108_SLICE_X106Y108_D5Q;
  assign CLBLL_R_X71Y108_SLICE_X107Y108_A = CLBLL_R_X71Y108_SLICE_X107Y108_AO6;
  assign CLBLL_R_X71Y108_SLICE_X107Y108_B = CLBLL_R_X71Y108_SLICE_X107Y108_BO6;
  assign CLBLL_R_X71Y108_SLICE_X107Y108_C = CLBLL_R_X71Y108_SLICE_X107Y108_CO6;
  assign CLBLL_R_X71Y108_SLICE_X107Y108_D = CLBLL_R_X71Y108_SLICE_X107Y108_DO6;
  assign CLBLL_R_X71Y108_SLICE_X107Y108_AMUX = CLBLL_R_X71Y108_SLICE_X107Y108_A5Q;
  assign CLBLL_R_X71Y109_SLICE_X106Y109_A = CLBLL_R_X71Y109_SLICE_X106Y109_AO6;
  assign CLBLL_R_X71Y109_SLICE_X106Y109_B = CLBLL_R_X71Y109_SLICE_X106Y109_BO6;
  assign CLBLL_R_X71Y109_SLICE_X106Y109_C = CLBLL_R_X71Y109_SLICE_X106Y109_CO6;
  assign CLBLL_R_X71Y109_SLICE_X106Y109_D = CLBLL_R_X71Y109_SLICE_X106Y109_DO6;
  assign CLBLL_R_X71Y109_SLICE_X106Y109_BMUX = CLBLL_R_X71Y109_SLICE_X106Y109_B5Q;
  assign CLBLL_R_X71Y109_SLICE_X106Y109_CMUX = CLBLL_R_X71Y109_SLICE_X106Y109_CO5;
  assign CLBLL_R_X71Y109_SLICE_X107Y109_A = CLBLL_R_X71Y109_SLICE_X107Y109_AO6;
  assign CLBLL_R_X71Y109_SLICE_X107Y109_B = CLBLL_R_X71Y109_SLICE_X107Y109_BO6;
  assign CLBLL_R_X71Y109_SLICE_X107Y109_C = CLBLL_R_X71Y109_SLICE_X107Y109_CO6;
  assign CLBLL_R_X71Y109_SLICE_X107Y109_D = CLBLL_R_X71Y109_SLICE_X107Y109_DO6;
  assign CLBLL_R_X71Y110_SLICE_X106Y110_A = CLBLL_R_X71Y110_SLICE_X106Y110_AO6;
  assign CLBLL_R_X71Y110_SLICE_X106Y110_B = CLBLL_R_X71Y110_SLICE_X106Y110_BO6;
  assign CLBLL_R_X71Y110_SLICE_X106Y110_C = CLBLL_R_X71Y110_SLICE_X106Y110_CO6;
  assign CLBLL_R_X71Y110_SLICE_X106Y110_D = CLBLL_R_X71Y110_SLICE_X106Y110_DO6;
  assign CLBLL_R_X71Y110_SLICE_X106Y110_AMUX = CLBLL_R_X71Y110_SLICE_X106Y110_A5Q;
  assign CLBLL_R_X71Y110_SLICE_X107Y110_A = CLBLL_R_X71Y110_SLICE_X107Y110_AO6;
  assign CLBLL_R_X71Y110_SLICE_X107Y110_B = CLBLL_R_X71Y110_SLICE_X107Y110_BO6;
  assign CLBLL_R_X71Y110_SLICE_X107Y110_C = CLBLL_R_X71Y110_SLICE_X107Y110_CO6;
  assign CLBLL_R_X71Y110_SLICE_X107Y110_D = CLBLL_R_X71Y110_SLICE_X107Y110_DO6;
  assign CLBLL_R_X71Y111_SLICE_X106Y111_A = CLBLL_R_X71Y111_SLICE_X106Y111_AO6;
  assign CLBLL_R_X71Y111_SLICE_X106Y111_B = CLBLL_R_X71Y111_SLICE_X106Y111_BO6;
  assign CLBLL_R_X71Y111_SLICE_X106Y111_C = CLBLL_R_X71Y111_SLICE_X106Y111_CO6;
  assign CLBLL_R_X71Y111_SLICE_X106Y111_D = CLBLL_R_X71Y111_SLICE_X106Y111_DO6;
  assign CLBLL_R_X71Y111_SLICE_X106Y111_AMUX = CLBLL_R_X71Y111_SLICE_X106Y111_A5Q;
  assign CLBLL_R_X71Y111_SLICE_X107Y111_A = CLBLL_R_X71Y111_SLICE_X107Y111_AO6;
  assign CLBLL_R_X71Y111_SLICE_X107Y111_B = CLBLL_R_X71Y111_SLICE_X107Y111_BO6;
  assign CLBLL_R_X71Y111_SLICE_X107Y111_C = CLBLL_R_X71Y111_SLICE_X107Y111_CO6;
  assign CLBLL_R_X71Y111_SLICE_X107Y111_D = CLBLL_R_X71Y111_SLICE_X107Y111_DO6;
  assign CLBLL_R_X71Y112_SLICE_X106Y112_A = CLBLL_R_X71Y112_SLICE_X106Y112_AO6;
  assign CLBLL_R_X71Y112_SLICE_X106Y112_B = CLBLL_R_X71Y112_SLICE_X106Y112_BO6;
  assign CLBLL_R_X71Y112_SLICE_X106Y112_C = CLBLL_R_X71Y112_SLICE_X106Y112_CO6;
  assign CLBLL_R_X71Y112_SLICE_X106Y112_D = CLBLL_R_X71Y112_SLICE_X106Y112_DO6;
  assign CLBLL_R_X71Y112_SLICE_X106Y112_BMUX = CLBLL_R_X71Y112_SLICE_X106Y112_B5Q;
  assign CLBLL_R_X71Y112_SLICE_X107Y112_A = CLBLL_R_X71Y112_SLICE_X107Y112_AO6;
  assign CLBLL_R_X71Y112_SLICE_X107Y112_B = CLBLL_R_X71Y112_SLICE_X107Y112_BO6;
  assign CLBLL_R_X71Y112_SLICE_X107Y112_C = CLBLL_R_X71Y112_SLICE_X107Y112_CO6;
  assign CLBLL_R_X71Y112_SLICE_X107Y112_D = CLBLL_R_X71Y112_SLICE_X107Y112_DO6;
  assign CLBLL_R_X71Y114_SLICE_X106Y114_A = CLBLL_R_X71Y114_SLICE_X106Y114_AO6;
  assign CLBLL_R_X71Y114_SLICE_X106Y114_B = CLBLL_R_X71Y114_SLICE_X106Y114_BO6;
  assign CLBLL_R_X71Y114_SLICE_X106Y114_C = CLBLL_R_X71Y114_SLICE_X106Y114_CO6;
  assign CLBLL_R_X71Y114_SLICE_X106Y114_D = CLBLL_R_X71Y114_SLICE_X106Y114_DO6;
  assign CLBLL_R_X71Y114_SLICE_X107Y114_A = CLBLL_R_X71Y114_SLICE_X107Y114_AO6;
  assign CLBLL_R_X71Y114_SLICE_X107Y114_B = CLBLL_R_X71Y114_SLICE_X107Y114_BO6;
  assign CLBLL_R_X71Y114_SLICE_X107Y114_C = CLBLL_R_X71Y114_SLICE_X107Y114_CO6;
  assign CLBLL_R_X71Y114_SLICE_X107Y114_D = CLBLL_R_X71Y114_SLICE_X107Y114_DO6;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_A = CLBLL_R_X71Y117_SLICE_X106Y117_AO6;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_B = CLBLL_R_X71Y117_SLICE_X106Y117_BO6;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_C = CLBLL_R_X71Y117_SLICE_X106Y117_CO6;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_D = CLBLL_R_X71Y117_SLICE_X106Y117_DO6;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_AMUX = CLBLL_R_X71Y117_SLICE_X106Y117_A5Q;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_BMUX = CLBLL_R_X71Y117_SLICE_X106Y117_B5Q;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_A = CLBLL_R_X71Y117_SLICE_X107Y117_AO6;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_B = CLBLL_R_X71Y117_SLICE_X107Y117_BO6;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_C = CLBLL_R_X71Y117_SLICE_X107Y117_CO6;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_D = CLBLL_R_X71Y117_SLICE_X107Y117_DO6;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_A = CLBLL_R_X71Y119_SLICE_X106Y119_AO6;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_B = CLBLL_R_X71Y119_SLICE_X106Y119_BO6;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_C = CLBLL_R_X71Y119_SLICE_X106Y119_CO6;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_D = CLBLL_R_X71Y119_SLICE_X106Y119_DO6;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_AMUX = CLBLL_R_X71Y119_SLICE_X106Y119_A5Q;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_A = CLBLL_R_X71Y119_SLICE_X107Y119_AO6;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_B = CLBLL_R_X71Y119_SLICE_X107Y119_BO6;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_C = CLBLL_R_X71Y119_SLICE_X107Y119_CO6;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_D = CLBLL_R_X71Y119_SLICE_X107Y119_DO6;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_A = CLBLL_R_X71Y121_SLICE_X106Y121_AO6;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_B = CLBLL_R_X71Y121_SLICE_X106Y121_BO6;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_C = CLBLL_R_X71Y121_SLICE_X106Y121_CO6;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_D = CLBLL_R_X71Y121_SLICE_X106Y121_DO6;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_AMUX = CLBLL_R_X71Y121_SLICE_X106Y121_A5Q;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_BMUX = CLBLL_R_X71Y121_SLICE_X106Y121_BO5;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_A = CLBLL_R_X71Y121_SLICE_X107Y121_AO6;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_B = CLBLL_R_X71Y121_SLICE_X107Y121_BO6;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_C = CLBLL_R_X71Y121_SLICE_X107Y121_CO6;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_D = CLBLL_R_X71Y121_SLICE_X107Y121_DO6;
  assign CLBLL_R_X71Y124_SLICE_X106Y124_A = CLBLL_R_X71Y124_SLICE_X106Y124_AO6;
  assign CLBLL_R_X71Y124_SLICE_X106Y124_B = CLBLL_R_X71Y124_SLICE_X106Y124_BO6;
  assign CLBLL_R_X71Y124_SLICE_X106Y124_C = CLBLL_R_X71Y124_SLICE_X106Y124_CO6;
  assign CLBLL_R_X71Y124_SLICE_X106Y124_D = CLBLL_R_X71Y124_SLICE_X106Y124_DO6;
  assign CLBLL_R_X71Y124_SLICE_X106Y124_AMUX = CLBLL_R_X71Y124_SLICE_X106Y124_A5Q;
  assign CLBLL_R_X71Y124_SLICE_X107Y124_A = CLBLL_R_X71Y124_SLICE_X107Y124_AO6;
  assign CLBLL_R_X71Y124_SLICE_X107Y124_B = CLBLL_R_X71Y124_SLICE_X107Y124_BO6;
  assign CLBLL_R_X71Y124_SLICE_X107Y124_C = CLBLL_R_X71Y124_SLICE_X107Y124_CO6;
  assign CLBLL_R_X71Y124_SLICE_X107Y124_D = CLBLL_R_X71Y124_SLICE_X107Y124_DO6;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_A = CLBLL_R_X71Y125_SLICE_X106Y125_AO6;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_B = CLBLL_R_X71Y125_SLICE_X106Y125_BO6;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_C = CLBLL_R_X71Y125_SLICE_X106Y125_CO6;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_D = CLBLL_R_X71Y125_SLICE_X106Y125_DO6;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_A = CLBLL_R_X71Y125_SLICE_X107Y125_AO6;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_B = CLBLL_R_X71Y125_SLICE_X107Y125_BO6;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_C = CLBLL_R_X71Y125_SLICE_X107Y125_CO6;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_D = CLBLL_R_X71Y125_SLICE_X107Y125_DO6;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_A = CLBLL_R_X71Y126_SLICE_X106Y126_AO6;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_B = CLBLL_R_X71Y126_SLICE_X106Y126_BO6;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_C = CLBLL_R_X71Y126_SLICE_X106Y126_CO6;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_D = CLBLL_R_X71Y126_SLICE_X106Y126_DO6;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_A = CLBLL_R_X71Y126_SLICE_X107Y126_AO6;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_B = CLBLL_R_X71Y126_SLICE_X107Y126_BO6;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_C = CLBLL_R_X71Y126_SLICE_X107Y126_CO6;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_D = CLBLL_R_X71Y126_SLICE_X107Y126_DO6;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_AMUX = CLBLL_R_X71Y126_SLICE_X107Y126_AO5;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_BMUX = CLBLL_R_X71Y126_SLICE_X107Y126_BO5;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_A = CLBLL_R_X71Y127_SLICE_X106Y127_AO6;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_B = CLBLL_R_X71Y127_SLICE_X106Y127_BO6;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_C = CLBLL_R_X71Y127_SLICE_X106Y127_CO6;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_D = CLBLL_R_X71Y127_SLICE_X106Y127_DO6;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_A = CLBLL_R_X71Y127_SLICE_X107Y127_AO6;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_B = CLBLL_R_X71Y127_SLICE_X107Y127_BO6;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_C = CLBLL_R_X71Y127_SLICE_X107Y127_CO6;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_D = CLBLL_R_X71Y127_SLICE_X107Y127_DO6;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_AMUX = CLBLL_R_X71Y127_SLICE_X107Y127_AO5;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_A = CLBLL_R_X71Y128_SLICE_X106Y128_AO6;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_B = CLBLL_R_X71Y128_SLICE_X106Y128_BO6;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_C = CLBLL_R_X71Y128_SLICE_X106Y128_CO6;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_D = CLBLL_R_X71Y128_SLICE_X106Y128_DO6;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_A = CLBLL_R_X71Y128_SLICE_X107Y128_AO6;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_B = CLBLL_R_X71Y128_SLICE_X107Y128_BO6;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_C = CLBLL_R_X71Y128_SLICE_X107Y128_CO6;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_D = CLBLL_R_X71Y128_SLICE_X107Y128_DO6;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_A = CLBLL_R_X71Y129_SLICE_X106Y129_AO6;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_B = CLBLL_R_X71Y129_SLICE_X106Y129_BO6;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_C = CLBLL_R_X71Y129_SLICE_X106Y129_CO6;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_D = CLBLL_R_X71Y129_SLICE_X106Y129_DO6;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_AMUX = CLBLL_R_X71Y129_SLICE_X106Y129_AO6;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_A = CLBLL_R_X71Y129_SLICE_X107Y129_AO6;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_B = CLBLL_R_X71Y129_SLICE_X107Y129_BO6;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_C = CLBLL_R_X71Y129_SLICE_X107Y129_CO6;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_D = CLBLL_R_X71Y129_SLICE_X107Y129_DO6;
  assign CLBLL_R_X71Y130_SLICE_X106Y130_A = CLBLL_R_X71Y130_SLICE_X106Y130_AO6;
  assign CLBLL_R_X71Y130_SLICE_X106Y130_B = CLBLL_R_X71Y130_SLICE_X106Y130_BO6;
  assign CLBLL_R_X71Y130_SLICE_X106Y130_C = CLBLL_R_X71Y130_SLICE_X106Y130_CO6;
  assign CLBLL_R_X71Y130_SLICE_X106Y130_D = CLBLL_R_X71Y130_SLICE_X106Y130_DO6;
  assign CLBLL_R_X71Y130_SLICE_X106Y130_DMUX = CLBLL_R_X71Y130_SLICE_X106Y130_DO5;
  assign CLBLL_R_X71Y130_SLICE_X107Y130_A = CLBLL_R_X71Y130_SLICE_X107Y130_AO6;
  assign CLBLL_R_X71Y130_SLICE_X107Y130_B = CLBLL_R_X71Y130_SLICE_X107Y130_BO6;
  assign CLBLL_R_X71Y130_SLICE_X107Y130_C = CLBLL_R_X71Y130_SLICE_X107Y130_CO6;
  assign CLBLL_R_X71Y130_SLICE_X107Y130_D = CLBLL_R_X71Y130_SLICE_X107Y130_DO6;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_A = CLBLL_R_X71Y131_SLICE_X106Y131_AO6;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_B = CLBLL_R_X71Y131_SLICE_X106Y131_BO6;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_C = CLBLL_R_X71Y131_SLICE_X106Y131_CO6;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_D = CLBLL_R_X71Y131_SLICE_X106Y131_DO6;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_A = CLBLL_R_X71Y131_SLICE_X107Y131_AO6;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_B = CLBLL_R_X71Y131_SLICE_X107Y131_BO6;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_C = CLBLL_R_X71Y131_SLICE_X107Y131_CO6;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_D = CLBLL_R_X71Y131_SLICE_X107Y131_DO6;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_AMUX = CLBLL_R_X71Y131_SLICE_X107Y131_A5Q;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_DMUX = CLBLL_R_X71Y131_SLICE_X107Y131_DO5;
  assign CLBLL_R_X71Y132_SLICE_X106Y132_A = CLBLL_R_X71Y132_SLICE_X106Y132_AO6;
  assign CLBLL_R_X71Y132_SLICE_X106Y132_B = CLBLL_R_X71Y132_SLICE_X106Y132_BO6;
  assign CLBLL_R_X71Y132_SLICE_X106Y132_C = CLBLL_R_X71Y132_SLICE_X106Y132_CO6;
  assign CLBLL_R_X71Y132_SLICE_X106Y132_D = CLBLL_R_X71Y132_SLICE_X106Y132_DO6;
  assign CLBLL_R_X71Y132_SLICE_X106Y132_AMUX = CLBLL_R_X71Y132_SLICE_X106Y132_AO5;
  assign CLBLL_R_X71Y132_SLICE_X107Y132_A = CLBLL_R_X71Y132_SLICE_X107Y132_AO6;
  assign CLBLL_R_X71Y132_SLICE_X107Y132_B = CLBLL_R_X71Y132_SLICE_X107Y132_BO6;
  assign CLBLL_R_X71Y132_SLICE_X107Y132_C = CLBLL_R_X71Y132_SLICE_X107Y132_CO6;
  assign CLBLL_R_X71Y132_SLICE_X107Y132_D = CLBLL_R_X71Y132_SLICE_X107Y132_DO6;
  assign CLBLL_R_X71Y133_SLICE_X106Y133_A = CLBLL_R_X71Y133_SLICE_X106Y133_AO6;
  assign CLBLL_R_X71Y133_SLICE_X106Y133_B = CLBLL_R_X71Y133_SLICE_X106Y133_BO6;
  assign CLBLL_R_X71Y133_SLICE_X106Y133_C = CLBLL_R_X71Y133_SLICE_X106Y133_CO6;
  assign CLBLL_R_X71Y133_SLICE_X106Y133_D = CLBLL_R_X71Y133_SLICE_X106Y133_DO6;
  assign CLBLL_R_X71Y133_SLICE_X107Y133_A = CLBLL_R_X71Y133_SLICE_X107Y133_AO6;
  assign CLBLL_R_X71Y133_SLICE_X107Y133_B = CLBLL_R_X71Y133_SLICE_X107Y133_BO6;
  assign CLBLL_R_X71Y133_SLICE_X107Y133_C = CLBLL_R_X71Y133_SLICE_X107Y133_CO6;
  assign CLBLL_R_X71Y133_SLICE_X107Y133_D = CLBLL_R_X71Y133_SLICE_X107Y133_DO6;
  assign CLBLL_R_X71Y133_SLICE_X107Y133_CMUX = CLBLL_R_X71Y133_SLICE_X107Y133_CO6;
  assign CLBLL_R_X71Y134_SLICE_X106Y134_A = CLBLL_R_X71Y134_SLICE_X106Y134_AO6;
  assign CLBLL_R_X71Y134_SLICE_X106Y134_B = CLBLL_R_X71Y134_SLICE_X106Y134_BO6;
  assign CLBLL_R_X71Y134_SLICE_X106Y134_C = CLBLL_R_X71Y134_SLICE_X106Y134_CO6;
  assign CLBLL_R_X71Y134_SLICE_X106Y134_D = CLBLL_R_X71Y134_SLICE_X106Y134_DO6;
  assign CLBLL_R_X71Y134_SLICE_X107Y134_A = CLBLL_R_X71Y134_SLICE_X107Y134_AO6;
  assign CLBLL_R_X71Y134_SLICE_X107Y134_B = CLBLL_R_X71Y134_SLICE_X107Y134_BO6;
  assign CLBLL_R_X71Y134_SLICE_X107Y134_C = CLBLL_R_X71Y134_SLICE_X107Y134_CO6;
  assign CLBLL_R_X71Y134_SLICE_X107Y134_D = CLBLL_R_X71Y134_SLICE_X107Y134_DO6;
  assign CLBLL_R_X73Y101_SLICE_X110Y101_A = CLBLL_R_X73Y101_SLICE_X110Y101_AO6;
  assign CLBLL_R_X73Y101_SLICE_X110Y101_B = CLBLL_R_X73Y101_SLICE_X110Y101_BO6;
  assign CLBLL_R_X73Y101_SLICE_X110Y101_C = CLBLL_R_X73Y101_SLICE_X110Y101_CO6;
  assign CLBLL_R_X73Y101_SLICE_X110Y101_D = CLBLL_R_X73Y101_SLICE_X110Y101_DO6;
  assign CLBLL_R_X73Y101_SLICE_X111Y101_A = CLBLL_R_X73Y101_SLICE_X111Y101_AO6;
  assign CLBLL_R_X73Y101_SLICE_X111Y101_B = CLBLL_R_X73Y101_SLICE_X111Y101_BO6;
  assign CLBLL_R_X73Y101_SLICE_X111Y101_C = CLBLL_R_X73Y101_SLICE_X111Y101_CO6;
  assign CLBLL_R_X73Y101_SLICE_X111Y101_D = CLBLL_R_X73Y101_SLICE_X111Y101_DO6;
  assign CLBLL_R_X73Y102_SLICE_X110Y102_A = CLBLL_R_X73Y102_SLICE_X110Y102_AO6;
  assign CLBLL_R_X73Y102_SLICE_X110Y102_B = CLBLL_R_X73Y102_SLICE_X110Y102_BO6;
  assign CLBLL_R_X73Y102_SLICE_X110Y102_C = CLBLL_R_X73Y102_SLICE_X110Y102_CO6;
  assign CLBLL_R_X73Y102_SLICE_X110Y102_D = CLBLL_R_X73Y102_SLICE_X110Y102_DO6;
  assign CLBLL_R_X73Y102_SLICE_X110Y102_AMUX = CLBLL_R_X73Y102_SLICE_X110Y102_A5Q;
  assign CLBLL_R_X73Y102_SLICE_X111Y102_A = CLBLL_R_X73Y102_SLICE_X111Y102_AO6;
  assign CLBLL_R_X73Y102_SLICE_X111Y102_B = CLBLL_R_X73Y102_SLICE_X111Y102_BO6;
  assign CLBLL_R_X73Y102_SLICE_X111Y102_C = CLBLL_R_X73Y102_SLICE_X111Y102_CO6;
  assign CLBLL_R_X73Y102_SLICE_X111Y102_D = CLBLL_R_X73Y102_SLICE_X111Y102_DO6;
  assign CLBLL_R_X73Y102_SLICE_X111Y102_AMUX = CLBLL_R_X73Y102_SLICE_X111Y102_A5Q;
  assign CLBLL_R_X73Y103_SLICE_X110Y103_A = CLBLL_R_X73Y103_SLICE_X110Y103_AO6;
  assign CLBLL_R_X73Y103_SLICE_X110Y103_B = CLBLL_R_X73Y103_SLICE_X110Y103_BO6;
  assign CLBLL_R_X73Y103_SLICE_X110Y103_C = CLBLL_R_X73Y103_SLICE_X110Y103_CO6;
  assign CLBLL_R_X73Y103_SLICE_X110Y103_D = CLBLL_R_X73Y103_SLICE_X110Y103_DO6;
  assign CLBLL_R_X73Y103_SLICE_X110Y103_AMUX = CLBLL_R_X73Y103_SLICE_X110Y103_A5Q;
  assign CLBLL_R_X73Y103_SLICE_X110Y103_BMUX = CLBLL_R_X73Y103_SLICE_X110Y103_B5Q;
  assign CLBLL_R_X73Y103_SLICE_X110Y103_CMUX = CLBLL_R_X73Y103_SLICE_X110Y103_CO5;
  assign CLBLL_R_X73Y103_SLICE_X110Y103_DMUX = CLBLL_R_X73Y103_SLICE_X110Y103_DO6;
  assign CLBLL_R_X73Y103_SLICE_X111Y103_A = CLBLL_R_X73Y103_SLICE_X111Y103_AO6;
  assign CLBLL_R_X73Y103_SLICE_X111Y103_B = CLBLL_R_X73Y103_SLICE_X111Y103_BO6;
  assign CLBLL_R_X73Y103_SLICE_X111Y103_C = CLBLL_R_X73Y103_SLICE_X111Y103_CO6;
  assign CLBLL_R_X73Y103_SLICE_X111Y103_D = CLBLL_R_X73Y103_SLICE_X111Y103_DO6;
  assign CLBLL_R_X73Y103_SLICE_X111Y103_AMUX = CLBLL_R_X73Y103_SLICE_X111Y103_A5Q;
  assign CLBLL_R_X73Y104_SLICE_X110Y104_A = CLBLL_R_X73Y104_SLICE_X110Y104_AO6;
  assign CLBLL_R_X73Y104_SLICE_X110Y104_B = CLBLL_R_X73Y104_SLICE_X110Y104_BO6;
  assign CLBLL_R_X73Y104_SLICE_X110Y104_C = CLBLL_R_X73Y104_SLICE_X110Y104_CO6;
  assign CLBLL_R_X73Y104_SLICE_X110Y104_D = CLBLL_R_X73Y104_SLICE_X110Y104_DO6;
  assign CLBLL_R_X73Y104_SLICE_X110Y104_AMUX = CLBLL_R_X73Y104_SLICE_X110Y104_A5Q;
  assign CLBLL_R_X73Y104_SLICE_X110Y104_BMUX = CLBLL_R_X73Y104_SLICE_X110Y104_BO5;
  assign CLBLL_R_X73Y104_SLICE_X110Y104_DMUX = CLBLL_R_X73Y104_SLICE_X110Y104_DO5;
  assign CLBLL_R_X73Y104_SLICE_X111Y104_A = CLBLL_R_X73Y104_SLICE_X111Y104_AO6;
  assign CLBLL_R_X73Y104_SLICE_X111Y104_B = CLBLL_R_X73Y104_SLICE_X111Y104_BO6;
  assign CLBLL_R_X73Y104_SLICE_X111Y104_C = CLBLL_R_X73Y104_SLICE_X111Y104_CO6;
  assign CLBLL_R_X73Y104_SLICE_X111Y104_D = CLBLL_R_X73Y104_SLICE_X111Y104_DO6;
  assign CLBLL_R_X73Y104_SLICE_X111Y104_DMUX = CLBLL_R_X73Y104_SLICE_X111Y104_DO6;
  assign CLBLL_R_X73Y106_SLICE_X110Y106_A = CLBLL_R_X73Y106_SLICE_X110Y106_AO6;
  assign CLBLL_R_X73Y106_SLICE_X110Y106_B = CLBLL_R_X73Y106_SLICE_X110Y106_BO6;
  assign CLBLL_R_X73Y106_SLICE_X110Y106_C = CLBLL_R_X73Y106_SLICE_X110Y106_CO6;
  assign CLBLL_R_X73Y106_SLICE_X110Y106_D = CLBLL_R_X73Y106_SLICE_X110Y106_DO6;
  assign CLBLL_R_X73Y106_SLICE_X111Y106_A = CLBLL_R_X73Y106_SLICE_X111Y106_AO6;
  assign CLBLL_R_X73Y106_SLICE_X111Y106_B = CLBLL_R_X73Y106_SLICE_X111Y106_BO6;
  assign CLBLL_R_X73Y106_SLICE_X111Y106_C = CLBLL_R_X73Y106_SLICE_X111Y106_CO6;
  assign CLBLL_R_X73Y106_SLICE_X111Y106_D = CLBLL_R_X73Y106_SLICE_X111Y106_DO6;
  assign CLBLL_R_X73Y107_SLICE_X110Y107_A = CLBLL_R_X73Y107_SLICE_X110Y107_AO6;
  assign CLBLL_R_X73Y107_SLICE_X110Y107_B = CLBLL_R_X73Y107_SLICE_X110Y107_BO6;
  assign CLBLL_R_X73Y107_SLICE_X110Y107_C = CLBLL_R_X73Y107_SLICE_X110Y107_CO6;
  assign CLBLL_R_X73Y107_SLICE_X110Y107_D = CLBLL_R_X73Y107_SLICE_X110Y107_DO6;
  assign CLBLL_R_X73Y107_SLICE_X111Y107_A = CLBLL_R_X73Y107_SLICE_X111Y107_AO6;
  assign CLBLL_R_X73Y107_SLICE_X111Y107_B = CLBLL_R_X73Y107_SLICE_X111Y107_BO6;
  assign CLBLL_R_X73Y107_SLICE_X111Y107_C = CLBLL_R_X73Y107_SLICE_X111Y107_CO6;
  assign CLBLL_R_X73Y107_SLICE_X111Y107_D = CLBLL_R_X73Y107_SLICE_X111Y107_DO6;
  assign CLBLL_R_X73Y108_SLICE_X110Y108_A = CLBLL_R_X73Y108_SLICE_X110Y108_AO6;
  assign CLBLL_R_X73Y108_SLICE_X110Y108_B = CLBLL_R_X73Y108_SLICE_X110Y108_BO6;
  assign CLBLL_R_X73Y108_SLICE_X110Y108_C = CLBLL_R_X73Y108_SLICE_X110Y108_CO6;
  assign CLBLL_R_X73Y108_SLICE_X110Y108_D = CLBLL_R_X73Y108_SLICE_X110Y108_DO6;
  assign CLBLL_R_X73Y108_SLICE_X110Y108_AMUX = CLBLL_R_X73Y108_SLICE_X110Y108_A5Q;
  assign CLBLL_R_X73Y108_SLICE_X111Y108_A = CLBLL_R_X73Y108_SLICE_X111Y108_AO6;
  assign CLBLL_R_X73Y108_SLICE_X111Y108_B = CLBLL_R_X73Y108_SLICE_X111Y108_BO6;
  assign CLBLL_R_X73Y108_SLICE_X111Y108_C = CLBLL_R_X73Y108_SLICE_X111Y108_CO6;
  assign CLBLL_R_X73Y108_SLICE_X111Y108_D = CLBLL_R_X73Y108_SLICE_X111Y108_DO6;
  assign CLBLL_R_X73Y109_SLICE_X110Y109_A = CLBLL_R_X73Y109_SLICE_X110Y109_AO6;
  assign CLBLL_R_X73Y109_SLICE_X110Y109_B = CLBLL_R_X73Y109_SLICE_X110Y109_BO6;
  assign CLBLL_R_X73Y109_SLICE_X110Y109_C = CLBLL_R_X73Y109_SLICE_X110Y109_CO6;
  assign CLBLL_R_X73Y109_SLICE_X110Y109_D = CLBLL_R_X73Y109_SLICE_X110Y109_DO6;
  assign CLBLL_R_X73Y109_SLICE_X111Y109_A = CLBLL_R_X73Y109_SLICE_X111Y109_AO6;
  assign CLBLL_R_X73Y109_SLICE_X111Y109_B = CLBLL_R_X73Y109_SLICE_X111Y109_BO6;
  assign CLBLL_R_X73Y109_SLICE_X111Y109_C = CLBLL_R_X73Y109_SLICE_X111Y109_CO6;
  assign CLBLL_R_X73Y109_SLICE_X111Y109_D = CLBLL_R_X73Y109_SLICE_X111Y109_DO6;
  assign CLBLL_R_X73Y111_SLICE_X110Y111_A = CLBLL_R_X73Y111_SLICE_X110Y111_AO6;
  assign CLBLL_R_X73Y111_SLICE_X110Y111_B = CLBLL_R_X73Y111_SLICE_X110Y111_BO6;
  assign CLBLL_R_X73Y111_SLICE_X110Y111_C = CLBLL_R_X73Y111_SLICE_X110Y111_CO6;
  assign CLBLL_R_X73Y111_SLICE_X110Y111_D = CLBLL_R_X73Y111_SLICE_X110Y111_DO6;
  assign CLBLL_R_X73Y111_SLICE_X110Y111_AMUX = CLBLL_R_X73Y111_SLICE_X110Y111_A5Q;
  assign CLBLL_R_X73Y111_SLICE_X111Y111_A = CLBLL_R_X73Y111_SLICE_X111Y111_AO6;
  assign CLBLL_R_X73Y111_SLICE_X111Y111_B = CLBLL_R_X73Y111_SLICE_X111Y111_BO6;
  assign CLBLL_R_X73Y111_SLICE_X111Y111_C = CLBLL_R_X73Y111_SLICE_X111Y111_CO6;
  assign CLBLL_R_X73Y111_SLICE_X111Y111_D = CLBLL_R_X73Y111_SLICE_X111Y111_DO6;
  assign CLBLL_R_X73Y113_SLICE_X110Y113_A = CLBLL_R_X73Y113_SLICE_X110Y113_AO6;
  assign CLBLL_R_X73Y113_SLICE_X110Y113_B = CLBLL_R_X73Y113_SLICE_X110Y113_BO6;
  assign CLBLL_R_X73Y113_SLICE_X110Y113_C = CLBLL_R_X73Y113_SLICE_X110Y113_CO6;
  assign CLBLL_R_X73Y113_SLICE_X110Y113_D = CLBLL_R_X73Y113_SLICE_X110Y113_DO6;
  assign CLBLL_R_X73Y113_SLICE_X110Y113_AMUX = CLBLL_R_X73Y113_SLICE_X110Y113_A5Q;
  assign CLBLL_R_X73Y113_SLICE_X111Y113_A = CLBLL_R_X73Y113_SLICE_X111Y113_AO6;
  assign CLBLL_R_X73Y113_SLICE_X111Y113_B = CLBLL_R_X73Y113_SLICE_X111Y113_BO6;
  assign CLBLL_R_X73Y113_SLICE_X111Y113_C = CLBLL_R_X73Y113_SLICE_X111Y113_CO6;
  assign CLBLL_R_X73Y113_SLICE_X111Y113_D = CLBLL_R_X73Y113_SLICE_X111Y113_DO6;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_A = CLBLL_R_X73Y118_SLICE_X110Y118_AO6;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_B = CLBLL_R_X73Y118_SLICE_X110Y118_BO6;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_C = CLBLL_R_X73Y118_SLICE_X110Y118_CO6;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_D = CLBLL_R_X73Y118_SLICE_X110Y118_DO6;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_BMUX = CLBLL_R_X73Y118_SLICE_X110Y118_B5Q;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_A = CLBLL_R_X73Y118_SLICE_X111Y118_AO6;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_B = CLBLL_R_X73Y118_SLICE_X111Y118_BO6;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_C = CLBLL_R_X73Y118_SLICE_X111Y118_CO6;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_D = CLBLL_R_X73Y118_SLICE_X111Y118_DO6;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_AMUX = CLBLL_R_X73Y118_SLICE_X111Y118_A5Q;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_A = CLBLL_R_X73Y119_SLICE_X110Y119_AO6;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_B = CLBLL_R_X73Y119_SLICE_X110Y119_BO6;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_C = CLBLL_R_X73Y119_SLICE_X110Y119_CO6;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_D = CLBLL_R_X73Y119_SLICE_X110Y119_DO6;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_AMUX = CLBLL_R_X73Y119_SLICE_X110Y119_A5Q;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_BMUX = CLBLL_R_X73Y119_SLICE_X110Y119_B5Q;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_CMUX = CLBLL_R_X73Y119_SLICE_X110Y119_CO6;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_A = CLBLL_R_X73Y119_SLICE_X111Y119_AO6;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_B = CLBLL_R_X73Y119_SLICE_X111Y119_BO6;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_C = CLBLL_R_X73Y119_SLICE_X111Y119_CO6;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_D = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_A = CLBLL_R_X73Y121_SLICE_X110Y121_AO6;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_B = CLBLL_R_X73Y121_SLICE_X110Y121_BO6;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_C = CLBLL_R_X73Y121_SLICE_X110Y121_CO6;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_D = CLBLL_R_X73Y121_SLICE_X110Y121_DO6;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_A = CLBLL_R_X73Y121_SLICE_X111Y121_AO6;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_B = CLBLL_R_X73Y121_SLICE_X111Y121_BO6;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_C = CLBLL_R_X73Y121_SLICE_X111Y121_CO6;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_D = CLBLL_R_X73Y121_SLICE_X111Y121_DO6;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_A = CLBLL_R_X73Y122_SLICE_X110Y122_AO6;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_B = CLBLL_R_X73Y122_SLICE_X110Y122_BO6;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_C = CLBLL_R_X73Y122_SLICE_X110Y122_CO6;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_D = CLBLL_R_X73Y122_SLICE_X110Y122_DO6;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_AMUX = CLBLL_R_X73Y122_SLICE_X110Y122_AO5;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_DMUX = CLBLL_R_X73Y122_SLICE_X110Y122_DO5;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_A = CLBLL_R_X73Y122_SLICE_X111Y122_AO6;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_B = CLBLL_R_X73Y122_SLICE_X111Y122_BO6;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_C = CLBLL_R_X73Y122_SLICE_X111Y122_CO6;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_D = CLBLL_R_X73Y122_SLICE_X111Y122_DO6;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_A = CLBLL_R_X73Y123_SLICE_X110Y123_AO6;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_B = CLBLL_R_X73Y123_SLICE_X110Y123_BO6;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_C = CLBLL_R_X73Y123_SLICE_X110Y123_CO6;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_D = CLBLL_R_X73Y123_SLICE_X110Y123_DO6;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_A = CLBLL_R_X73Y123_SLICE_X111Y123_AO6;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_B = CLBLL_R_X73Y123_SLICE_X111Y123_BO6;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_C = CLBLL_R_X73Y123_SLICE_X111Y123_CO6;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_D = CLBLL_R_X73Y123_SLICE_X111Y123_DO6;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_AMUX = CLBLL_R_X73Y123_SLICE_X111Y123_AO5;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_A = CLBLL_R_X73Y124_SLICE_X110Y124_AO6;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_B = CLBLL_R_X73Y124_SLICE_X110Y124_BO6;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_C = CLBLL_R_X73Y124_SLICE_X110Y124_CO6;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_D = CLBLL_R_X73Y124_SLICE_X110Y124_DO6;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_AMUX = CLBLL_R_X73Y124_SLICE_X110Y124_A5Q;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_CMUX = CLBLL_R_X73Y124_SLICE_X110Y124_CO5;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_A = CLBLL_R_X73Y124_SLICE_X111Y124_AO6;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_B = CLBLL_R_X73Y124_SLICE_X111Y124_BO6;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_C = CLBLL_R_X73Y124_SLICE_X111Y124_CO6;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_D = CLBLL_R_X73Y124_SLICE_X111Y124_DO6;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_A = CLBLL_R_X73Y125_SLICE_X110Y125_AO6;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_B = CLBLL_R_X73Y125_SLICE_X110Y125_BO6;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_C = CLBLL_R_X73Y125_SLICE_X110Y125_CO6;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_D = CLBLL_R_X73Y125_SLICE_X110Y125_DO6;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_BMUX = CLBLL_R_X73Y125_SLICE_X110Y125_BO6;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_A = CLBLL_R_X73Y125_SLICE_X111Y125_AO6;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_B = CLBLL_R_X73Y125_SLICE_X111Y125_BO6;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_C = CLBLL_R_X73Y125_SLICE_X111Y125_CO6;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_D = CLBLL_R_X73Y125_SLICE_X111Y125_DO6;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_AMUX = CLBLL_R_X73Y125_SLICE_X111Y125_A5Q;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_A = CLBLL_R_X73Y126_SLICE_X110Y126_AO6;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_B = CLBLL_R_X73Y126_SLICE_X110Y126_BO6;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_C = CLBLL_R_X73Y126_SLICE_X110Y126_CO6;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_D = CLBLL_R_X73Y126_SLICE_X110Y126_DO6;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_AMUX = CLBLL_R_X73Y126_SLICE_X110Y126_A5Q;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_CMUX = CLBLL_R_X73Y126_SLICE_X110Y126_CO5;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_A = CLBLL_R_X73Y126_SLICE_X111Y126_AO6;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_B = CLBLL_R_X73Y126_SLICE_X111Y126_BO6;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_C = CLBLL_R_X73Y126_SLICE_X111Y126_CO6;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_D = CLBLL_R_X73Y126_SLICE_X111Y126_DO6;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_BMUX = CLBLL_R_X73Y126_SLICE_X111Y126_BO5;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_A = CLBLL_R_X73Y127_SLICE_X110Y127_AO6;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_B = CLBLL_R_X73Y127_SLICE_X110Y127_BO6;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_C = CLBLL_R_X73Y127_SLICE_X110Y127_CO6;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_D = CLBLL_R_X73Y127_SLICE_X110Y127_DO6;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_AMUX = CLBLL_R_X73Y127_SLICE_X110Y127_A5Q;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_CMUX = CLBLL_R_X73Y127_SLICE_X110Y127_CO5;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_A = CLBLL_R_X73Y127_SLICE_X111Y127_AO6;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_B = CLBLL_R_X73Y127_SLICE_X111Y127_BO6;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_C = CLBLL_R_X73Y127_SLICE_X111Y127_CO6;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_D = CLBLL_R_X73Y127_SLICE_X111Y127_DO6;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_BMUX = CLBLL_R_X73Y127_SLICE_X111Y127_BO5;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_A = CLBLL_R_X73Y128_SLICE_X110Y128_AO6;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_B = CLBLL_R_X73Y128_SLICE_X110Y128_BO6;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_C = CLBLL_R_X73Y128_SLICE_X110Y128_CO6;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_D = CLBLL_R_X73Y128_SLICE_X110Y128_DO6;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_A = CLBLL_R_X73Y128_SLICE_X111Y128_AO6;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_B = CLBLL_R_X73Y128_SLICE_X111Y128_BO6;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_C = CLBLL_R_X73Y128_SLICE_X111Y128_CO6;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_D = CLBLL_R_X73Y128_SLICE_X111Y128_DO6;
  assign CLBLL_R_X73Y131_SLICE_X110Y131_A = CLBLL_R_X73Y131_SLICE_X110Y131_AO6;
  assign CLBLL_R_X73Y131_SLICE_X110Y131_B = CLBLL_R_X73Y131_SLICE_X110Y131_BO6;
  assign CLBLL_R_X73Y131_SLICE_X110Y131_C = CLBLL_R_X73Y131_SLICE_X110Y131_CO6;
  assign CLBLL_R_X73Y131_SLICE_X110Y131_D = CLBLL_R_X73Y131_SLICE_X110Y131_DO6;
  assign CLBLL_R_X73Y131_SLICE_X111Y131_A = CLBLL_R_X73Y131_SLICE_X111Y131_AO6;
  assign CLBLL_R_X73Y131_SLICE_X111Y131_B = CLBLL_R_X73Y131_SLICE_X111Y131_BO6;
  assign CLBLL_R_X73Y131_SLICE_X111Y131_C = CLBLL_R_X73Y131_SLICE_X111Y131_CO6;
  assign CLBLL_R_X73Y131_SLICE_X111Y131_D = CLBLL_R_X73Y131_SLICE_X111Y131_DO6;
  assign CLBLL_R_X73Y132_SLICE_X110Y132_A = CLBLL_R_X73Y132_SLICE_X110Y132_AO6;
  assign CLBLL_R_X73Y132_SLICE_X110Y132_B = CLBLL_R_X73Y132_SLICE_X110Y132_BO6;
  assign CLBLL_R_X73Y132_SLICE_X110Y132_C = CLBLL_R_X73Y132_SLICE_X110Y132_CO6;
  assign CLBLL_R_X73Y132_SLICE_X110Y132_D = CLBLL_R_X73Y132_SLICE_X110Y132_DO6;
  assign CLBLL_R_X73Y132_SLICE_X110Y132_AMUX = CLBLL_R_X73Y132_SLICE_X110Y132_AO5;
  assign CLBLL_R_X73Y132_SLICE_X111Y132_A = CLBLL_R_X73Y132_SLICE_X111Y132_AO6;
  assign CLBLL_R_X73Y132_SLICE_X111Y132_B = CLBLL_R_X73Y132_SLICE_X111Y132_BO6;
  assign CLBLL_R_X73Y132_SLICE_X111Y132_C = CLBLL_R_X73Y132_SLICE_X111Y132_CO6;
  assign CLBLL_R_X73Y132_SLICE_X111Y132_D = CLBLL_R_X73Y132_SLICE_X111Y132_DO6;
  assign CLBLL_R_X73Y132_SLICE_X111Y132_AMUX = CLBLL_R_X73Y132_SLICE_X111Y132_AO5;
  assign CLBLL_R_X73Y132_SLICE_X111Y132_CMUX = CLBLL_R_X73Y132_SLICE_X111Y132_CO6;
  assign CLBLL_R_X73Y133_SLICE_X110Y133_A = CLBLL_R_X73Y133_SLICE_X110Y133_AO6;
  assign CLBLL_R_X73Y133_SLICE_X110Y133_B = CLBLL_R_X73Y133_SLICE_X110Y133_BO6;
  assign CLBLL_R_X73Y133_SLICE_X110Y133_C = CLBLL_R_X73Y133_SLICE_X110Y133_CO6;
  assign CLBLL_R_X73Y133_SLICE_X110Y133_D = CLBLL_R_X73Y133_SLICE_X110Y133_DO6;
  assign CLBLL_R_X73Y133_SLICE_X110Y133_AMUX = CLBLL_R_X73Y133_SLICE_X110Y133_A5Q;
  assign CLBLL_R_X73Y133_SLICE_X111Y133_A = CLBLL_R_X73Y133_SLICE_X111Y133_AO6;
  assign CLBLL_R_X73Y133_SLICE_X111Y133_B = CLBLL_R_X73Y133_SLICE_X111Y133_BO6;
  assign CLBLL_R_X73Y133_SLICE_X111Y133_C = CLBLL_R_X73Y133_SLICE_X111Y133_CO6;
  assign CLBLL_R_X73Y133_SLICE_X111Y133_D = CLBLL_R_X73Y133_SLICE_X111Y133_DO6;
  assign CLBLL_R_X73Y133_SLICE_X111Y133_AMUX = CLBLL_R_X73Y133_SLICE_X111Y133_A5Q;
  assign CLBLL_R_X73Y133_SLICE_X111Y133_BMUX = CLBLL_R_X73Y133_SLICE_X111Y133_BO6;
  assign CLBLL_R_X73Y134_SLICE_X110Y134_A = CLBLL_R_X73Y134_SLICE_X110Y134_AO6;
  assign CLBLL_R_X73Y134_SLICE_X110Y134_B = CLBLL_R_X73Y134_SLICE_X110Y134_BO6;
  assign CLBLL_R_X73Y134_SLICE_X110Y134_C = CLBLL_R_X73Y134_SLICE_X110Y134_CO6;
  assign CLBLL_R_X73Y134_SLICE_X110Y134_D = CLBLL_R_X73Y134_SLICE_X110Y134_DO6;
  assign CLBLL_R_X73Y134_SLICE_X110Y134_AMUX = CLBLL_R_X73Y134_SLICE_X110Y134_AO5;
  assign CLBLL_R_X73Y134_SLICE_X111Y134_A = CLBLL_R_X73Y134_SLICE_X111Y134_AO6;
  assign CLBLL_R_X73Y134_SLICE_X111Y134_B = CLBLL_R_X73Y134_SLICE_X111Y134_BO6;
  assign CLBLL_R_X73Y134_SLICE_X111Y134_C = CLBLL_R_X73Y134_SLICE_X111Y134_CO6;
  assign CLBLL_R_X73Y134_SLICE_X111Y134_D = CLBLL_R_X73Y134_SLICE_X111Y134_DO6;
  assign CLBLL_R_X75Y103_SLICE_X114Y103_A = CLBLL_R_X75Y103_SLICE_X114Y103_AO6;
  assign CLBLL_R_X75Y103_SLICE_X114Y103_B = CLBLL_R_X75Y103_SLICE_X114Y103_BO6;
  assign CLBLL_R_X75Y103_SLICE_X114Y103_C = CLBLL_R_X75Y103_SLICE_X114Y103_CO6;
  assign CLBLL_R_X75Y103_SLICE_X114Y103_D = CLBLL_R_X75Y103_SLICE_X114Y103_DO6;
  assign CLBLL_R_X75Y103_SLICE_X115Y103_A = CLBLL_R_X75Y103_SLICE_X115Y103_AO6;
  assign CLBLL_R_X75Y103_SLICE_X115Y103_B = CLBLL_R_X75Y103_SLICE_X115Y103_BO6;
  assign CLBLL_R_X75Y103_SLICE_X115Y103_C = CLBLL_R_X75Y103_SLICE_X115Y103_CO6;
  assign CLBLL_R_X75Y103_SLICE_X115Y103_D = CLBLL_R_X75Y103_SLICE_X115Y103_DO6;
  assign CLBLL_R_X75Y107_SLICE_X114Y107_A = CLBLL_R_X75Y107_SLICE_X114Y107_AO6;
  assign CLBLL_R_X75Y107_SLICE_X114Y107_B = CLBLL_R_X75Y107_SLICE_X114Y107_BO6;
  assign CLBLL_R_X75Y107_SLICE_X114Y107_C = CLBLL_R_X75Y107_SLICE_X114Y107_CO6;
  assign CLBLL_R_X75Y107_SLICE_X114Y107_D = CLBLL_R_X75Y107_SLICE_X114Y107_DO6;
  assign CLBLL_R_X75Y107_SLICE_X115Y107_A = CLBLL_R_X75Y107_SLICE_X115Y107_AO6;
  assign CLBLL_R_X75Y107_SLICE_X115Y107_B = CLBLL_R_X75Y107_SLICE_X115Y107_BO6;
  assign CLBLL_R_X75Y107_SLICE_X115Y107_C = CLBLL_R_X75Y107_SLICE_X115Y107_CO6;
  assign CLBLL_R_X75Y107_SLICE_X115Y107_D = CLBLL_R_X75Y107_SLICE_X115Y107_DO6;
  assign CLBLL_R_X75Y113_SLICE_X114Y113_A = CLBLL_R_X75Y113_SLICE_X114Y113_AO6;
  assign CLBLL_R_X75Y113_SLICE_X114Y113_B = CLBLL_R_X75Y113_SLICE_X114Y113_BO6;
  assign CLBLL_R_X75Y113_SLICE_X114Y113_C = CLBLL_R_X75Y113_SLICE_X114Y113_CO6;
  assign CLBLL_R_X75Y113_SLICE_X114Y113_D = CLBLL_R_X75Y113_SLICE_X114Y113_DO6;
  assign CLBLL_R_X75Y113_SLICE_X115Y113_A = CLBLL_R_X75Y113_SLICE_X115Y113_AO6;
  assign CLBLL_R_X75Y113_SLICE_X115Y113_B = CLBLL_R_X75Y113_SLICE_X115Y113_BO6;
  assign CLBLL_R_X75Y113_SLICE_X115Y113_C = CLBLL_R_X75Y113_SLICE_X115Y113_CO6;
  assign CLBLL_R_X75Y113_SLICE_X115Y113_D = CLBLL_R_X75Y113_SLICE_X115Y113_DO6;
  assign CLBLL_R_X75Y121_SLICE_X114Y121_A = CLBLL_R_X75Y121_SLICE_X114Y121_AO6;
  assign CLBLL_R_X75Y121_SLICE_X114Y121_B = CLBLL_R_X75Y121_SLICE_X114Y121_BO6;
  assign CLBLL_R_X75Y121_SLICE_X114Y121_C = CLBLL_R_X75Y121_SLICE_X114Y121_CO6;
  assign CLBLL_R_X75Y121_SLICE_X114Y121_D = CLBLL_R_X75Y121_SLICE_X114Y121_DO6;
  assign CLBLL_R_X75Y121_SLICE_X114Y121_AMUX = CLBLL_R_X75Y121_SLICE_X114Y121_AO5;
  assign CLBLL_R_X75Y121_SLICE_X115Y121_A = CLBLL_R_X75Y121_SLICE_X115Y121_AO6;
  assign CLBLL_R_X75Y121_SLICE_X115Y121_B = CLBLL_R_X75Y121_SLICE_X115Y121_BO6;
  assign CLBLL_R_X75Y121_SLICE_X115Y121_C = CLBLL_R_X75Y121_SLICE_X115Y121_CO6;
  assign CLBLL_R_X75Y121_SLICE_X115Y121_D = CLBLL_R_X75Y121_SLICE_X115Y121_DO6;
  assign CLBLL_R_X75Y122_SLICE_X114Y122_A = CLBLL_R_X75Y122_SLICE_X114Y122_AO6;
  assign CLBLL_R_X75Y122_SLICE_X114Y122_B = CLBLL_R_X75Y122_SLICE_X114Y122_BO6;
  assign CLBLL_R_X75Y122_SLICE_X114Y122_C = CLBLL_R_X75Y122_SLICE_X114Y122_CO6;
  assign CLBLL_R_X75Y122_SLICE_X114Y122_D = CLBLL_R_X75Y122_SLICE_X114Y122_DO6;
  assign CLBLL_R_X75Y122_SLICE_X115Y122_A = CLBLL_R_X75Y122_SLICE_X115Y122_AO6;
  assign CLBLL_R_X75Y122_SLICE_X115Y122_B = CLBLL_R_X75Y122_SLICE_X115Y122_BO6;
  assign CLBLL_R_X75Y122_SLICE_X115Y122_C = CLBLL_R_X75Y122_SLICE_X115Y122_CO6;
  assign CLBLL_R_X75Y122_SLICE_X115Y122_D = CLBLL_R_X75Y122_SLICE_X115Y122_DO6;
  assign CLBLL_R_X75Y122_SLICE_X115Y122_AMUX = CLBLL_R_X75Y122_SLICE_X115Y122_A5Q;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_A = CLBLL_R_X75Y123_SLICE_X114Y123_AO6;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_B = CLBLL_R_X75Y123_SLICE_X114Y123_BO6;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_C = CLBLL_R_X75Y123_SLICE_X114Y123_CO6;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_D = CLBLL_R_X75Y123_SLICE_X114Y123_DO6;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_AMUX = CLBLL_R_X75Y123_SLICE_X114Y123_AO5;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_A = CLBLL_R_X75Y123_SLICE_X115Y123_AO6;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_B = CLBLL_R_X75Y123_SLICE_X115Y123_BO6;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_C = CLBLL_R_X75Y123_SLICE_X115Y123_CO6;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_D = CLBLL_R_X75Y123_SLICE_X115Y123_DO6;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_AMUX = CLBLL_R_X75Y123_SLICE_X115Y123_AO5;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_A = CLBLL_R_X75Y124_SLICE_X114Y124_AO6;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_B = CLBLL_R_X75Y124_SLICE_X114Y124_BO6;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_C = CLBLL_R_X75Y124_SLICE_X114Y124_CO6;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_D = CLBLL_R_X75Y124_SLICE_X114Y124_DO6;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_CMUX = CLBLL_R_X75Y124_SLICE_X114Y124_C5Q;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_DMUX = CLBLL_R_X75Y124_SLICE_X114Y124_D5Q;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_A = CLBLL_R_X75Y124_SLICE_X115Y124_AO6;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_B = CLBLL_R_X75Y124_SLICE_X115Y124_BO6;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_C = CLBLL_R_X75Y124_SLICE_X115Y124_CO6;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_D = CLBLL_R_X75Y124_SLICE_X115Y124_DO6;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_BMUX = CLBLL_R_X75Y124_SLICE_X115Y124_B5Q;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_A = CLBLL_R_X75Y127_SLICE_X114Y127_AO6;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_B = CLBLL_R_X75Y127_SLICE_X114Y127_BO6;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_C = CLBLL_R_X75Y127_SLICE_X114Y127_CO6;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_D = CLBLL_R_X75Y127_SLICE_X114Y127_DO6;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_AMUX = CLBLL_R_X75Y127_SLICE_X114Y127_A5Q;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_CMUX = CLBLL_R_X75Y127_SLICE_X114Y127_CO5;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_A = CLBLL_R_X75Y127_SLICE_X115Y127_AO6;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_B = CLBLL_R_X75Y127_SLICE_X115Y127_BO6;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_C = CLBLL_R_X75Y127_SLICE_X115Y127_CO6;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_D = CLBLL_R_X75Y127_SLICE_X115Y127_DO6;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_A = CLBLL_R_X75Y128_SLICE_X114Y128_AO6;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_B = CLBLL_R_X75Y128_SLICE_X114Y128_BO6;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_C = CLBLL_R_X75Y128_SLICE_X114Y128_CO6;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_D = CLBLL_R_X75Y128_SLICE_X114Y128_DO6;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_AMUX = CLBLL_R_X75Y128_SLICE_X114Y128_AO5;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_BMUX = CLBLL_R_X75Y128_SLICE_X114Y128_BO5;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_DMUX = CLBLL_R_X75Y128_SLICE_X114Y128_DO5;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_A = CLBLL_R_X75Y128_SLICE_X115Y128_AO6;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_B = CLBLL_R_X75Y128_SLICE_X115Y128_BO6;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_C = CLBLL_R_X75Y128_SLICE_X115Y128_CO6;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_D = CLBLL_R_X75Y128_SLICE_X115Y128_DO6;
  assign CLBLL_R_X75Y129_SLICE_X114Y129_A = CLBLL_R_X75Y129_SLICE_X114Y129_AO6;
  assign CLBLL_R_X75Y129_SLICE_X114Y129_B = CLBLL_R_X75Y129_SLICE_X114Y129_BO6;
  assign CLBLL_R_X75Y129_SLICE_X114Y129_C = CLBLL_R_X75Y129_SLICE_X114Y129_CO6;
  assign CLBLL_R_X75Y129_SLICE_X114Y129_D = CLBLL_R_X75Y129_SLICE_X114Y129_DO6;
  assign CLBLL_R_X75Y129_SLICE_X114Y129_CMUX = CLBLL_R_X75Y129_SLICE_X114Y129_CO5;
  assign CLBLL_R_X75Y129_SLICE_X115Y129_A = CLBLL_R_X75Y129_SLICE_X115Y129_AO6;
  assign CLBLL_R_X75Y129_SLICE_X115Y129_B = CLBLL_R_X75Y129_SLICE_X115Y129_BO6;
  assign CLBLL_R_X75Y129_SLICE_X115Y129_C = CLBLL_R_X75Y129_SLICE_X115Y129_CO6;
  assign CLBLL_R_X75Y129_SLICE_X115Y129_D = CLBLL_R_X75Y129_SLICE_X115Y129_DO6;
  assign CLBLL_R_X75Y130_SLICE_X114Y130_A = CLBLL_R_X75Y130_SLICE_X114Y130_AO6;
  assign CLBLL_R_X75Y130_SLICE_X114Y130_B = CLBLL_R_X75Y130_SLICE_X114Y130_BO6;
  assign CLBLL_R_X75Y130_SLICE_X114Y130_C = CLBLL_R_X75Y130_SLICE_X114Y130_CO6;
  assign CLBLL_R_X75Y130_SLICE_X114Y130_D = CLBLL_R_X75Y130_SLICE_X114Y130_DO6;
  assign CLBLL_R_X75Y130_SLICE_X115Y130_A = CLBLL_R_X75Y130_SLICE_X115Y130_AO6;
  assign CLBLL_R_X75Y130_SLICE_X115Y130_B = CLBLL_R_X75Y130_SLICE_X115Y130_BO6;
  assign CLBLL_R_X75Y130_SLICE_X115Y130_C = CLBLL_R_X75Y130_SLICE_X115Y130_CO6;
  assign CLBLL_R_X75Y130_SLICE_X115Y130_D = CLBLL_R_X75Y130_SLICE_X115Y130_DO6;
  assign CLBLL_R_X75Y130_SLICE_X115Y130_BMUX = CLBLL_R_X75Y130_SLICE_X115Y130_BO5;
  assign CLBLL_R_X75Y133_SLICE_X114Y133_A = CLBLL_R_X75Y133_SLICE_X114Y133_AO6;
  assign CLBLL_R_X75Y133_SLICE_X114Y133_B = CLBLL_R_X75Y133_SLICE_X114Y133_BO6;
  assign CLBLL_R_X75Y133_SLICE_X114Y133_C = CLBLL_R_X75Y133_SLICE_X114Y133_CO6;
  assign CLBLL_R_X75Y133_SLICE_X114Y133_D = CLBLL_R_X75Y133_SLICE_X114Y133_DO6;
  assign CLBLL_R_X75Y133_SLICE_X114Y133_CMUX = CLBLL_R_X75Y133_SLICE_X114Y133_CO5;
  assign CLBLL_R_X75Y133_SLICE_X115Y133_A = CLBLL_R_X75Y133_SLICE_X115Y133_AO6;
  assign CLBLL_R_X75Y133_SLICE_X115Y133_B = CLBLL_R_X75Y133_SLICE_X115Y133_BO6;
  assign CLBLL_R_X75Y133_SLICE_X115Y133_C = CLBLL_R_X75Y133_SLICE_X115Y133_CO6;
  assign CLBLL_R_X75Y133_SLICE_X115Y133_D = CLBLL_R_X75Y133_SLICE_X115Y133_DO6;
  assign CLBLL_R_X75Y134_SLICE_X114Y134_A = CLBLL_R_X75Y134_SLICE_X114Y134_AO6;
  assign CLBLL_R_X75Y134_SLICE_X114Y134_B = CLBLL_R_X75Y134_SLICE_X114Y134_BO6;
  assign CLBLL_R_X75Y134_SLICE_X114Y134_C = CLBLL_R_X75Y134_SLICE_X114Y134_CO6;
  assign CLBLL_R_X75Y134_SLICE_X114Y134_D = CLBLL_R_X75Y134_SLICE_X114Y134_DO6;
  assign CLBLL_R_X75Y134_SLICE_X114Y134_AMUX = CLBLL_R_X75Y134_SLICE_X114Y134_A5Q;
  assign CLBLL_R_X75Y134_SLICE_X114Y134_BMUX = CLBLL_R_X75Y134_SLICE_X114Y134_BO5;
  assign CLBLL_R_X75Y134_SLICE_X114Y134_CMUX = CLBLL_R_X75Y134_SLICE_X114Y134_CO5;
  assign CLBLL_R_X75Y134_SLICE_X115Y134_A = CLBLL_R_X75Y134_SLICE_X115Y134_AO6;
  assign CLBLL_R_X75Y134_SLICE_X115Y134_B = CLBLL_R_X75Y134_SLICE_X115Y134_BO6;
  assign CLBLL_R_X75Y134_SLICE_X115Y134_C = CLBLL_R_X75Y134_SLICE_X115Y134_CO6;
  assign CLBLL_R_X75Y134_SLICE_X115Y134_D = CLBLL_R_X75Y134_SLICE_X115Y134_DO6;
  assign CLBLL_R_X75Y134_SLICE_X115Y134_AMUX = CLBLL_R_X75Y134_SLICE_X115Y134_AO5;
  assign CLBLL_R_X75Y134_SLICE_X115Y134_DMUX = CLBLL_R_X75Y134_SLICE_X115Y134_DO5;
  assign CLBLL_R_X77Y104_SLICE_X118Y104_A = CLBLL_R_X77Y104_SLICE_X118Y104_AO6;
  assign CLBLL_R_X77Y104_SLICE_X118Y104_B = CLBLL_R_X77Y104_SLICE_X118Y104_BO6;
  assign CLBLL_R_X77Y104_SLICE_X118Y104_C = CLBLL_R_X77Y104_SLICE_X118Y104_CO6;
  assign CLBLL_R_X77Y104_SLICE_X118Y104_D = CLBLL_R_X77Y104_SLICE_X118Y104_DO6;
  assign CLBLL_R_X77Y104_SLICE_X119Y104_A = CLBLL_R_X77Y104_SLICE_X119Y104_AO6;
  assign CLBLL_R_X77Y104_SLICE_X119Y104_B = CLBLL_R_X77Y104_SLICE_X119Y104_BO6;
  assign CLBLL_R_X77Y104_SLICE_X119Y104_C = CLBLL_R_X77Y104_SLICE_X119Y104_CO6;
  assign CLBLL_R_X77Y104_SLICE_X119Y104_D = CLBLL_R_X77Y104_SLICE_X119Y104_DO6;
  assign CLBLL_R_X77Y104_SLICE_X119Y104_AMUX = CLBLL_R_X77Y104_SLICE_X119Y104_A5Q;
  assign CLBLL_R_X77Y108_SLICE_X118Y108_A = CLBLL_R_X77Y108_SLICE_X118Y108_AO6;
  assign CLBLL_R_X77Y108_SLICE_X118Y108_B = CLBLL_R_X77Y108_SLICE_X118Y108_BO6;
  assign CLBLL_R_X77Y108_SLICE_X118Y108_C = CLBLL_R_X77Y108_SLICE_X118Y108_CO6;
  assign CLBLL_R_X77Y108_SLICE_X118Y108_D = CLBLL_R_X77Y108_SLICE_X118Y108_DO6;
  assign CLBLL_R_X77Y108_SLICE_X119Y108_A = CLBLL_R_X77Y108_SLICE_X119Y108_AO6;
  assign CLBLL_R_X77Y108_SLICE_X119Y108_B = CLBLL_R_X77Y108_SLICE_X119Y108_BO6;
  assign CLBLL_R_X77Y108_SLICE_X119Y108_C = CLBLL_R_X77Y108_SLICE_X119Y108_CO6;
  assign CLBLL_R_X77Y108_SLICE_X119Y108_D = CLBLL_R_X77Y108_SLICE_X119Y108_DO6;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_A = CLBLL_R_X77Y113_SLICE_X118Y113_AO6;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_B = CLBLL_R_X77Y113_SLICE_X118Y113_BO6;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_C = CLBLL_R_X77Y113_SLICE_X118Y113_CO6;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_D = CLBLL_R_X77Y113_SLICE_X118Y113_DO6;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_A = CLBLL_R_X77Y113_SLICE_X119Y113_AO6;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_B = CLBLL_R_X77Y113_SLICE_X119Y113_BO6;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_C = CLBLL_R_X77Y113_SLICE_X119Y113_CO6;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_D = CLBLL_R_X77Y113_SLICE_X119Y113_DO6;
  assign CLBLL_R_X77Y121_SLICE_X118Y121_A = CLBLL_R_X77Y121_SLICE_X118Y121_AO6;
  assign CLBLL_R_X77Y121_SLICE_X118Y121_B = CLBLL_R_X77Y121_SLICE_X118Y121_BO6;
  assign CLBLL_R_X77Y121_SLICE_X118Y121_C = CLBLL_R_X77Y121_SLICE_X118Y121_CO6;
  assign CLBLL_R_X77Y121_SLICE_X118Y121_D = CLBLL_R_X77Y121_SLICE_X118Y121_DO6;
  assign CLBLL_R_X77Y121_SLICE_X119Y121_A = CLBLL_R_X77Y121_SLICE_X119Y121_AO6;
  assign CLBLL_R_X77Y121_SLICE_X119Y121_B = CLBLL_R_X77Y121_SLICE_X119Y121_BO6;
  assign CLBLL_R_X77Y121_SLICE_X119Y121_C = CLBLL_R_X77Y121_SLICE_X119Y121_CO6;
  assign CLBLL_R_X77Y121_SLICE_X119Y121_D = CLBLL_R_X77Y121_SLICE_X119Y121_DO6;
  assign CLBLL_R_X77Y121_SLICE_X119Y121_BMUX = CLBLL_R_X77Y121_SLICE_X119Y121_BO5;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_A = CLBLL_R_X77Y122_SLICE_X118Y122_AO6;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_B = CLBLL_R_X77Y122_SLICE_X118Y122_BO6;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_C = CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_D = CLBLL_R_X77Y122_SLICE_X118Y122_DO6;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_A = CLBLL_R_X77Y122_SLICE_X119Y122_AO6;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_B = CLBLL_R_X77Y122_SLICE_X119Y122_BO6;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_C = CLBLL_R_X77Y122_SLICE_X119Y122_CO6;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_D = CLBLL_R_X77Y122_SLICE_X119Y122_DO6;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_AMUX = CLBLL_R_X77Y122_SLICE_X119Y122_AO5;
  assign CLBLL_R_X77Y123_SLICE_X118Y123_A = CLBLL_R_X77Y123_SLICE_X118Y123_AO6;
  assign CLBLL_R_X77Y123_SLICE_X118Y123_B = CLBLL_R_X77Y123_SLICE_X118Y123_BO6;
  assign CLBLL_R_X77Y123_SLICE_X118Y123_C = CLBLL_R_X77Y123_SLICE_X118Y123_CO6;
  assign CLBLL_R_X77Y123_SLICE_X118Y123_D = CLBLL_R_X77Y123_SLICE_X118Y123_DO6;
  assign CLBLL_R_X77Y123_SLICE_X118Y123_BMUX = CLBLL_R_X77Y123_SLICE_X118Y123_BO5;
  assign CLBLL_R_X77Y123_SLICE_X119Y123_A = CLBLL_R_X77Y123_SLICE_X119Y123_AO6;
  assign CLBLL_R_X77Y123_SLICE_X119Y123_B = CLBLL_R_X77Y123_SLICE_X119Y123_BO6;
  assign CLBLL_R_X77Y123_SLICE_X119Y123_C = CLBLL_R_X77Y123_SLICE_X119Y123_CO6;
  assign CLBLL_R_X77Y123_SLICE_X119Y123_D = CLBLL_R_X77Y123_SLICE_X119Y123_DO6;
  assign CLBLL_R_X77Y123_SLICE_X119Y123_BMUX = CLBLL_R_X77Y123_SLICE_X119Y123_BO5;
  assign CLBLL_R_X77Y124_SLICE_X118Y124_A = CLBLL_R_X77Y124_SLICE_X118Y124_AO6;
  assign CLBLL_R_X77Y124_SLICE_X118Y124_B = CLBLL_R_X77Y124_SLICE_X118Y124_BO6;
  assign CLBLL_R_X77Y124_SLICE_X118Y124_C = CLBLL_R_X77Y124_SLICE_X118Y124_CO6;
  assign CLBLL_R_X77Y124_SLICE_X118Y124_D = CLBLL_R_X77Y124_SLICE_X118Y124_DO6;
  assign CLBLL_R_X77Y124_SLICE_X118Y124_AMUX = CLBLL_R_X77Y124_SLICE_X118Y124_AO5;
  assign CLBLL_R_X77Y124_SLICE_X119Y124_A = CLBLL_R_X77Y124_SLICE_X119Y124_AO6;
  assign CLBLL_R_X77Y124_SLICE_X119Y124_B = CLBLL_R_X77Y124_SLICE_X119Y124_BO6;
  assign CLBLL_R_X77Y124_SLICE_X119Y124_C = CLBLL_R_X77Y124_SLICE_X119Y124_CO6;
  assign CLBLL_R_X77Y124_SLICE_X119Y124_D = CLBLL_R_X77Y124_SLICE_X119Y124_DO6;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_A = CLBLL_R_X77Y125_SLICE_X118Y125_AO6;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_B = CLBLL_R_X77Y125_SLICE_X118Y125_BO6;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_C = CLBLL_R_X77Y125_SLICE_X118Y125_CO6;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_D = CLBLL_R_X77Y125_SLICE_X118Y125_DO6;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_AMUX = CLBLL_R_X77Y125_SLICE_X118Y125_A5Q;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_BMUX = CLBLL_R_X77Y125_SLICE_X118Y125_BO5;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_A = CLBLL_R_X77Y125_SLICE_X119Y125_AO6;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_B = CLBLL_R_X77Y125_SLICE_X119Y125_BO6;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_C = CLBLL_R_X77Y125_SLICE_X119Y125_CO6;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_D = CLBLL_R_X77Y125_SLICE_X119Y125_DO6;
  assign CLBLL_R_X77Y126_SLICE_X118Y126_A = CLBLL_R_X77Y126_SLICE_X118Y126_AO6;
  assign CLBLL_R_X77Y126_SLICE_X118Y126_B = CLBLL_R_X77Y126_SLICE_X118Y126_BO6;
  assign CLBLL_R_X77Y126_SLICE_X118Y126_C = CLBLL_R_X77Y126_SLICE_X118Y126_CO6;
  assign CLBLL_R_X77Y126_SLICE_X118Y126_D = CLBLL_R_X77Y126_SLICE_X118Y126_DO6;
  assign CLBLL_R_X77Y126_SLICE_X118Y126_AMUX = CLBLL_R_X77Y126_SLICE_X118Y126_AO5;
  assign CLBLL_R_X77Y126_SLICE_X119Y126_A = CLBLL_R_X77Y126_SLICE_X119Y126_AO6;
  assign CLBLL_R_X77Y126_SLICE_X119Y126_B = CLBLL_R_X77Y126_SLICE_X119Y126_BO6;
  assign CLBLL_R_X77Y126_SLICE_X119Y126_C = CLBLL_R_X77Y126_SLICE_X119Y126_CO6;
  assign CLBLL_R_X77Y126_SLICE_X119Y126_D = CLBLL_R_X77Y126_SLICE_X119Y126_DO6;
  assign CLBLL_R_X77Y127_SLICE_X118Y127_A = CLBLL_R_X77Y127_SLICE_X118Y127_AO6;
  assign CLBLL_R_X77Y127_SLICE_X118Y127_B = CLBLL_R_X77Y127_SLICE_X118Y127_BO6;
  assign CLBLL_R_X77Y127_SLICE_X118Y127_C = CLBLL_R_X77Y127_SLICE_X118Y127_CO6;
  assign CLBLL_R_X77Y127_SLICE_X118Y127_D = CLBLL_R_X77Y127_SLICE_X118Y127_DO6;
  assign CLBLL_R_X77Y127_SLICE_X119Y127_A = CLBLL_R_X77Y127_SLICE_X119Y127_AO6;
  assign CLBLL_R_X77Y127_SLICE_X119Y127_B = CLBLL_R_X77Y127_SLICE_X119Y127_BO6;
  assign CLBLL_R_X77Y127_SLICE_X119Y127_C = CLBLL_R_X77Y127_SLICE_X119Y127_CO6;
  assign CLBLL_R_X77Y127_SLICE_X119Y127_D = CLBLL_R_X77Y127_SLICE_X119Y127_DO6;
  assign CLBLL_R_X77Y127_SLICE_X119Y127_AMUX = CLBLL_R_X77Y127_SLICE_X119Y127_AO5;
  assign CLBLL_R_X77Y128_SLICE_X118Y128_A = CLBLL_R_X77Y128_SLICE_X118Y128_AO6;
  assign CLBLL_R_X77Y128_SLICE_X118Y128_B = CLBLL_R_X77Y128_SLICE_X118Y128_BO6;
  assign CLBLL_R_X77Y128_SLICE_X118Y128_C = CLBLL_R_X77Y128_SLICE_X118Y128_CO6;
  assign CLBLL_R_X77Y128_SLICE_X118Y128_D = CLBLL_R_X77Y128_SLICE_X118Y128_DO6;
  assign CLBLL_R_X77Y128_SLICE_X118Y128_AMUX = CLBLL_R_X77Y128_SLICE_X118Y128_AO5;
  assign CLBLL_R_X77Y128_SLICE_X118Y128_BMUX = CLBLL_R_X77Y128_SLICE_X118Y128_B5Q;
  assign CLBLL_R_X77Y128_SLICE_X118Y128_CMUX = CLBLL_R_X77Y128_SLICE_X118Y128_CO5;
  assign CLBLL_R_X77Y128_SLICE_X119Y128_A = CLBLL_R_X77Y128_SLICE_X119Y128_AO6;
  assign CLBLL_R_X77Y128_SLICE_X119Y128_B = CLBLL_R_X77Y128_SLICE_X119Y128_BO6;
  assign CLBLL_R_X77Y128_SLICE_X119Y128_C = CLBLL_R_X77Y128_SLICE_X119Y128_CO6;
  assign CLBLL_R_X77Y128_SLICE_X119Y128_D = CLBLL_R_X77Y128_SLICE_X119Y128_DO6;
  assign CLBLL_R_X77Y128_SLICE_X119Y128_AMUX = CLBLL_R_X77Y128_SLICE_X119Y128_A5Q;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_A = CLBLL_R_X77Y129_SLICE_X118Y129_AO6;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_B = CLBLL_R_X77Y129_SLICE_X118Y129_BO6;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_C = CLBLL_R_X77Y129_SLICE_X118Y129_CO6;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_D = CLBLL_R_X77Y129_SLICE_X118Y129_DO6;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_A = CLBLL_R_X77Y129_SLICE_X119Y129_AO6;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_B = CLBLL_R_X77Y129_SLICE_X119Y129_BO6;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_C = CLBLL_R_X77Y129_SLICE_X119Y129_CO6;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_D = CLBLL_R_X77Y129_SLICE_X119Y129_DO6;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_AMUX = CLBLL_R_X77Y129_SLICE_X119Y129_AO5;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_CMUX = CLBLL_R_X77Y129_SLICE_X119Y129_CO6;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_A = CLBLL_R_X77Y130_SLICE_X118Y130_AO6;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_B = CLBLL_R_X77Y130_SLICE_X118Y130_BO6;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_C = CLBLL_R_X77Y130_SLICE_X118Y130_CO6;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_D = CLBLL_R_X77Y130_SLICE_X118Y130_DO6;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_AMUX = CLBLL_R_X77Y130_SLICE_X118Y130_AO5;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_DMUX = CLBLL_R_X77Y130_SLICE_X118Y130_DO5;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_A = CLBLL_R_X77Y130_SLICE_X119Y130_AO6;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_B = CLBLL_R_X77Y130_SLICE_X119Y130_BO6;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_C = CLBLL_R_X77Y130_SLICE_X119Y130_CO6;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_D = CLBLL_R_X77Y130_SLICE_X119Y130_DO6;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_AMUX = CLBLL_R_X77Y130_SLICE_X119Y130_AO5;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_A = CLBLL_R_X77Y131_SLICE_X118Y131_AO6;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_B = CLBLL_R_X77Y131_SLICE_X118Y131_BO6;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_C = CLBLL_R_X77Y131_SLICE_X118Y131_CO6;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_D = CLBLL_R_X77Y131_SLICE_X118Y131_DO6;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_A = CLBLL_R_X77Y131_SLICE_X119Y131_AO6;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_B = CLBLL_R_X77Y131_SLICE_X119Y131_BO6;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_C = CLBLL_R_X77Y131_SLICE_X119Y131_CO6;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_D = CLBLL_R_X77Y131_SLICE_X119Y131_DO6;
  assign CLBLL_R_X79Y96_SLICE_X122Y96_A = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLL_R_X79Y96_SLICE_X122Y96_B = CLBLL_R_X79Y96_SLICE_X122Y96_BO6;
  assign CLBLL_R_X79Y96_SLICE_X122Y96_C = CLBLL_R_X79Y96_SLICE_X122Y96_CO6;
  assign CLBLL_R_X79Y96_SLICE_X122Y96_D = CLBLL_R_X79Y96_SLICE_X122Y96_DO6;
  assign CLBLL_R_X79Y96_SLICE_X123Y96_A = CLBLL_R_X79Y96_SLICE_X123Y96_AO6;
  assign CLBLL_R_X79Y96_SLICE_X123Y96_B = CLBLL_R_X79Y96_SLICE_X123Y96_BO6;
  assign CLBLL_R_X79Y96_SLICE_X123Y96_C = CLBLL_R_X79Y96_SLICE_X123Y96_CO6;
  assign CLBLL_R_X79Y96_SLICE_X123Y96_D = CLBLL_R_X79Y96_SLICE_X123Y96_DO6;
  assign CLBLL_R_X79Y99_SLICE_X122Y99_A = CLBLL_R_X79Y99_SLICE_X122Y99_AO6;
  assign CLBLL_R_X79Y99_SLICE_X122Y99_B = CLBLL_R_X79Y99_SLICE_X122Y99_BO6;
  assign CLBLL_R_X79Y99_SLICE_X122Y99_C = CLBLL_R_X79Y99_SLICE_X122Y99_CO6;
  assign CLBLL_R_X79Y99_SLICE_X122Y99_D = CLBLL_R_X79Y99_SLICE_X122Y99_DO6;
  assign CLBLL_R_X79Y99_SLICE_X123Y99_A = CLBLL_R_X79Y99_SLICE_X123Y99_AO6;
  assign CLBLL_R_X79Y99_SLICE_X123Y99_B = CLBLL_R_X79Y99_SLICE_X123Y99_BO6;
  assign CLBLL_R_X79Y99_SLICE_X123Y99_C = CLBLL_R_X79Y99_SLICE_X123Y99_CO6;
  assign CLBLL_R_X79Y99_SLICE_X123Y99_D = CLBLL_R_X79Y99_SLICE_X123Y99_DO6;
  assign CLBLL_R_X79Y104_SLICE_X122Y104_A = CLBLL_R_X79Y104_SLICE_X122Y104_AO6;
  assign CLBLL_R_X79Y104_SLICE_X122Y104_B = CLBLL_R_X79Y104_SLICE_X122Y104_BO6;
  assign CLBLL_R_X79Y104_SLICE_X122Y104_C = CLBLL_R_X79Y104_SLICE_X122Y104_CO6;
  assign CLBLL_R_X79Y104_SLICE_X122Y104_D = CLBLL_R_X79Y104_SLICE_X122Y104_DO6;
  assign CLBLL_R_X79Y104_SLICE_X122Y104_AMUX = CLBLL_R_X79Y104_SLICE_X122Y104_A5Q;
  assign CLBLL_R_X79Y104_SLICE_X123Y104_A = CLBLL_R_X79Y104_SLICE_X123Y104_AO6;
  assign CLBLL_R_X79Y104_SLICE_X123Y104_B = CLBLL_R_X79Y104_SLICE_X123Y104_BO6;
  assign CLBLL_R_X79Y104_SLICE_X123Y104_C = CLBLL_R_X79Y104_SLICE_X123Y104_CO6;
  assign CLBLL_R_X79Y104_SLICE_X123Y104_D = CLBLL_R_X79Y104_SLICE_X123Y104_DO6;
  assign CLBLL_R_X79Y127_SLICE_X122Y127_A = CLBLL_R_X79Y127_SLICE_X122Y127_AO6;
  assign CLBLL_R_X79Y127_SLICE_X122Y127_B = CLBLL_R_X79Y127_SLICE_X122Y127_BO6;
  assign CLBLL_R_X79Y127_SLICE_X122Y127_C = CLBLL_R_X79Y127_SLICE_X122Y127_CO6;
  assign CLBLL_R_X79Y127_SLICE_X122Y127_D = CLBLL_R_X79Y127_SLICE_X122Y127_DO6;
  assign CLBLL_R_X79Y127_SLICE_X122Y127_AMUX = CLBLL_R_X79Y127_SLICE_X122Y127_A5Q;
  assign CLBLL_R_X79Y127_SLICE_X123Y127_A = CLBLL_R_X79Y127_SLICE_X123Y127_AO6;
  assign CLBLL_R_X79Y127_SLICE_X123Y127_B = CLBLL_R_X79Y127_SLICE_X123Y127_BO6;
  assign CLBLL_R_X79Y127_SLICE_X123Y127_C = CLBLL_R_X79Y127_SLICE_X123Y127_CO6;
  assign CLBLL_R_X79Y127_SLICE_X123Y127_D = CLBLL_R_X79Y127_SLICE_X123Y127_DO6;
  assign CLBLL_R_X79Y128_SLICE_X122Y128_A = CLBLL_R_X79Y128_SLICE_X122Y128_AO6;
  assign CLBLL_R_X79Y128_SLICE_X122Y128_B = CLBLL_R_X79Y128_SLICE_X122Y128_BO6;
  assign CLBLL_R_X79Y128_SLICE_X122Y128_C = CLBLL_R_X79Y128_SLICE_X122Y128_CO6;
  assign CLBLL_R_X79Y128_SLICE_X122Y128_D = CLBLL_R_X79Y128_SLICE_X122Y128_DO6;
  assign CLBLL_R_X79Y128_SLICE_X123Y128_A = CLBLL_R_X79Y128_SLICE_X123Y128_AO6;
  assign CLBLL_R_X79Y128_SLICE_X123Y128_B = CLBLL_R_X79Y128_SLICE_X123Y128_BO6;
  assign CLBLL_R_X79Y128_SLICE_X123Y128_C = CLBLL_R_X79Y128_SLICE_X123Y128_CO6;
  assign CLBLL_R_X79Y128_SLICE_X123Y128_D = CLBLL_R_X79Y128_SLICE_X123Y128_DO6;
  assign CLBLL_R_X79Y135_SLICE_X122Y135_A = CLBLL_R_X79Y135_SLICE_X122Y135_AO6;
  assign CLBLL_R_X79Y135_SLICE_X122Y135_B = CLBLL_R_X79Y135_SLICE_X122Y135_BO6;
  assign CLBLL_R_X79Y135_SLICE_X122Y135_C = CLBLL_R_X79Y135_SLICE_X122Y135_CO6;
  assign CLBLL_R_X79Y135_SLICE_X122Y135_D = CLBLL_R_X79Y135_SLICE_X122Y135_DO6;
  assign CLBLL_R_X79Y135_SLICE_X123Y135_A = CLBLL_R_X79Y135_SLICE_X123Y135_AO6;
  assign CLBLL_R_X79Y135_SLICE_X123Y135_B = CLBLL_R_X79Y135_SLICE_X123Y135_BO6;
  assign CLBLL_R_X79Y135_SLICE_X123Y135_C = CLBLL_R_X79Y135_SLICE_X123Y135_CO6;
  assign CLBLL_R_X79Y135_SLICE_X123Y135_D = CLBLL_R_X79Y135_SLICE_X123Y135_DO6;
  assign CLBLL_R_X83Y94_SLICE_X130Y94_A = CLBLL_R_X83Y94_SLICE_X130Y94_AO6;
  assign CLBLL_R_X83Y94_SLICE_X130Y94_B = CLBLL_R_X83Y94_SLICE_X130Y94_BO6;
  assign CLBLL_R_X83Y94_SLICE_X130Y94_C = CLBLL_R_X83Y94_SLICE_X130Y94_CO6;
  assign CLBLL_R_X83Y94_SLICE_X130Y94_D = CLBLL_R_X83Y94_SLICE_X130Y94_DO6;
  assign CLBLL_R_X83Y94_SLICE_X130Y94_AMUX = CLBLL_R_X83Y94_SLICE_X130Y94_A5Q;
  assign CLBLL_R_X83Y94_SLICE_X131Y94_A = CLBLL_R_X83Y94_SLICE_X131Y94_AO6;
  assign CLBLL_R_X83Y94_SLICE_X131Y94_B = CLBLL_R_X83Y94_SLICE_X131Y94_BO6;
  assign CLBLL_R_X83Y94_SLICE_X131Y94_C = CLBLL_R_X83Y94_SLICE_X131Y94_CO6;
  assign CLBLL_R_X83Y94_SLICE_X131Y94_D = CLBLL_R_X83Y94_SLICE_X131Y94_DO6;
  assign CLBLL_R_X83Y130_SLICE_X130Y130_A = CLBLL_R_X83Y130_SLICE_X130Y130_AO6;
  assign CLBLL_R_X83Y130_SLICE_X130Y130_B = CLBLL_R_X83Y130_SLICE_X130Y130_BO6;
  assign CLBLL_R_X83Y130_SLICE_X130Y130_C = CLBLL_R_X83Y130_SLICE_X130Y130_CO6;
  assign CLBLL_R_X83Y130_SLICE_X130Y130_D = CLBLL_R_X83Y130_SLICE_X130Y130_DO6;
  assign CLBLL_R_X83Y130_SLICE_X131Y130_A = CLBLL_R_X83Y130_SLICE_X131Y130_AO6;
  assign CLBLL_R_X83Y130_SLICE_X131Y130_B = CLBLL_R_X83Y130_SLICE_X131Y130_BO6;
  assign CLBLL_R_X83Y130_SLICE_X131Y130_C = CLBLL_R_X83Y130_SLICE_X131Y130_CO6;
  assign CLBLL_R_X83Y130_SLICE_X131Y130_D = CLBLL_R_X83Y130_SLICE_X131Y130_DO6;
  assign CLBLL_R_X83Y132_SLICE_X130Y132_A = CLBLL_R_X83Y132_SLICE_X130Y132_AO6;
  assign CLBLL_R_X83Y132_SLICE_X130Y132_B = CLBLL_R_X83Y132_SLICE_X130Y132_BO6;
  assign CLBLL_R_X83Y132_SLICE_X130Y132_C = CLBLL_R_X83Y132_SLICE_X130Y132_CO6;
  assign CLBLL_R_X83Y132_SLICE_X130Y132_D = CLBLL_R_X83Y132_SLICE_X130Y132_DO6;
  assign CLBLL_R_X83Y132_SLICE_X131Y132_A = CLBLL_R_X83Y132_SLICE_X131Y132_AO6;
  assign CLBLL_R_X83Y132_SLICE_X131Y132_B = CLBLL_R_X83Y132_SLICE_X131Y132_BO6;
  assign CLBLL_R_X83Y132_SLICE_X131Y132_C = CLBLL_R_X83Y132_SLICE_X131Y132_CO6;
  assign CLBLL_R_X83Y132_SLICE_X131Y132_D = CLBLL_R_X83Y132_SLICE_X131Y132_DO6;
  assign CLBLM_L_X60Y92_SLICE_X90Y92_A = CLBLM_L_X60Y92_SLICE_X90Y92_AO6;
  assign CLBLM_L_X60Y92_SLICE_X90Y92_B = CLBLM_L_X60Y92_SLICE_X90Y92_BO6;
  assign CLBLM_L_X60Y92_SLICE_X90Y92_C = CLBLM_L_X60Y92_SLICE_X90Y92_CO6;
  assign CLBLM_L_X60Y92_SLICE_X90Y92_D = CLBLM_L_X60Y92_SLICE_X90Y92_DO6;
  assign CLBLM_L_X60Y92_SLICE_X91Y92_A = CLBLM_L_X60Y92_SLICE_X91Y92_AO6;
  assign CLBLM_L_X60Y92_SLICE_X91Y92_B = CLBLM_L_X60Y92_SLICE_X91Y92_BO6;
  assign CLBLM_L_X60Y92_SLICE_X91Y92_C = CLBLM_L_X60Y92_SLICE_X91Y92_CO6;
  assign CLBLM_L_X60Y92_SLICE_X91Y92_D = CLBLM_L_X60Y92_SLICE_X91Y92_DO6;
  assign CLBLM_L_X60Y94_SLICE_X90Y94_A = CLBLM_L_X60Y94_SLICE_X90Y94_AO6;
  assign CLBLM_L_X60Y94_SLICE_X90Y94_B = CLBLM_L_X60Y94_SLICE_X90Y94_BO6;
  assign CLBLM_L_X60Y94_SLICE_X90Y94_C = CLBLM_L_X60Y94_SLICE_X90Y94_CO6;
  assign CLBLM_L_X60Y94_SLICE_X90Y94_D = CLBLM_L_X60Y94_SLICE_X90Y94_DO6;
  assign CLBLM_L_X60Y94_SLICE_X91Y94_A = CLBLM_L_X60Y94_SLICE_X91Y94_AO6;
  assign CLBLM_L_X60Y94_SLICE_X91Y94_B = CLBLM_L_X60Y94_SLICE_X91Y94_BO6;
  assign CLBLM_L_X60Y94_SLICE_X91Y94_C = CLBLM_L_X60Y94_SLICE_X91Y94_CO6;
  assign CLBLM_L_X60Y94_SLICE_X91Y94_D = CLBLM_L_X60Y94_SLICE_X91Y94_DO6;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_A = CLBLM_L_X60Y97_SLICE_X90Y97_AO6;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_B = CLBLM_L_X60Y97_SLICE_X90Y97_BO6;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_C = CLBLM_L_X60Y97_SLICE_X90Y97_CO6;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_D = CLBLM_L_X60Y97_SLICE_X90Y97_DO6;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_A = CLBLM_L_X60Y97_SLICE_X91Y97_AO6;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_B = CLBLM_L_X60Y97_SLICE_X91Y97_BO6;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_C = CLBLM_L_X60Y97_SLICE_X91Y97_CO6;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_D = CLBLM_L_X60Y97_SLICE_X91Y97_DO6;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_A = CLBLM_L_X60Y99_SLICE_X90Y99_AO6;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_B = CLBLM_L_X60Y99_SLICE_X90Y99_BO6;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_C = CLBLM_L_X60Y99_SLICE_X90Y99_CO6;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_D = CLBLM_L_X60Y99_SLICE_X90Y99_DO6;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_A = CLBLM_L_X60Y99_SLICE_X91Y99_AO6;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_B = CLBLM_L_X60Y99_SLICE_X91Y99_BO6;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_C = CLBLM_L_X60Y99_SLICE_X91Y99_CO6;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_D = CLBLM_L_X60Y99_SLICE_X91Y99_DO6;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_A = CLBLM_L_X60Y101_SLICE_X90Y101_AO6;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_B = CLBLM_L_X60Y101_SLICE_X90Y101_BO6;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_C = CLBLM_L_X60Y101_SLICE_X90Y101_CO6;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_D = CLBLM_L_X60Y101_SLICE_X90Y101_DO6;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_A = CLBLM_L_X60Y101_SLICE_X91Y101_AO6;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_B = CLBLM_L_X60Y101_SLICE_X91Y101_BO6;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_C = CLBLM_L_X60Y101_SLICE_X91Y101_CO6;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_D = CLBLM_L_X60Y101_SLICE_X91Y101_DO6;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_A = CLBLM_L_X60Y104_SLICE_X90Y104_AO6;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_B = CLBLM_L_X60Y104_SLICE_X90Y104_BO6;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_C = CLBLM_L_X60Y104_SLICE_X90Y104_CO6;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_D = CLBLM_L_X60Y104_SLICE_X90Y104_DO6;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_A = CLBLM_L_X60Y104_SLICE_X91Y104_AO6;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_B = CLBLM_L_X60Y104_SLICE_X91Y104_BO6;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_C = CLBLM_L_X60Y104_SLICE_X91Y104_CO6;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_D = CLBLM_L_X60Y104_SLICE_X91Y104_DO6;
  assign CLBLM_L_X62Y90_SLICE_X92Y90_A = CLBLM_L_X62Y90_SLICE_X92Y90_AO6;
  assign CLBLM_L_X62Y90_SLICE_X92Y90_B = CLBLM_L_X62Y90_SLICE_X92Y90_BO6;
  assign CLBLM_L_X62Y90_SLICE_X92Y90_C = CLBLM_L_X62Y90_SLICE_X92Y90_CO6;
  assign CLBLM_L_X62Y90_SLICE_X92Y90_D = CLBLM_L_X62Y90_SLICE_X92Y90_DO6;
  assign CLBLM_L_X62Y90_SLICE_X93Y90_A = CLBLM_L_X62Y90_SLICE_X93Y90_AO6;
  assign CLBLM_L_X62Y90_SLICE_X93Y90_B = CLBLM_L_X62Y90_SLICE_X93Y90_BO6;
  assign CLBLM_L_X62Y90_SLICE_X93Y90_C = CLBLM_L_X62Y90_SLICE_X93Y90_CO6;
  assign CLBLM_L_X62Y90_SLICE_X93Y90_D = CLBLM_L_X62Y90_SLICE_X93Y90_DO6;
  assign CLBLM_L_X62Y92_SLICE_X92Y92_A = CLBLM_L_X62Y92_SLICE_X92Y92_AO6;
  assign CLBLM_L_X62Y92_SLICE_X92Y92_B = CLBLM_L_X62Y92_SLICE_X92Y92_BO6;
  assign CLBLM_L_X62Y92_SLICE_X92Y92_C = CLBLM_L_X62Y92_SLICE_X92Y92_CO6;
  assign CLBLM_L_X62Y92_SLICE_X92Y92_D = CLBLM_L_X62Y92_SLICE_X92Y92_DO6;
  assign CLBLM_L_X62Y92_SLICE_X93Y92_A = CLBLM_L_X62Y92_SLICE_X93Y92_AO6;
  assign CLBLM_L_X62Y92_SLICE_X93Y92_B = CLBLM_L_X62Y92_SLICE_X93Y92_BO6;
  assign CLBLM_L_X62Y92_SLICE_X93Y92_C = CLBLM_L_X62Y92_SLICE_X93Y92_CO6;
  assign CLBLM_L_X62Y92_SLICE_X93Y92_D = CLBLM_L_X62Y92_SLICE_X93Y92_DO6;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_A = CLBLM_L_X62Y95_SLICE_X92Y95_AO6;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_B = CLBLM_L_X62Y95_SLICE_X92Y95_BO6;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_C = CLBLM_L_X62Y95_SLICE_X92Y95_CO6;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_D = CLBLM_L_X62Y95_SLICE_X92Y95_DO6;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_A = CLBLM_L_X62Y95_SLICE_X93Y95_AO6;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_B = CLBLM_L_X62Y95_SLICE_X93Y95_BO6;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_C = CLBLM_L_X62Y95_SLICE_X93Y95_CO6;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_D = CLBLM_L_X62Y95_SLICE_X93Y95_DO6;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_A = CLBLM_L_X62Y97_SLICE_X92Y97_AO6;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_B = CLBLM_L_X62Y97_SLICE_X92Y97_BO6;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_C = CLBLM_L_X62Y97_SLICE_X92Y97_CO6;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_D = CLBLM_L_X62Y97_SLICE_X92Y97_DO6;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_A = CLBLM_L_X62Y97_SLICE_X93Y97_AO6;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_B = CLBLM_L_X62Y97_SLICE_X93Y97_BO6;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_C = CLBLM_L_X62Y97_SLICE_X93Y97_CO6;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_D = CLBLM_L_X62Y97_SLICE_X93Y97_DO6;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_A = CLBLM_L_X62Y98_SLICE_X92Y98_AO6;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_B = CLBLM_L_X62Y98_SLICE_X92Y98_BO6;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_C = CLBLM_L_X62Y98_SLICE_X92Y98_CO6;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_D = CLBLM_L_X62Y98_SLICE_X92Y98_DO6;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_A = CLBLM_L_X62Y98_SLICE_X93Y98_AO6;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_B = CLBLM_L_X62Y98_SLICE_X93Y98_BO6;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_C = CLBLM_L_X62Y98_SLICE_X93Y98_CO6;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_D = CLBLM_L_X62Y98_SLICE_X93Y98_DO6;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_A = CLBLM_L_X62Y99_SLICE_X92Y99_AO6;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_B = CLBLM_L_X62Y99_SLICE_X92Y99_BO6;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_C = CLBLM_L_X62Y99_SLICE_X92Y99_CO6;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_D = CLBLM_L_X62Y99_SLICE_X92Y99_DO6;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_A = CLBLM_L_X62Y99_SLICE_X93Y99_AO6;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_B = CLBLM_L_X62Y99_SLICE_X93Y99_BO6;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_C = CLBLM_L_X62Y99_SLICE_X93Y99_CO6;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_D = CLBLM_L_X62Y99_SLICE_X93Y99_DO6;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_A = CLBLM_L_X62Y100_SLICE_X92Y100_AO6;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_B = CLBLM_L_X62Y100_SLICE_X92Y100_BO6;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_C = CLBLM_L_X62Y100_SLICE_X92Y100_CO6;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_D = CLBLM_L_X62Y100_SLICE_X92Y100_DO6;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_A = CLBLM_L_X62Y100_SLICE_X93Y100_AO6;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_B = CLBLM_L_X62Y100_SLICE_X93Y100_BO6;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_C = CLBLM_L_X62Y100_SLICE_X93Y100_CO6;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_D = CLBLM_L_X62Y100_SLICE_X93Y100_DO6;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_A = CLBLM_L_X62Y101_SLICE_X92Y101_AO6;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_B = CLBLM_L_X62Y101_SLICE_X92Y101_BO6;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_C = CLBLM_L_X62Y101_SLICE_X92Y101_CO6;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_D = CLBLM_L_X62Y101_SLICE_X92Y101_DO6;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_A = CLBLM_L_X62Y101_SLICE_X93Y101_AO6;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_B = CLBLM_L_X62Y101_SLICE_X93Y101_BO6;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_C = CLBLM_L_X62Y101_SLICE_X93Y101_CO6;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_D = CLBLM_L_X62Y101_SLICE_X93Y101_DO6;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_AMUX = CLBLM_L_X62Y101_SLICE_X93Y101_AO5;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_A = CLBLM_L_X62Y102_SLICE_X92Y102_AO6;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_B = CLBLM_L_X62Y102_SLICE_X92Y102_BO6;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_C = CLBLM_L_X62Y102_SLICE_X92Y102_CO6;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_D = CLBLM_L_X62Y102_SLICE_X92Y102_DO6;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_A = CLBLM_L_X62Y102_SLICE_X93Y102_AO6;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_B = CLBLM_L_X62Y102_SLICE_X93Y102_BO6;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_C = CLBLM_L_X62Y102_SLICE_X93Y102_CO6;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_D = CLBLM_L_X62Y102_SLICE_X93Y102_DO6;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_A = CLBLM_L_X62Y103_SLICE_X92Y103_AO6;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_B = CLBLM_L_X62Y103_SLICE_X92Y103_BO6;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_C = CLBLM_L_X62Y103_SLICE_X92Y103_CO6;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_D = CLBLM_L_X62Y103_SLICE_X92Y103_DO6;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_AMUX = CLBLM_L_X62Y103_SLICE_X92Y103_A5Q;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_BMUX = CLBLM_L_X62Y103_SLICE_X92Y103_B5Q;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_A = CLBLM_L_X62Y103_SLICE_X93Y103_AO6;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_B = CLBLM_L_X62Y103_SLICE_X93Y103_BO6;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_C = CLBLM_L_X62Y103_SLICE_X93Y103_CO6;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_D = CLBLM_L_X62Y103_SLICE_X93Y103_DO6;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_A = CLBLM_L_X62Y105_SLICE_X92Y105_AO6;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_B = CLBLM_L_X62Y105_SLICE_X92Y105_BO6;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_C = CLBLM_L_X62Y105_SLICE_X92Y105_CO6;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_D = CLBLM_L_X62Y105_SLICE_X92Y105_DO6;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_A = CLBLM_L_X62Y105_SLICE_X93Y105_AO6;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_B = CLBLM_L_X62Y105_SLICE_X93Y105_BO6;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_C = CLBLM_L_X62Y105_SLICE_X93Y105_CO6;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_D = CLBLM_L_X62Y105_SLICE_X93Y105_DO6;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_AMUX = CLBLM_L_X62Y105_SLICE_X93Y105_A5Q;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_A = CLBLM_L_X62Y106_SLICE_X92Y106_AO6;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_B = CLBLM_L_X62Y106_SLICE_X92Y106_BO6;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_C = CLBLM_L_X62Y106_SLICE_X92Y106_CO6;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_D = CLBLM_L_X62Y106_SLICE_X92Y106_DO6;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_A = CLBLM_L_X62Y106_SLICE_X93Y106_AO6;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_B = CLBLM_L_X62Y106_SLICE_X93Y106_BO6;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_C = CLBLM_L_X62Y106_SLICE_X93Y106_CO6;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_D = CLBLM_L_X62Y106_SLICE_X93Y106_DO6;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_AMUX = CLBLM_L_X62Y106_SLICE_X93Y106_AO5;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_A = CLBLM_L_X62Y107_SLICE_X92Y107_AO6;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_B = CLBLM_L_X62Y107_SLICE_X92Y107_BO6;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_C = CLBLM_L_X62Y107_SLICE_X92Y107_CO6;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_D = CLBLM_L_X62Y107_SLICE_X92Y107_DO6;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_AMUX = CLBLM_L_X62Y107_SLICE_X92Y107_AO5;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_A = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_B = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_C = CLBLM_L_X62Y107_SLICE_X93Y107_CO6;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_D = CLBLM_L_X62Y107_SLICE_X93Y107_DO6;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_AMUX = CLBLM_L_X62Y107_SLICE_X93Y107_A5Q;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_CMUX = CLBLM_L_X62Y107_SLICE_X93Y107_CO5;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_A = CLBLM_L_X64Y96_SLICE_X96Y96_AO6;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_B = CLBLM_L_X64Y96_SLICE_X96Y96_BO6;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_C = CLBLM_L_X64Y96_SLICE_X96Y96_CO6;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_D = CLBLM_L_X64Y96_SLICE_X96Y96_DO6;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_A = CLBLM_L_X64Y96_SLICE_X97Y96_AO6;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_B = CLBLM_L_X64Y96_SLICE_X97Y96_BO6;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_C = CLBLM_L_X64Y96_SLICE_X97Y96_CO6;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_D = CLBLM_L_X64Y96_SLICE_X97Y96_DO6;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_AMUX = CLBLM_L_X64Y96_SLICE_X97Y96_A5Q;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_A = CLBLM_L_X64Y97_SLICE_X96Y97_AO6;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_B = CLBLM_L_X64Y97_SLICE_X96Y97_BO6;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_C = CLBLM_L_X64Y97_SLICE_X96Y97_CO6;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_D = CLBLM_L_X64Y97_SLICE_X96Y97_DO6;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_A = CLBLM_L_X64Y97_SLICE_X97Y97_AO6;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_B = CLBLM_L_X64Y97_SLICE_X97Y97_BO6;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_C = CLBLM_L_X64Y97_SLICE_X97Y97_CO6;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_D = CLBLM_L_X64Y97_SLICE_X97Y97_DO6;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_AMUX = CLBLM_L_X64Y97_SLICE_X97Y97_A5Q;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_BMUX = CLBLM_L_X64Y97_SLICE_X97Y97_BO5;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_A = CLBLM_L_X64Y98_SLICE_X96Y98_AO6;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_B = CLBLM_L_X64Y98_SLICE_X96Y98_BO6;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_C = CLBLM_L_X64Y98_SLICE_X96Y98_CO6;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_D = CLBLM_L_X64Y98_SLICE_X96Y98_DO6;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_AMUX = CLBLM_L_X64Y98_SLICE_X96Y98_AO5;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_A = CLBLM_L_X64Y98_SLICE_X97Y98_AO6;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_B = CLBLM_L_X64Y98_SLICE_X97Y98_BO6;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_C = CLBLM_L_X64Y98_SLICE_X97Y98_CO6;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_D = CLBLM_L_X64Y98_SLICE_X97Y98_DO6;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_A = CLBLM_L_X64Y99_SLICE_X96Y99_AO6;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_B = CLBLM_L_X64Y99_SLICE_X96Y99_BO6;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_C = CLBLM_L_X64Y99_SLICE_X96Y99_CO6;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_D = CLBLM_L_X64Y99_SLICE_X96Y99_DO6;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_AMUX = CLBLM_L_X64Y99_SLICE_X96Y99_A5Q;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_BMUX = CLBLM_L_X64Y99_SLICE_X96Y99_BO5;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_A = CLBLM_L_X64Y99_SLICE_X97Y99_AO6;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_B = CLBLM_L_X64Y99_SLICE_X97Y99_BO6;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_C = CLBLM_L_X64Y99_SLICE_X97Y99_CO6;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_D = CLBLM_L_X64Y99_SLICE_X97Y99_DO6;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_AMUX = CLBLM_L_X64Y99_SLICE_X97Y99_A5Q;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_BMUX = CLBLM_L_X64Y99_SLICE_X97Y99_B5Q;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_A = CLBLM_L_X64Y100_SLICE_X96Y100_AO6;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_B = CLBLM_L_X64Y100_SLICE_X96Y100_BO6;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_C = CLBLM_L_X64Y100_SLICE_X96Y100_CO6;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_D = CLBLM_L_X64Y100_SLICE_X96Y100_DO6;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_A = CLBLM_L_X64Y100_SLICE_X97Y100_AO6;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_B = CLBLM_L_X64Y100_SLICE_X97Y100_BO6;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_C = CLBLM_L_X64Y100_SLICE_X97Y100_CO6;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_D = CLBLM_L_X64Y100_SLICE_X97Y100_DO6;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_A = CLBLM_L_X64Y101_SLICE_X96Y101_AO6;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_B = CLBLM_L_X64Y101_SLICE_X96Y101_BO6;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_C = CLBLM_L_X64Y101_SLICE_X96Y101_CO6;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_D = CLBLM_L_X64Y101_SLICE_X96Y101_DO6;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_AMUX = CLBLM_L_X64Y101_SLICE_X96Y101_A5Q;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_BMUX = CLBLM_L_X64Y101_SLICE_X96Y101_B5Q;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_CMUX = CLBLM_L_X64Y101_SLICE_X96Y101_C5Q;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_A = CLBLM_L_X64Y101_SLICE_X97Y101_AO6;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_B = CLBLM_L_X64Y101_SLICE_X97Y101_BO6;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_C = CLBLM_L_X64Y101_SLICE_X97Y101_CO6;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_D = CLBLM_L_X64Y101_SLICE_X97Y101_DO6;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_A = CLBLM_L_X64Y102_SLICE_X96Y102_AO6;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_B = CLBLM_L_X64Y102_SLICE_X96Y102_BO6;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_C = CLBLM_L_X64Y102_SLICE_X96Y102_CO6;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_D = CLBLM_L_X64Y102_SLICE_X96Y102_DO6;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_AMUX = CLBLM_L_X64Y102_SLICE_X96Y102_A5Q;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_BMUX = CLBLM_L_X64Y102_SLICE_X96Y102_BO5;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_A = CLBLM_L_X64Y102_SLICE_X97Y102_AO6;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_B = CLBLM_L_X64Y102_SLICE_X97Y102_BO6;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_C = CLBLM_L_X64Y102_SLICE_X97Y102_CO6;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_D = CLBLM_L_X64Y102_SLICE_X97Y102_DO6;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_A = CLBLM_L_X64Y103_SLICE_X96Y103_AO6;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_B = CLBLM_L_X64Y103_SLICE_X96Y103_BO6;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_C = CLBLM_L_X64Y103_SLICE_X96Y103_CO6;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_D = CLBLM_L_X64Y103_SLICE_X96Y103_DO6;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_A = CLBLM_L_X64Y103_SLICE_X97Y103_AO6;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_B = CLBLM_L_X64Y103_SLICE_X97Y103_BO6;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_C = CLBLM_L_X64Y103_SLICE_X97Y103_CO6;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_D = CLBLM_L_X64Y103_SLICE_X97Y103_DO6;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_DMUX = CLBLM_L_X64Y103_SLICE_X97Y103_DO6;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_A = CLBLM_L_X64Y104_SLICE_X96Y104_AO6;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_B = CLBLM_L_X64Y104_SLICE_X96Y104_BO6;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_C = CLBLM_L_X64Y104_SLICE_X96Y104_CO6;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_D = CLBLM_L_X64Y104_SLICE_X96Y104_DO6;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_A = CLBLM_L_X64Y104_SLICE_X97Y104_AO6;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_B = CLBLM_L_X64Y104_SLICE_X97Y104_BO6;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_C = CLBLM_L_X64Y104_SLICE_X97Y104_CO6;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_D = CLBLM_L_X64Y104_SLICE_X97Y104_DO6;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_A = CLBLM_L_X64Y105_SLICE_X96Y105_AO6;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_B = CLBLM_L_X64Y105_SLICE_X96Y105_BO6;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_C = CLBLM_L_X64Y105_SLICE_X96Y105_CO6;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_D = CLBLM_L_X64Y105_SLICE_X96Y105_DO6;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_AMUX = CLBLM_L_X64Y105_SLICE_X96Y105_AO5;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_BMUX = CLBLM_L_X64Y105_SLICE_X96Y105_BO5;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_CMUX = CLBLM_L_X64Y105_SLICE_X96Y105_C5Q;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_A = CLBLM_L_X64Y105_SLICE_X97Y105_AO6;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_B = CLBLM_L_X64Y105_SLICE_X97Y105_BO6;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_C = CLBLM_L_X64Y105_SLICE_X97Y105_CO6;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_D = CLBLM_L_X64Y105_SLICE_X97Y105_DO6;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_A = CLBLM_L_X64Y106_SLICE_X96Y106_AO6;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_B = CLBLM_L_X64Y106_SLICE_X96Y106_BO6;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_C = CLBLM_L_X64Y106_SLICE_X96Y106_CO6;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_D = CLBLM_L_X64Y106_SLICE_X96Y106_DO6;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_AMUX = CLBLM_L_X64Y106_SLICE_X96Y106_A5Q;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_BMUX = CLBLM_L_X64Y106_SLICE_X96Y106_BO5;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_DMUX = CLBLM_L_X64Y106_SLICE_X96Y106_DO5;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_A = CLBLM_L_X64Y106_SLICE_X97Y106_AO6;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_B = CLBLM_L_X64Y106_SLICE_X97Y106_BO6;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_C = CLBLM_L_X64Y106_SLICE_X97Y106_CO6;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_D = CLBLM_L_X64Y106_SLICE_X97Y106_DO6;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_BMUX = CLBLM_L_X64Y106_SLICE_X97Y106_B5Q;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_CMUX = CLBLM_L_X64Y106_SLICE_X97Y106_C5Q;
  assign CLBLM_L_X64Y122_SLICE_X96Y122_A = CLBLM_L_X64Y122_SLICE_X96Y122_AO6;
  assign CLBLM_L_X64Y122_SLICE_X96Y122_B = CLBLM_L_X64Y122_SLICE_X96Y122_BO6;
  assign CLBLM_L_X64Y122_SLICE_X96Y122_C = CLBLM_L_X64Y122_SLICE_X96Y122_CO6;
  assign CLBLM_L_X64Y122_SLICE_X96Y122_D = CLBLM_L_X64Y122_SLICE_X96Y122_DO6;
  assign CLBLM_L_X64Y122_SLICE_X97Y122_A = CLBLM_L_X64Y122_SLICE_X97Y122_AO6;
  assign CLBLM_L_X64Y122_SLICE_X97Y122_B = CLBLM_L_X64Y122_SLICE_X97Y122_BO6;
  assign CLBLM_L_X64Y122_SLICE_X97Y122_C = CLBLM_L_X64Y122_SLICE_X97Y122_CO6;
  assign CLBLM_L_X64Y122_SLICE_X97Y122_D = CLBLM_L_X64Y122_SLICE_X97Y122_DO6;
  assign CLBLM_L_X68Y95_SLICE_X102Y95_A = CLBLM_L_X68Y95_SLICE_X102Y95_AO6;
  assign CLBLM_L_X68Y95_SLICE_X102Y95_B = CLBLM_L_X68Y95_SLICE_X102Y95_BO6;
  assign CLBLM_L_X68Y95_SLICE_X102Y95_C = CLBLM_L_X68Y95_SLICE_X102Y95_CO6;
  assign CLBLM_L_X68Y95_SLICE_X102Y95_D = CLBLM_L_X68Y95_SLICE_X102Y95_DO6;
  assign CLBLM_L_X68Y95_SLICE_X102Y95_AMUX = CLBLM_L_X68Y95_SLICE_X102Y95_A5Q;
  assign CLBLM_L_X68Y95_SLICE_X103Y95_A = CLBLM_L_X68Y95_SLICE_X103Y95_AO6;
  assign CLBLM_L_X68Y95_SLICE_X103Y95_B = CLBLM_L_X68Y95_SLICE_X103Y95_BO6;
  assign CLBLM_L_X68Y95_SLICE_X103Y95_C = CLBLM_L_X68Y95_SLICE_X103Y95_CO6;
  assign CLBLM_L_X68Y95_SLICE_X103Y95_D = CLBLM_L_X68Y95_SLICE_X103Y95_DO6;
  assign CLBLM_L_X68Y96_SLICE_X102Y96_A = CLBLM_L_X68Y96_SLICE_X102Y96_AO6;
  assign CLBLM_L_X68Y96_SLICE_X102Y96_B = CLBLM_L_X68Y96_SLICE_X102Y96_BO6;
  assign CLBLM_L_X68Y96_SLICE_X102Y96_C = CLBLM_L_X68Y96_SLICE_X102Y96_CO6;
  assign CLBLM_L_X68Y96_SLICE_X102Y96_D = CLBLM_L_X68Y96_SLICE_X102Y96_DO6;
  assign CLBLM_L_X68Y96_SLICE_X102Y96_CMUX = CLBLM_L_X68Y96_SLICE_X102Y96_CO6;
  assign CLBLM_L_X68Y96_SLICE_X103Y96_A = CLBLM_L_X68Y96_SLICE_X103Y96_AO6;
  assign CLBLM_L_X68Y96_SLICE_X103Y96_B = CLBLM_L_X68Y96_SLICE_X103Y96_BO6;
  assign CLBLM_L_X68Y96_SLICE_X103Y96_C = CLBLM_L_X68Y96_SLICE_X103Y96_CO6;
  assign CLBLM_L_X68Y96_SLICE_X103Y96_D = CLBLM_L_X68Y96_SLICE_X103Y96_DO6;
  assign CLBLM_L_X68Y96_SLICE_X103Y96_AMUX = CLBLM_L_X68Y96_SLICE_X103Y96_AO6;
  assign CLBLM_L_X68Y97_SLICE_X102Y97_A = CLBLM_L_X68Y97_SLICE_X102Y97_AO6;
  assign CLBLM_L_X68Y97_SLICE_X102Y97_B = CLBLM_L_X68Y97_SLICE_X102Y97_BO6;
  assign CLBLM_L_X68Y97_SLICE_X102Y97_C = CLBLM_L_X68Y97_SLICE_X102Y97_CO6;
  assign CLBLM_L_X68Y97_SLICE_X102Y97_D = CLBLM_L_X68Y97_SLICE_X102Y97_DO6;
  assign CLBLM_L_X68Y97_SLICE_X102Y97_AMUX = CLBLM_L_X68Y97_SLICE_X102Y97_AO5;
  assign CLBLM_L_X68Y97_SLICE_X103Y97_A = CLBLM_L_X68Y97_SLICE_X103Y97_AO6;
  assign CLBLM_L_X68Y97_SLICE_X103Y97_B = CLBLM_L_X68Y97_SLICE_X103Y97_BO6;
  assign CLBLM_L_X68Y97_SLICE_X103Y97_C = CLBLM_L_X68Y97_SLICE_X103Y97_CO6;
  assign CLBLM_L_X68Y97_SLICE_X103Y97_D = CLBLM_L_X68Y97_SLICE_X103Y97_DO6;
  assign CLBLM_L_X68Y98_SLICE_X102Y98_A = CLBLM_L_X68Y98_SLICE_X102Y98_AO6;
  assign CLBLM_L_X68Y98_SLICE_X102Y98_B = CLBLM_L_X68Y98_SLICE_X102Y98_BO6;
  assign CLBLM_L_X68Y98_SLICE_X102Y98_C = CLBLM_L_X68Y98_SLICE_X102Y98_CO6;
  assign CLBLM_L_X68Y98_SLICE_X102Y98_D = CLBLM_L_X68Y98_SLICE_X102Y98_DO6;
  assign CLBLM_L_X68Y98_SLICE_X103Y98_A = CLBLM_L_X68Y98_SLICE_X103Y98_AO6;
  assign CLBLM_L_X68Y98_SLICE_X103Y98_B = CLBLM_L_X68Y98_SLICE_X103Y98_BO6;
  assign CLBLM_L_X68Y98_SLICE_X103Y98_C = CLBLM_L_X68Y98_SLICE_X103Y98_CO6;
  assign CLBLM_L_X68Y98_SLICE_X103Y98_D = CLBLM_L_X68Y98_SLICE_X103Y98_DO6;
  assign CLBLM_L_X68Y98_SLICE_X103Y98_AMUX = CLBLM_L_X68Y98_SLICE_X103Y98_A5Q;
  assign CLBLM_L_X68Y99_SLICE_X102Y99_A = CLBLM_L_X68Y99_SLICE_X102Y99_AO6;
  assign CLBLM_L_X68Y99_SLICE_X102Y99_B = CLBLM_L_X68Y99_SLICE_X102Y99_BO6;
  assign CLBLM_L_X68Y99_SLICE_X102Y99_C = CLBLM_L_X68Y99_SLICE_X102Y99_CO6;
  assign CLBLM_L_X68Y99_SLICE_X102Y99_D = CLBLM_L_X68Y99_SLICE_X102Y99_DO6;
  assign CLBLM_L_X68Y99_SLICE_X102Y99_AMUX = CLBLM_L_X68Y99_SLICE_X102Y99_AO5;
  assign CLBLM_L_X68Y99_SLICE_X102Y99_BMUX = CLBLM_L_X68Y99_SLICE_X102Y99_BO5;
  assign CLBLM_L_X68Y99_SLICE_X102Y99_DMUX = CLBLM_L_X68Y99_SLICE_X102Y99_DO6;
  assign CLBLM_L_X68Y99_SLICE_X103Y99_A = CLBLM_L_X68Y99_SLICE_X103Y99_AO6;
  assign CLBLM_L_X68Y99_SLICE_X103Y99_B = CLBLM_L_X68Y99_SLICE_X103Y99_BO6;
  assign CLBLM_L_X68Y99_SLICE_X103Y99_C = CLBLM_L_X68Y99_SLICE_X103Y99_CO6;
  assign CLBLM_L_X68Y99_SLICE_X103Y99_D = CLBLM_L_X68Y99_SLICE_X103Y99_DO6;
  assign CLBLM_L_X68Y99_SLICE_X103Y99_CMUX = CLBLM_L_X68Y99_SLICE_X103Y99_C5Q;
  assign CLBLM_L_X68Y99_SLICE_X103Y99_DMUX = CLBLM_L_X68Y99_SLICE_X103Y99_D5Q;
  assign CLBLM_L_X68Y100_SLICE_X102Y100_A = CLBLM_L_X68Y100_SLICE_X102Y100_AO6;
  assign CLBLM_L_X68Y100_SLICE_X102Y100_B = CLBLM_L_X68Y100_SLICE_X102Y100_BO6;
  assign CLBLM_L_X68Y100_SLICE_X102Y100_C = CLBLM_L_X68Y100_SLICE_X102Y100_CO6;
  assign CLBLM_L_X68Y100_SLICE_X102Y100_D = CLBLM_L_X68Y100_SLICE_X102Y100_DO6;
  assign CLBLM_L_X68Y100_SLICE_X103Y100_A = CLBLM_L_X68Y100_SLICE_X103Y100_AO6;
  assign CLBLM_L_X68Y100_SLICE_X103Y100_B = CLBLM_L_X68Y100_SLICE_X103Y100_BO6;
  assign CLBLM_L_X68Y100_SLICE_X103Y100_C = CLBLM_L_X68Y100_SLICE_X103Y100_CO6;
  assign CLBLM_L_X68Y100_SLICE_X103Y100_D = CLBLM_L_X68Y100_SLICE_X103Y100_DO6;
  assign CLBLM_L_X68Y101_SLICE_X102Y101_A = CLBLM_L_X68Y101_SLICE_X102Y101_AO6;
  assign CLBLM_L_X68Y101_SLICE_X102Y101_B = CLBLM_L_X68Y101_SLICE_X102Y101_BO6;
  assign CLBLM_L_X68Y101_SLICE_X102Y101_C = CLBLM_L_X68Y101_SLICE_X102Y101_CO6;
  assign CLBLM_L_X68Y101_SLICE_X102Y101_D = CLBLM_L_X68Y101_SLICE_X102Y101_DO6;
  assign CLBLM_L_X68Y101_SLICE_X102Y101_AMUX = CLBLM_L_X68Y101_SLICE_X102Y101_A5Q;
  assign CLBLM_L_X68Y101_SLICE_X102Y101_BMUX = CLBLM_L_X68Y101_SLICE_X102Y101_BO5;
  assign CLBLM_L_X68Y101_SLICE_X103Y101_A = CLBLM_L_X68Y101_SLICE_X103Y101_AO6;
  assign CLBLM_L_X68Y101_SLICE_X103Y101_B = CLBLM_L_X68Y101_SLICE_X103Y101_BO6;
  assign CLBLM_L_X68Y101_SLICE_X103Y101_C = CLBLM_L_X68Y101_SLICE_X103Y101_CO6;
  assign CLBLM_L_X68Y101_SLICE_X103Y101_D = CLBLM_L_X68Y101_SLICE_X103Y101_DO6;
  assign CLBLM_L_X68Y102_SLICE_X102Y102_A = CLBLM_L_X68Y102_SLICE_X102Y102_AO6;
  assign CLBLM_L_X68Y102_SLICE_X102Y102_B = CLBLM_L_X68Y102_SLICE_X102Y102_BO6;
  assign CLBLM_L_X68Y102_SLICE_X102Y102_C = CLBLM_L_X68Y102_SLICE_X102Y102_CO6;
  assign CLBLM_L_X68Y102_SLICE_X102Y102_D = CLBLM_L_X68Y102_SLICE_X102Y102_DO6;
  assign CLBLM_L_X68Y102_SLICE_X103Y102_A = CLBLM_L_X68Y102_SLICE_X103Y102_AO6;
  assign CLBLM_L_X68Y102_SLICE_X103Y102_B = CLBLM_L_X68Y102_SLICE_X103Y102_BO6;
  assign CLBLM_L_X68Y102_SLICE_X103Y102_C = CLBLM_L_X68Y102_SLICE_X103Y102_CO6;
  assign CLBLM_L_X68Y102_SLICE_X103Y102_D = CLBLM_L_X68Y102_SLICE_X103Y102_DO6;
  assign CLBLM_L_X68Y103_SLICE_X102Y103_A = CLBLM_L_X68Y103_SLICE_X102Y103_AO6;
  assign CLBLM_L_X68Y103_SLICE_X102Y103_B = CLBLM_L_X68Y103_SLICE_X102Y103_BO6;
  assign CLBLM_L_X68Y103_SLICE_X102Y103_C = CLBLM_L_X68Y103_SLICE_X102Y103_CO6;
  assign CLBLM_L_X68Y103_SLICE_X102Y103_D = CLBLM_L_X68Y103_SLICE_X102Y103_DO6;
  assign CLBLM_L_X68Y103_SLICE_X102Y103_BMUX = CLBLM_L_X68Y103_SLICE_X102Y103_B5Q;
  assign CLBLM_L_X68Y103_SLICE_X103Y103_A = CLBLM_L_X68Y103_SLICE_X103Y103_AO6;
  assign CLBLM_L_X68Y103_SLICE_X103Y103_B = CLBLM_L_X68Y103_SLICE_X103Y103_BO6;
  assign CLBLM_L_X68Y103_SLICE_X103Y103_C = CLBLM_L_X68Y103_SLICE_X103Y103_CO6;
  assign CLBLM_L_X68Y103_SLICE_X103Y103_D = CLBLM_L_X68Y103_SLICE_X103Y103_DO6;
  assign CLBLM_L_X68Y105_SLICE_X102Y105_A = CLBLM_L_X68Y105_SLICE_X102Y105_AO6;
  assign CLBLM_L_X68Y105_SLICE_X102Y105_B = CLBLM_L_X68Y105_SLICE_X102Y105_BO6;
  assign CLBLM_L_X68Y105_SLICE_X102Y105_C = CLBLM_L_X68Y105_SLICE_X102Y105_CO6;
  assign CLBLM_L_X68Y105_SLICE_X102Y105_D = CLBLM_L_X68Y105_SLICE_X102Y105_DO6;
  assign CLBLM_L_X68Y105_SLICE_X102Y105_AMUX = CLBLM_L_X68Y105_SLICE_X102Y105_AO5;
  assign CLBLM_L_X68Y105_SLICE_X103Y105_A = CLBLM_L_X68Y105_SLICE_X103Y105_AO6;
  assign CLBLM_L_X68Y105_SLICE_X103Y105_B = CLBLM_L_X68Y105_SLICE_X103Y105_BO6;
  assign CLBLM_L_X68Y105_SLICE_X103Y105_C = CLBLM_L_X68Y105_SLICE_X103Y105_CO6;
  assign CLBLM_L_X68Y105_SLICE_X103Y105_D = CLBLM_L_X68Y105_SLICE_X103Y105_DO6;
  assign CLBLM_L_X68Y106_SLICE_X102Y106_A = CLBLM_L_X68Y106_SLICE_X102Y106_AO6;
  assign CLBLM_L_X68Y106_SLICE_X102Y106_B = CLBLM_L_X68Y106_SLICE_X102Y106_BO6;
  assign CLBLM_L_X68Y106_SLICE_X102Y106_C = CLBLM_L_X68Y106_SLICE_X102Y106_CO6;
  assign CLBLM_L_X68Y106_SLICE_X102Y106_D = CLBLM_L_X68Y106_SLICE_X102Y106_DO6;
  assign CLBLM_L_X68Y106_SLICE_X102Y106_AMUX = CLBLM_L_X68Y106_SLICE_X102Y106_AO5;
  assign CLBLM_L_X68Y106_SLICE_X103Y106_A = CLBLM_L_X68Y106_SLICE_X103Y106_AO6;
  assign CLBLM_L_X68Y106_SLICE_X103Y106_B = CLBLM_L_X68Y106_SLICE_X103Y106_BO6;
  assign CLBLM_L_X68Y106_SLICE_X103Y106_C = CLBLM_L_X68Y106_SLICE_X103Y106_CO6;
  assign CLBLM_L_X68Y106_SLICE_X103Y106_D = CLBLM_L_X68Y106_SLICE_X103Y106_DO6;
  assign CLBLM_L_X68Y106_SLICE_X103Y106_AMUX = CLBLM_L_X68Y106_SLICE_X103Y106_AO5;
  assign CLBLM_L_X68Y106_SLICE_X103Y106_BMUX = CLBLM_L_X68Y106_SLICE_X103Y106_B5Q;
  assign CLBLM_L_X68Y107_SLICE_X102Y107_A = CLBLM_L_X68Y107_SLICE_X102Y107_AO6;
  assign CLBLM_L_X68Y107_SLICE_X102Y107_B = CLBLM_L_X68Y107_SLICE_X102Y107_BO6;
  assign CLBLM_L_X68Y107_SLICE_X102Y107_C = CLBLM_L_X68Y107_SLICE_X102Y107_CO6;
  assign CLBLM_L_X68Y107_SLICE_X102Y107_D = CLBLM_L_X68Y107_SLICE_X102Y107_DO6;
  assign CLBLM_L_X68Y107_SLICE_X102Y107_AMUX = CLBLM_L_X68Y107_SLICE_X102Y107_AO5;
  assign CLBLM_L_X68Y107_SLICE_X103Y107_A = CLBLM_L_X68Y107_SLICE_X103Y107_AO6;
  assign CLBLM_L_X68Y107_SLICE_X103Y107_B = CLBLM_L_X68Y107_SLICE_X103Y107_BO6;
  assign CLBLM_L_X68Y107_SLICE_X103Y107_C = CLBLM_L_X68Y107_SLICE_X103Y107_CO6;
  assign CLBLM_L_X68Y107_SLICE_X103Y107_D = CLBLM_L_X68Y107_SLICE_X103Y107_DO6;
  assign CLBLM_L_X68Y107_SLICE_X103Y107_CMUX = CLBLM_L_X68Y107_SLICE_X103Y107_CO6;
  assign CLBLM_L_X68Y108_SLICE_X102Y108_A = CLBLM_L_X68Y108_SLICE_X102Y108_AO6;
  assign CLBLM_L_X68Y108_SLICE_X102Y108_B = CLBLM_L_X68Y108_SLICE_X102Y108_BO6;
  assign CLBLM_L_X68Y108_SLICE_X102Y108_C = CLBLM_L_X68Y108_SLICE_X102Y108_CO6;
  assign CLBLM_L_X68Y108_SLICE_X102Y108_D = CLBLM_L_X68Y108_SLICE_X102Y108_DO6;
  assign CLBLM_L_X68Y108_SLICE_X102Y108_AMUX = CLBLM_L_X68Y108_SLICE_X102Y108_A5Q;
  assign CLBLM_L_X68Y108_SLICE_X102Y108_BMUX = CLBLM_L_X68Y108_SLICE_X102Y108_B5Q;
  assign CLBLM_L_X68Y108_SLICE_X102Y108_CMUX = CLBLM_L_X68Y108_SLICE_X102Y108_CO6;
  assign CLBLM_L_X68Y108_SLICE_X103Y108_A = CLBLM_L_X68Y108_SLICE_X103Y108_AO6;
  assign CLBLM_L_X68Y108_SLICE_X103Y108_B = CLBLM_L_X68Y108_SLICE_X103Y108_BO6;
  assign CLBLM_L_X68Y108_SLICE_X103Y108_C = CLBLM_L_X68Y108_SLICE_X103Y108_CO6;
  assign CLBLM_L_X68Y108_SLICE_X103Y108_D = CLBLM_L_X68Y108_SLICE_X103Y108_DO6;
  assign CLBLM_L_X68Y108_SLICE_X103Y108_AMUX = CLBLM_L_X68Y108_SLICE_X103Y108_A5Q;
  assign CLBLM_L_X68Y109_SLICE_X102Y109_A = CLBLM_L_X68Y109_SLICE_X102Y109_AO6;
  assign CLBLM_L_X68Y109_SLICE_X102Y109_B = CLBLM_L_X68Y109_SLICE_X102Y109_BO6;
  assign CLBLM_L_X68Y109_SLICE_X102Y109_C = CLBLM_L_X68Y109_SLICE_X102Y109_CO6;
  assign CLBLM_L_X68Y109_SLICE_X102Y109_D = CLBLM_L_X68Y109_SLICE_X102Y109_DO6;
  assign CLBLM_L_X68Y109_SLICE_X102Y109_AMUX = CLBLM_L_X68Y109_SLICE_X102Y109_A5Q;
  assign CLBLM_L_X68Y109_SLICE_X102Y109_BMUX = CLBLM_L_X68Y109_SLICE_X102Y109_BO5;
  assign CLBLM_L_X68Y109_SLICE_X102Y109_CMUX = CLBLM_L_X68Y109_SLICE_X102Y109_CO6;
  assign CLBLM_L_X68Y109_SLICE_X103Y109_A = CLBLM_L_X68Y109_SLICE_X103Y109_AO6;
  assign CLBLM_L_X68Y109_SLICE_X103Y109_B = CLBLM_L_X68Y109_SLICE_X103Y109_BO6;
  assign CLBLM_L_X68Y109_SLICE_X103Y109_C = CLBLM_L_X68Y109_SLICE_X103Y109_CO6;
  assign CLBLM_L_X68Y109_SLICE_X103Y109_D = CLBLM_L_X68Y109_SLICE_X103Y109_DO6;
  assign CLBLM_L_X68Y109_SLICE_X103Y109_BMUX = CLBLM_L_X68Y109_SLICE_X103Y109_B5Q;
  assign CLBLM_L_X68Y112_SLICE_X102Y112_A = CLBLM_L_X68Y112_SLICE_X102Y112_AO6;
  assign CLBLM_L_X68Y112_SLICE_X102Y112_B = CLBLM_L_X68Y112_SLICE_X102Y112_BO6;
  assign CLBLM_L_X68Y112_SLICE_X102Y112_C = CLBLM_L_X68Y112_SLICE_X102Y112_CO6;
  assign CLBLM_L_X68Y112_SLICE_X102Y112_D = CLBLM_L_X68Y112_SLICE_X102Y112_DO6;
  assign CLBLM_L_X68Y112_SLICE_X103Y112_A = CLBLM_L_X68Y112_SLICE_X103Y112_AO6;
  assign CLBLM_L_X68Y112_SLICE_X103Y112_B = CLBLM_L_X68Y112_SLICE_X103Y112_BO6;
  assign CLBLM_L_X68Y112_SLICE_X103Y112_C = CLBLM_L_X68Y112_SLICE_X103Y112_CO6;
  assign CLBLM_L_X68Y112_SLICE_X103Y112_D = CLBLM_L_X68Y112_SLICE_X103Y112_DO6;
  assign CLBLM_L_X68Y121_SLICE_X102Y121_A = CLBLM_L_X68Y121_SLICE_X102Y121_AO6;
  assign CLBLM_L_X68Y121_SLICE_X102Y121_B = CLBLM_L_X68Y121_SLICE_X102Y121_BO6;
  assign CLBLM_L_X68Y121_SLICE_X102Y121_C = CLBLM_L_X68Y121_SLICE_X102Y121_CO6;
  assign CLBLM_L_X68Y121_SLICE_X102Y121_D = CLBLM_L_X68Y121_SLICE_X102Y121_DO6;
  assign CLBLM_L_X68Y121_SLICE_X103Y121_A = CLBLM_L_X68Y121_SLICE_X103Y121_AO6;
  assign CLBLM_L_X68Y121_SLICE_X103Y121_B = CLBLM_L_X68Y121_SLICE_X103Y121_BO6;
  assign CLBLM_L_X68Y121_SLICE_X103Y121_C = CLBLM_L_X68Y121_SLICE_X103Y121_CO6;
  assign CLBLM_L_X68Y121_SLICE_X103Y121_D = CLBLM_L_X68Y121_SLICE_X103Y121_DO6;
  assign CLBLM_L_X70Y98_SLICE_X104Y98_A = CLBLM_L_X70Y98_SLICE_X104Y98_AO6;
  assign CLBLM_L_X70Y98_SLICE_X104Y98_B = CLBLM_L_X70Y98_SLICE_X104Y98_BO6;
  assign CLBLM_L_X70Y98_SLICE_X104Y98_C = CLBLM_L_X70Y98_SLICE_X104Y98_CO6;
  assign CLBLM_L_X70Y98_SLICE_X104Y98_D = CLBLM_L_X70Y98_SLICE_X104Y98_DO6;
  assign CLBLM_L_X70Y98_SLICE_X105Y98_A = CLBLM_L_X70Y98_SLICE_X105Y98_AO6;
  assign CLBLM_L_X70Y98_SLICE_X105Y98_B = CLBLM_L_X70Y98_SLICE_X105Y98_BO6;
  assign CLBLM_L_X70Y98_SLICE_X105Y98_C = CLBLM_L_X70Y98_SLICE_X105Y98_CO6;
  assign CLBLM_L_X70Y98_SLICE_X105Y98_D = CLBLM_L_X70Y98_SLICE_X105Y98_DO6;
  assign CLBLM_L_X70Y99_SLICE_X104Y99_A = CLBLM_L_X70Y99_SLICE_X104Y99_AO6;
  assign CLBLM_L_X70Y99_SLICE_X104Y99_B = CLBLM_L_X70Y99_SLICE_X104Y99_BO6;
  assign CLBLM_L_X70Y99_SLICE_X104Y99_C = CLBLM_L_X70Y99_SLICE_X104Y99_CO6;
  assign CLBLM_L_X70Y99_SLICE_X104Y99_D = CLBLM_L_X70Y99_SLICE_X104Y99_DO6;
  assign CLBLM_L_X70Y99_SLICE_X105Y99_A = CLBLM_L_X70Y99_SLICE_X105Y99_AO6;
  assign CLBLM_L_X70Y99_SLICE_X105Y99_B = CLBLM_L_X70Y99_SLICE_X105Y99_BO6;
  assign CLBLM_L_X70Y99_SLICE_X105Y99_C = CLBLM_L_X70Y99_SLICE_X105Y99_CO6;
  assign CLBLM_L_X70Y99_SLICE_X105Y99_D = CLBLM_L_X70Y99_SLICE_X105Y99_DO6;
  assign CLBLM_L_X70Y99_SLICE_X105Y99_AMUX = CLBLM_L_X70Y99_SLICE_X105Y99_AO5;
  assign CLBLM_L_X70Y100_SLICE_X104Y100_A = CLBLM_L_X70Y100_SLICE_X104Y100_AO6;
  assign CLBLM_L_X70Y100_SLICE_X104Y100_B = CLBLM_L_X70Y100_SLICE_X104Y100_BO6;
  assign CLBLM_L_X70Y100_SLICE_X104Y100_C = CLBLM_L_X70Y100_SLICE_X104Y100_CO6;
  assign CLBLM_L_X70Y100_SLICE_X104Y100_D = CLBLM_L_X70Y100_SLICE_X104Y100_DO6;
  assign CLBLM_L_X70Y100_SLICE_X104Y100_AMUX = CLBLM_L_X70Y100_SLICE_X104Y100_A5Q;
  assign CLBLM_L_X70Y100_SLICE_X105Y100_A = CLBLM_L_X70Y100_SLICE_X105Y100_AO6;
  assign CLBLM_L_X70Y100_SLICE_X105Y100_B = CLBLM_L_X70Y100_SLICE_X105Y100_BO6;
  assign CLBLM_L_X70Y100_SLICE_X105Y100_C = CLBLM_L_X70Y100_SLICE_X105Y100_CO6;
  assign CLBLM_L_X70Y100_SLICE_X105Y100_D = CLBLM_L_X70Y100_SLICE_X105Y100_DO6;
  assign CLBLM_L_X70Y100_SLICE_X105Y100_AMUX = CLBLM_L_X70Y100_SLICE_X105Y100_A5Q;
  assign CLBLM_L_X70Y100_SLICE_X105Y100_BMUX = CLBLM_L_X70Y100_SLICE_X105Y100_B5Q;
  assign CLBLM_L_X70Y101_SLICE_X104Y101_A = CLBLM_L_X70Y101_SLICE_X104Y101_AO6;
  assign CLBLM_L_X70Y101_SLICE_X104Y101_B = CLBLM_L_X70Y101_SLICE_X104Y101_BO6;
  assign CLBLM_L_X70Y101_SLICE_X104Y101_C = CLBLM_L_X70Y101_SLICE_X104Y101_CO6;
  assign CLBLM_L_X70Y101_SLICE_X104Y101_D = CLBLM_L_X70Y101_SLICE_X104Y101_DO6;
  assign CLBLM_L_X70Y101_SLICE_X104Y101_AMUX = CLBLM_L_X70Y101_SLICE_X104Y101_AO5;
  assign CLBLM_L_X70Y101_SLICE_X105Y101_A = CLBLM_L_X70Y101_SLICE_X105Y101_AO6;
  assign CLBLM_L_X70Y101_SLICE_X105Y101_B = CLBLM_L_X70Y101_SLICE_X105Y101_BO6;
  assign CLBLM_L_X70Y101_SLICE_X105Y101_C = CLBLM_L_X70Y101_SLICE_X105Y101_CO6;
  assign CLBLM_L_X70Y101_SLICE_X105Y101_D = CLBLM_L_X70Y101_SLICE_X105Y101_DO6;
  assign CLBLM_L_X70Y101_SLICE_X105Y101_AMUX = CLBLM_L_X70Y101_SLICE_X105Y101_AO5;
  assign CLBLM_L_X70Y102_SLICE_X104Y102_A = CLBLM_L_X70Y102_SLICE_X104Y102_AO6;
  assign CLBLM_L_X70Y102_SLICE_X104Y102_B = CLBLM_L_X70Y102_SLICE_X104Y102_BO6;
  assign CLBLM_L_X70Y102_SLICE_X104Y102_C = CLBLM_L_X70Y102_SLICE_X104Y102_CO6;
  assign CLBLM_L_X70Y102_SLICE_X104Y102_D = CLBLM_L_X70Y102_SLICE_X104Y102_DO6;
  assign CLBLM_L_X70Y102_SLICE_X105Y102_A = CLBLM_L_X70Y102_SLICE_X105Y102_AO6;
  assign CLBLM_L_X70Y102_SLICE_X105Y102_B = CLBLM_L_X70Y102_SLICE_X105Y102_BO6;
  assign CLBLM_L_X70Y102_SLICE_X105Y102_C = CLBLM_L_X70Y102_SLICE_X105Y102_CO6;
  assign CLBLM_L_X70Y102_SLICE_X105Y102_D = CLBLM_L_X70Y102_SLICE_X105Y102_DO6;
  assign CLBLM_L_X70Y103_SLICE_X104Y103_A = CLBLM_L_X70Y103_SLICE_X104Y103_AO6;
  assign CLBLM_L_X70Y103_SLICE_X104Y103_B = CLBLM_L_X70Y103_SLICE_X104Y103_BO6;
  assign CLBLM_L_X70Y103_SLICE_X104Y103_C = CLBLM_L_X70Y103_SLICE_X104Y103_CO6;
  assign CLBLM_L_X70Y103_SLICE_X104Y103_D = CLBLM_L_X70Y103_SLICE_X104Y103_DO6;
  assign CLBLM_L_X70Y103_SLICE_X104Y103_BMUX = CLBLM_L_X70Y103_SLICE_X104Y103_B5Q;
  assign CLBLM_L_X70Y103_SLICE_X104Y103_CMUX = CLBLM_L_X70Y103_SLICE_X104Y103_C5Q;
  assign CLBLM_L_X70Y103_SLICE_X104Y103_DMUX = CLBLM_L_X70Y103_SLICE_X104Y103_DO5;
  assign CLBLM_L_X70Y103_SLICE_X105Y103_A = CLBLM_L_X70Y103_SLICE_X105Y103_AO6;
  assign CLBLM_L_X70Y103_SLICE_X105Y103_B = CLBLM_L_X70Y103_SLICE_X105Y103_BO6;
  assign CLBLM_L_X70Y103_SLICE_X105Y103_C = CLBLM_L_X70Y103_SLICE_X105Y103_CO6;
  assign CLBLM_L_X70Y103_SLICE_X105Y103_D = CLBLM_L_X70Y103_SLICE_X105Y103_DO6;
  assign CLBLM_L_X70Y103_SLICE_X105Y103_CMUX = CLBLM_L_X70Y103_SLICE_X105Y103_CO5;
  assign CLBLM_L_X70Y103_SLICE_X105Y103_DMUX = CLBLM_L_X70Y103_SLICE_X105Y103_DO5;
  assign CLBLM_L_X70Y104_SLICE_X104Y104_A = CLBLM_L_X70Y104_SLICE_X104Y104_AO6;
  assign CLBLM_L_X70Y104_SLICE_X104Y104_B = CLBLM_L_X70Y104_SLICE_X104Y104_BO6;
  assign CLBLM_L_X70Y104_SLICE_X104Y104_C = CLBLM_L_X70Y104_SLICE_X104Y104_CO6;
  assign CLBLM_L_X70Y104_SLICE_X104Y104_D = CLBLM_L_X70Y104_SLICE_X104Y104_DO6;
  assign CLBLM_L_X70Y104_SLICE_X104Y104_AMUX = CLBLM_L_X70Y104_SLICE_X104Y104_A5Q;
  assign CLBLM_L_X70Y104_SLICE_X104Y104_CMUX = CLBLM_L_X70Y104_SLICE_X104Y104_CO5;
  assign CLBLM_L_X70Y104_SLICE_X105Y104_A = CLBLM_L_X70Y104_SLICE_X105Y104_AO6;
  assign CLBLM_L_X70Y104_SLICE_X105Y104_B = CLBLM_L_X70Y104_SLICE_X105Y104_BO6;
  assign CLBLM_L_X70Y104_SLICE_X105Y104_C = CLBLM_L_X70Y104_SLICE_X105Y104_CO6;
  assign CLBLM_L_X70Y104_SLICE_X105Y104_D = CLBLM_L_X70Y104_SLICE_X105Y104_DO6;
  assign CLBLM_L_X70Y104_SLICE_X105Y104_DMUX = CLBLM_L_X70Y104_SLICE_X105Y104_D5Q;
  assign CLBLM_L_X70Y105_SLICE_X104Y105_A = CLBLM_L_X70Y105_SLICE_X104Y105_AO6;
  assign CLBLM_L_X70Y105_SLICE_X104Y105_B = CLBLM_L_X70Y105_SLICE_X104Y105_BO6;
  assign CLBLM_L_X70Y105_SLICE_X104Y105_C = CLBLM_L_X70Y105_SLICE_X104Y105_CO6;
  assign CLBLM_L_X70Y105_SLICE_X104Y105_D = CLBLM_L_X70Y105_SLICE_X104Y105_DO6;
  assign CLBLM_L_X70Y105_SLICE_X105Y105_A = CLBLM_L_X70Y105_SLICE_X105Y105_AO6;
  assign CLBLM_L_X70Y105_SLICE_X105Y105_B = CLBLM_L_X70Y105_SLICE_X105Y105_BO6;
  assign CLBLM_L_X70Y105_SLICE_X105Y105_C = CLBLM_L_X70Y105_SLICE_X105Y105_CO6;
  assign CLBLM_L_X70Y105_SLICE_X105Y105_D = CLBLM_L_X70Y105_SLICE_X105Y105_DO6;
  assign CLBLM_L_X70Y105_SLICE_X105Y105_AMUX = CLBLM_L_X70Y105_SLICE_X105Y105_A5Q;
  assign CLBLM_L_X70Y106_SLICE_X104Y106_A = CLBLM_L_X70Y106_SLICE_X104Y106_AO6;
  assign CLBLM_L_X70Y106_SLICE_X104Y106_B = CLBLM_L_X70Y106_SLICE_X104Y106_BO6;
  assign CLBLM_L_X70Y106_SLICE_X104Y106_C = CLBLM_L_X70Y106_SLICE_X104Y106_CO6;
  assign CLBLM_L_X70Y106_SLICE_X104Y106_D = CLBLM_L_X70Y106_SLICE_X104Y106_DO6;
  assign CLBLM_L_X70Y106_SLICE_X104Y106_AMUX = CLBLM_L_X70Y106_SLICE_X104Y106_A5Q;
  assign CLBLM_L_X70Y106_SLICE_X105Y106_A = CLBLM_L_X70Y106_SLICE_X105Y106_AO6;
  assign CLBLM_L_X70Y106_SLICE_X105Y106_B = CLBLM_L_X70Y106_SLICE_X105Y106_BO6;
  assign CLBLM_L_X70Y106_SLICE_X105Y106_C = CLBLM_L_X70Y106_SLICE_X105Y106_CO6;
  assign CLBLM_L_X70Y106_SLICE_X105Y106_D = CLBLM_L_X70Y106_SLICE_X105Y106_DO6;
  assign CLBLM_L_X70Y106_SLICE_X105Y106_AMUX = CLBLM_L_X70Y106_SLICE_X105Y106_A5Q;
  assign CLBLM_L_X70Y107_SLICE_X104Y107_A = CLBLM_L_X70Y107_SLICE_X104Y107_AO6;
  assign CLBLM_L_X70Y107_SLICE_X104Y107_B = CLBLM_L_X70Y107_SLICE_X104Y107_BO6;
  assign CLBLM_L_X70Y107_SLICE_X104Y107_C = CLBLM_L_X70Y107_SLICE_X104Y107_CO6;
  assign CLBLM_L_X70Y107_SLICE_X104Y107_D = CLBLM_L_X70Y107_SLICE_X104Y107_DO6;
  assign CLBLM_L_X70Y107_SLICE_X105Y107_A = CLBLM_L_X70Y107_SLICE_X105Y107_AO6;
  assign CLBLM_L_X70Y107_SLICE_X105Y107_B = CLBLM_L_X70Y107_SLICE_X105Y107_BO6;
  assign CLBLM_L_X70Y107_SLICE_X105Y107_C = CLBLM_L_X70Y107_SLICE_X105Y107_CO6;
  assign CLBLM_L_X70Y107_SLICE_X105Y107_D = CLBLM_L_X70Y107_SLICE_X105Y107_DO6;
  assign CLBLM_L_X70Y108_SLICE_X104Y108_A = CLBLM_L_X70Y108_SLICE_X104Y108_AO6;
  assign CLBLM_L_X70Y108_SLICE_X104Y108_B = CLBLM_L_X70Y108_SLICE_X104Y108_BO6;
  assign CLBLM_L_X70Y108_SLICE_X104Y108_C = CLBLM_L_X70Y108_SLICE_X104Y108_CO6;
  assign CLBLM_L_X70Y108_SLICE_X104Y108_D = CLBLM_L_X70Y108_SLICE_X104Y108_DO6;
  assign CLBLM_L_X70Y108_SLICE_X105Y108_A = CLBLM_L_X70Y108_SLICE_X105Y108_AO6;
  assign CLBLM_L_X70Y108_SLICE_X105Y108_B = CLBLM_L_X70Y108_SLICE_X105Y108_BO6;
  assign CLBLM_L_X70Y108_SLICE_X105Y108_C = CLBLM_L_X70Y108_SLICE_X105Y108_CO6;
  assign CLBLM_L_X70Y108_SLICE_X105Y108_D = CLBLM_L_X70Y108_SLICE_X105Y108_DO6;
  assign CLBLM_L_X70Y108_SLICE_X105Y108_AMUX = CLBLM_L_X70Y108_SLICE_X105Y108_AO5;
  assign CLBLM_L_X70Y109_SLICE_X104Y109_A = CLBLM_L_X70Y109_SLICE_X104Y109_AO6;
  assign CLBLM_L_X70Y109_SLICE_X104Y109_B = CLBLM_L_X70Y109_SLICE_X104Y109_BO6;
  assign CLBLM_L_X70Y109_SLICE_X104Y109_C = CLBLM_L_X70Y109_SLICE_X104Y109_CO6;
  assign CLBLM_L_X70Y109_SLICE_X104Y109_D = CLBLM_L_X70Y109_SLICE_X104Y109_DO6;
  assign CLBLM_L_X70Y109_SLICE_X104Y109_AMUX = CLBLM_L_X70Y109_SLICE_X104Y109_A5Q;
  assign CLBLM_L_X70Y109_SLICE_X104Y109_BMUX = CLBLM_L_X70Y109_SLICE_X104Y109_B5Q;
  assign CLBLM_L_X70Y109_SLICE_X105Y109_A = CLBLM_L_X70Y109_SLICE_X105Y109_AO6;
  assign CLBLM_L_X70Y109_SLICE_X105Y109_B = CLBLM_L_X70Y109_SLICE_X105Y109_BO6;
  assign CLBLM_L_X70Y109_SLICE_X105Y109_C = CLBLM_L_X70Y109_SLICE_X105Y109_CO6;
  assign CLBLM_L_X70Y109_SLICE_X105Y109_D = CLBLM_L_X70Y109_SLICE_X105Y109_DO6;
  assign CLBLM_L_X70Y110_SLICE_X104Y110_A = CLBLM_L_X70Y110_SLICE_X104Y110_AO6;
  assign CLBLM_L_X70Y110_SLICE_X104Y110_B = CLBLM_L_X70Y110_SLICE_X104Y110_BO6;
  assign CLBLM_L_X70Y110_SLICE_X104Y110_C = CLBLM_L_X70Y110_SLICE_X104Y110_CO6;
  assign CLBLM_L_X70Y110_SLICE_X104Y110_D = CLBLM_L_X70Y110_SLICE_X104Y110_DO6;
  assign CLBLM_L_X70Y110_SLICE_X104Y110_AMUX = CLBLM_L_X70Y110_SLICE_X104Y110_AO5;
  assign CLBLM_L_X70Y110_SLICE_X104Y110_BMUX = CLBLM_L_X70Y110_SLICE_X104Y110_B5Q;
  assign CLBLM_L_X70Y110_SLICE_X105Y110_A = CLBLM_L_X70Y110_SLICE_X105Y110_AO6;
  assign CLBLM_L_X70Y110_SLICE_X105Y110_B = CLBLM_L_X70Y110_SLICE_X105Y110_BO6;
  assign CLBLM_L_X70Y110_SLICE_X105Y110_C = CLBLM_L_X70Y110_SLICE_X105Y110_CO6;
  assign CLBLM_L_X70Y110_SLICE_X105Y110_D = CLBLM_L_X70Y110_SLICE_X105Y110_DO6;
  assign CLBLM_L_X70Y111_SLICE_X104Y111_A = CLBLM_L_X70Y111_SLICE_X104Y111_AO6;
  assign CLBLM_L_X70Y111_SLICE_X104Y111_B = CLBLM_L_X70Y111_SLICE_X104Y111_BO6;
  assign CLBLM_L_X70Y111_SLICE_X104Y111_C = CLBLM_L_X70Y111_SLICE_X104Y111_CO6;
  assign CLBLM_L_X70Y111_SLICE_X104Y111_D = CLBLM_L_X70Y111_SLICE_X104Y111_DO6;
  assign CLBLM_L_X70Y111_SLICE_X104Y111_AMUX = CLBLM_L_X70Y111_SLICE_X104Y111_AO5;
  assign CLBLM_L_X70Y111_SLICE_X104Y111_BMUX = CLBLM_L_X70Y111_SLICE_X104Y111_BO5;
  assign CLBLM_L_X70Y111_SLICE_X104Y111_CMUX = CLBLM_L_X70Y111_SLICE_X104Y111_CO6;
  assign CLBLM_L_X70Y111_SLICE_X105Y111_A = CLBLM_L_X70Y111_SLICE_X105Y111_AO6;
  assign CLBLM_L_X70Y111_SLICE_X105Y111_B = CLBLM_L_X70Y111_SLICE_X105Y111_BO6;
  assign CLBLM_L_X70Y111_SLICE_X105Y111_C = CLBLM_L_X70Y111_SLICE_X105Y111_CO6;
  assign CLBLM_L_X70Y111_SLICE_X105Y111_D = CLBLM_L_X70Y111_SLICE_X105Y111_DO6;
  assign CLBLM_L_X70Y112_SLICE_X104Y112_A = CLBLM_L_X70Y112_SLICE_X104Y112_AO6;
  assign CLBLM_L_X70Y112_SLICE_X104Y112_B = CLBLM_L_X70Y112_SLICE_X104Y112_BO6;
  assign CLBLM_L_X70Y112_SLICE_X104Y112_C = CLBLM_L_X70Y112_SLICE_X104Y112_CO6;
  assign CLBLM_L_X70Y112_SLICE_X104Y112_D = CLBLM_L_X70Y112_SLICE_X104Y112_DO6;
  assign CLBLM_L_X70Y112_SLICE_X104Y112_AMUX = CLBLM_L_X70Y112_SLICE_X104Y112_A5Q;
  assign CLBLM_L_X70Y112_SLICE_X104Y112_BMUX = CLBLM_L_X70Y112_SLICE_X104Y112_BO5;
  assign CLBLM_L_X70Y112_SLICE_X104Y112_CMUX = CLBLM_L_X70Y112_SLICE_X104Y112_C5Q;
  assign CLBLM_L_X70Y112_SLICE_X105Y112_A = CLBLM_L_X70Y112_SLICE_X105Y112_AO6;
  assign CLBLM_L_X70Y112_SLICE_X105Y112_B = CLBLM_L_X70Y112_SLICE_X105Y112_BO6;
  assign CLBLM_L_X70Y112_SLICE_X105Y112_C = CLBLM_L_X70Y112_SLICE_X105Y112_CO6;
  assign CLBLM_L_X70Y112_SLICE_X105Y112_D = CLBLM_L_X70Y112_SLICE_X105Y112_DO6;
  assign CLBLM_L_X70Y112_SLICE_X105Y112_AMUX = CLBLM_L_X70Y112_SLICE_X105Y112_A5Q;
  assign CLBLM_L_X70Y112_SLICE_X105Y112_BMUX = CLBLM_L_X70Y112_SLICE_X105Y112_B5Q;
  assign CLBLM_L_X70Y112_SLICE_X105Y112_CMUX = CLBLM_L_X70Y112_SLICE_X105Y112_C5Q;
  assign CLBLM_L_X70Y112_SLICE_X105Y112_DMUX = CLBLM_L_X70Y112_SLICE_X105Y112_D5Q;
  assign CLBLM_L_X70Y113_SLICE_X104Y113_A = CLBLM_L_X70Y113_SLICE_X104Y113_AO6;
  assign CLBLM_L_X70Y113_SLICE_X104Y113_B = CLBLM_L_X70Y113_SLICE_X104Y113_BO6;
  assign CLBLM_L_X70Y113_SLICE_X104Y113_C = CLBLM_L_X70Y113_SLICE_X104Y113_CO6;
  assign CLBLM_L_X70Y113_SLICE_X104Y113_D = CLBLM_L_X70Y113_SLICE_X104Y113_DO6;
  assign CLBLM_L_X70Y113_SLICE_X104Y113_AMUX = CLBLM_L_X70Y113_SLICE_X104Y113_A5Q;
  assign CLBLM_L_X70Y113_SLICE_X104Y113_BMUX = CLBLM_L_X70Y113_SLICE_X104Y113_B5Q;
  assign CLBLM_L_X70Y113_SLICE_X105Y113_A = CLBLM_L_X70Y113_SLICE_X105Y113_AO6;
  assign CLBLM_L_X70Y113_SLICE_X105Y113_B = CLBLM_L_X70Y113_SLICE_X105Y113_BO6;
  assign CLBLM_L_X70Y113_SLICE_X105Y113_C = CLBLM_L_X70Y113_SLICE_X105Y113_CO6;
  assign CLBLM_L_X70Y113_SLICE_X105Y113_D = CLBLM_L_X70Y113_SLICE_X105Y113_DO6;
  assign CLBLM_L_X70Y114_SLICE_X104Y114_A = CLBLM_L_X70Y114_SLICE_X104Y114_AO6;
  assign CLBLM_L_X70Y114_SLICE_X104Y114_B = CLBLM_L_X70Y114_SLICE_X104Y114_BO6;
  assign CLBLM_L_X70Y114_SLICE_X104Y114_C = CLBLM_L_X70Y114_SLICE_X104Y114_CO6;
  assign CLBLM_L_X70Y114_SLICE_X104Y114_D = CLBLM_L_X70Y114_SLICE_X104Y114_DO6;
  assign CLBLM_L_X70Y114_SLICE_X104Y114_AMUX = CLBLM_L_X70Y114_SLICE_X104Y114_A5Q;
  assign CLBLM_L_X70Y114_SLICE_X105Y114_A = CLBLM_L_X70Y114_SLICE_X105Y114_AO6;
  assign CLBLM_L_X70Y114_SLICE_X105Y114_B = CLBLM_L_X70Y114_SLICE_X105Y114_BO6;
  assign CLBLM_L_X70Y114_SLICE_X105Y114_C = CLBLM_L_X70Y114_SLICE_X105Y114_CO6;
  assign CLBLM_L_X70Y114_SLICE_X105Y114_D = CLBLM_L_X70Y114_SLICE_X105Y114_DO6;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_A = CLBLM_L_X70Y119_SLICE_X104Y119_AO6;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_B = CLBLM_L_X70Y119_SLICE_X104Y119_BO6;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_C = CLBLM_L_X70Y119_SLICE_X104Y119_CO6;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_D = CLBLM_L_X70Y119_SLICE_X104Y119_DO6;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_A = CLBLM_L_X70Y119_SLICE_X105Y119_AO6;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_B = CLBLM_L_X70Y119_SLICE_X105Y119_BO6;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_C = CLBLM_L_X70Y119_SLICE_X105Y119_CO6;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_D = CLBLM_L_X70Y119_SLICE_X105Y119_DO6;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_AMUX = CLBLM_L_X70Y119_SLICE_X105Y119_A5Q;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_A = CLBLM_L_X70Y123_SLICE_X104Y123_AO6;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_B = CLBLM_L_X70Y123_SLICE_X104Y123_BO6;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_C = CLBLM_L_X70Y123_SLICE_X104Y123_CO6;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_D = CLBLM_L_X70Y123_SLICE_X104Y123_DO6;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_AMUX = CLBLM_L_X70Y123_SLICE_X104Y123_A5Q;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_A = CLBLM_L_X70Y123_SLICE_X105Y123_AO6;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_B = CLBLM_L_X70Y123_SLICE_X105Y123_BO6;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_C = CLBLM_L_X70Y123_SLICE_X105Y123_CO6;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_D = CLBLM_L_X70Y123_SLICE_X105Y123_DO6;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_A = CLBLM_L_X70Y124_SLICE_X104Y124_AO6;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_B = CLBLM_L_X70Y124_SLICE_X104Y124_BO6;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_C = CLBLM_L_X70Y124_SLICE_X104Y124_CO6;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_D = CLBLM_L_X70Y124_SLICE_X104Y124_DO6;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_A = CLBLM_L_X70Y124_SLICE_X105Y124_AO6;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_B = CLBLM_L_X70Y124_SLICE_X105Y124_BO6;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_C = CLBLM_L_X70Y124_SLICE_X105Y124_CO6;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_D = CLBLM_L_X70Y124_SLICE_X105Y124_DO6;
  assign CLBLM_L_X70Y125_SLICE_X104Y125_A = CLBLM_L_X70Y125_SLICE_X104Y125_AO6;
  assign CLBLM_L_X70Y125_SLICE_X104Y125_B = CLBLM_L_X70Y125_SLICE_X104Y125_BO6;
  assign CLBLM_L_X70Y125_SLICE_X104Y125_C = CLBLM_L_X70Y125_SLICE_X104Y125_CO6;
  assign CLBLM_L_X70Y125_SLICE_X104Y125_D = CLBLM_L_X70Y125_SLICE_X104Y125_DO6;
  assign CLBLM_L_X70Y125_SLICE_X104Y125_AMUX = CLBLM_L_X70Y125_SLICE_X104Y125_A5Q;
  assign CLBLM_L_X70Y125_SLICE_X105Y125_A = CLBLM_L_X70Y125_SLICE_X105Y125_AO6;
  assign CLBLM_L_X70Y125_SLICE_X105Y125_B = CLBLM_L_X70Y125_SLICE_X105Y125_BO6;
  assign CLBLM_L_X70Y125_SLICE_X105Y125_C = CLBLM_L_X70Y125_SLICE_X105Y125_CO6;
  assign CLBLM_L_X70Y125_SLICE_X105Y125_D = CLBLM_L_X70Y125_SLICE_X105Y125_DO6;
  assign CLBLM_L_X70Y125_SLICE_X105Y125_AMUX = CLBLM_L_X70Y125_SLICE_X105Y125_AO5;
  assign CLBLM_L_X70Y125_SLICE_X105Y125_BMUX = CLBLM_L_X70Y125_SLICE_X105Y125_BO5;
  assign CLBLM_L_X70Y125_SLICE_X105Y125_CMUX = CLBLM_L_X70Y125_SLICE_X105Y125_CO6;
  assign CLBLM_L_X70Y126_SLICE_X104Y126_A = CLBLM_L_X70Y126_SLICE_X104Y126_AO6;
  assign CLBLM_L_X70Y126_SLICE_X104Y126_B = CLBLM_L_X70Y126_SLICE_X104Y126_BO6;
  assign CLBLM_L_X70Y126_SLICE_X104Y126_C = CLBLM_L_X70Y126_SLICE_X104Y126_CO6;
  assign CLBLM_L_X70Y126_SLICE_X104Y126_D = CLBLM_L_X70Y126_SLICE_X104Y126_DO6;
  assign CLBLM_L_X70Y126_SLICE_X105Y126_A = CLBLM_L_X70Y126_SLICE_X105Y126_AO6;
  assign CLBLM_L_X70Y126_SLICE_X105Y126_B = CLBLM_L_X70Y126_SLICE_X105Y126_BO6;
  assign CLBLM_L_X70Y126_SLICE_X105Y126_C = CLBLM_L_X70Y126_SLICE_X105Y126_CO6;
  assign CLBLM_L_X70Y126_SLICE_X105Y126_D = CLBLM_L_X70Y126_SLICE_X105Y126_DO6;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_A = CLBLM_L_X70Y128_SLICE_X104Y128_AO6;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_B = CLBLM_L_X70Y128_SLICE_X104Y128_BO6;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_C = CLBLM_L_X70Y128_SLICE_X104Y128_CO6;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_D = CLBLM_L_X70Y128_SLICE_X104Y128_DO6;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_AMUX = CLBLM_L_X70Y128_SLICE_X104Y128_AO5;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_BMUX = CLBLM_L_X70Y128_SLICE_X104Y128_BO5;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_A = CLBLM_L_X70Y128_SLICE_X105Y128_AO6;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_B = CLBLM_L_X70Y128_SLICE_X105Y128_BO6;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_C = CLBLM_L_X70Y128_SLICE_X105Y128_CO6;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_D = CLBLM_L_X70Y128_SLICE_X105Y128_DO6;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_BMUX = CLBLM_L_X70Y128_SLICE_X105Y128_BO6;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_A = CLBLM_L_X70Y129_SLICE_X104Y129_AO6;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_B = CLBLM_L_X70Y129_SLICE_X104Y129_BO6;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_C = CLBLM_L_X70Y129_SLICE_X104Y129_CO6;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_D = CLBLM_L_X70Y129_SLICE_X104Y129_DO6;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_A = CLBLM_L_X70Y129_SLICE_X105Y129_AO6;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_B = CLBLM_L_X70Y129_SLICE_X105Y129_BO6;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_C = CLBLM_L_X70Y129_SLICE_X105Y129_CO6;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_D = CLBLM_L_X70Y129_SLICE_X105Y129_DO6;
  assign CLBLM_L_X70Y130_SLICE_X104Y130_A = CLBLM_L_X70Y130_SLICE_X104Y130_AO6;
  assign CLBLM_L_X70Y130_SLICE_X104Y130_B = CLBLM_L_X70Y130_SLICE_X104Y130_BO6;
  assign CLBLM_L_X70Y130_SLICE_X104Y130_C = CLBLM_L_X70Y130_SLICE_X104Y130_CO6;
  assign CLBLM_L_X70Y130_SLICE_X104Y130_D = CLBLM_L_X70Y130_SLICE_X104Y130_DO6;
  assign CLBLM_L_X70Y130_SLICE_X104Y130_AMUX = CLBLM_L_X70Y130_SLICE_X104Y130_AO5;
  assign CLBLM_L_X70Y130_SLICE_X105Y130_A = CLBLM_L_X70Y130_SLICE_X105Y130_AO6;
  assign CLBLM_L_X70Y130_SLICE_X105Y130_B = CLBLM_L_X70Y130_SLICE_X105Y130_BO6;
  assign CLBLM_L_X70Y130_SLICE_X105Y130_C = CLBLM_L_X70Y130_SLICE_X105Y130_CO6;
  assign CLBLM_L_X70Y130_SLICE_X105Y130_D = CLBLM_L_X70Y130_SLICE_X105Y130_DO6;
  assign CLBLM_L_X70Y130_SLICE_X105Y130_AMUX = CLBLM_L_X70Y130_SLICE_X105Y130_A5Q;
  assign CLBLM_L_X70Y130_SLICE_X105Y130_DMUX = CLBLM_L_X70Y130_SLICE_X105Y130_DO5;
  assign CLBLM_L_X70Y131_SLICE_X104Y131_A = CLBLM_L_X70Y131_SLICE_X104Y131_AO6;
  assign CLBLM_L_X70Y131_SLICE_X104Y131_B = CLBLM_L_X70Y131_SLICE_X104Y131_BO6;
  assign CLBLM_L_X70Y131_SLICE_X104Y131_C = CLBLM_L_X70Y131_SLICE_X104Y131_CO6;
  assign CLBLM_L_X70Y131_SLICE_X104Y131_D = CLBLM_L_X70Y131_SLICE_X104Y131_DO6;
  assign CLBLM_L_X70Y131_SLICE_X105Y131_A = CLBLM_L_X70Y131_SLICE_X105Y131_AO6;
  assign CLBLM_L_X70Y131_SLICE_X105Y131_B = CLBLM_L_X70Y131_SLICE_X105Y131_BO6;
  assign CLBLM_L_X70Y131_SLICE_X105Y131_C = CLBLM_L_X70Y131_SLICE_X105Y131_CO6;
  assign CLBLM_L_X70Y131_SLICE_X105Y131_D = CLBLM_L_X70Y131_SLICE_X105Y131_DO6;
  assign CLBLM_L_X70Y132_SLICE_X104Y132_A = CLBLM_L_X70Y132_SLICE_X104Y132_AO6;
  assign CLBLM_L_X70Y132_SLICE_X104Y132_B = CLBLM_L_X70Y132_SLICE_X104Y132_BO6;
  assign CLBLM_L_X70Y132_SLICE_X104Y132_C = CLBLM_L_X70Y132_SLICE_X104Y132_CO6;
  assign CLBLM_L_X70Y132_SLICE_X104Y132_D = CLBLM_L_X70Y132_SLICE_X104Y132_DO6;
  assign CLBLM_L_X70Y132_SLICE_X105Y132_A = CLBLM_L_X70Y132_SLICE_X105Y132_AO6;
  assign CLBLM_L_X70Y132_SLICE_X105Y132_B = CLBLM_L_X70Y132_SLICE_X105Y132_BO6;
  assign CLBLM_L_X70Y132_SLICE_X105Y132_C = CLBLM_L_X70Y132_SLICE_X105Y132_CO6;
  assign CLBLM_L_X70Y132_SLICE_X105Y132_D = CLBLM_L_X70Y132_SLICE_X105Y132_DO6;
  assign CLBLM_L_X70Y133_SLICE_X104Y133_A = CLBLM_L_X70Y133_SLICE_X104Y133_AO6;
  assign CLBLM_L_X70Y133_SLICE_X104Y133_B = CLBLM_L_X70Y133_SLICE_X104Y133_BO6;
  assign CLBLM_L_X70Y133_SLICE_X104Y133_C = CLBLM_L_X70Y133_SLICE_X104Y133_CO6;
  assign CLBLM_L_X70Y133_SLICE_X104Y133_D = CLBLM_L_X70Y133_SLICE_X104Y133_DO6;
  assign CLBLM_L_X70Y133_SLICE_X104Y133_AMUX = CLBLM_L_X70Y133_SLICE_X104Y133_A5Q;
  assign CLBLM_L_X70Y133_SLICE_X104Y133_CMUX = CLBLM_L_X70Y133_SLICE_X104Y133_CO5;
  assign CLBLM_L_X70Y133_SLICE_X105Y133_A = CLBLM_L_X70Y133_SLICE_X105Y133_AO6;
  assign CLBLM_L_X70Y133_SLICE_X105Y133_B = CLBLM_L_X70Y133_SLICE_X105Y133_BO6;
  assign CLBLM_L_X70Y133_SLICE_X105Y133_C = CLBLM_L_X70Y133_SLICE_X105Y133_CO6;
  assign CLBLM_L_X70Y133_SLICE_X105Y133_D = CLBLM_L_X70Y133_SLICE_X105Y133_DO6;
  assign CLBLM_L_X70Y134_SLICE_X104Y134_A = CLBLM_L_X70Y134_SLICE_X104Y134_AO6;
  assign CLBLM_L_X70Y134_SLICE_X104Y134_B = CLBLM_L_X70Y134_SLICE_X104Y134_BO6;
  assign CLBLM_L_X70Y134_SLICE_X104Y134_C = CLBLM_L_X70Y134_SLICE_X104Y134_CO6;
  assign CLBLM_L_X70Y134_SLICE_X104Y134_D = CLBLM_L_X70Y134_SLICE_X104Y134_DO6;
  assign CLBLM_L_X70Y134_SLICE_X104Y134_CMUX = CLBLM_L_X70Y134_SLICE_X104Y134_CO5;
  assign CLBLM_L_X70Y134_SLICE_X105Y134_A = CLBLM_L_X70Y134_SLICE_X105Y134_AO6;
  assign CLBLM_L_X70Y134_SLICE_X105Y134_B = CLBLM_L_X70Y134_SLICE_X105Y134_BO6;
  assign CLBLM_L_X70Y134_SLICE_X105Y134_C = CLBLM_L_X70Y134_SLICE_X105Y134_CO6;
  assign CLBLM_L_X70Y134_SLICE_X105Y134_D = CLBLM_L_X70Y134_SLICE_X105Y134_DO6;
  assign CLBLM_L_X70Y134_SLICE_X105Y134_DMUX = CLBLM_L_X70Y134_SLICE_X105Y134_DO5;
  assign CLBLM_L_X70Y135_SLICE_X104Y135_A = CLBLM_L_X70Y135_SLICE_X104Y135_AO6;
  assign CLBLM_L_X70Y135_SLICE_X104Y135_B = CLBLM_L_X70Y135_SLICE_X104Y135_BO6;
  assign CLBLM_L_X70Y135_SLICE_X104Y135_C = CLBLM_L_X70Y135_SLICE_X104Y135_CO6;
  assign CLBLM_L_X70Y135_SLICE_X104Y135_D = CLBLM_L_X70Y135_SLICE_X104Y135_DO6;
  assign CLBLM_L_X70Y135_SLICE_X104Y135_CMUX = CLBLM_L_X70Y135_SLICE_X104Y135_CO5;
  assign CLBLM_L_X70Y135_SLICE_X105Y135_A = CLBLM_L_X70Y135_SLICE_X105Y135_AO6;
  assign CLBLM_L_X70Y135_SLICE_X105Y135_B = CLBLM_L_X70Y135_SLICE_X105Y135_BO6;
  assign CLBLM_L_X70Y135_SLICE_X105Y135_C = CLBLM_L_X70Y135_SLICE_X105Y135_CO6;
  assign CLBLM_L_X70Y135_SLICE_X105Y135_D = CLBLM_L_X70Y135_SLICE_X105Y135_DO6;
  assign CLBLM_L_X70Y135_SLICE_X105Y135_AMUX = CLBLM_L_X70Y135_SLICE_X105Y135_A5Q;
  assign CLBLM_L_X70Y136_SLICE_X104Y136_A = CLBLM_L_X70Y136_SLICE_X104Y136_AO6;
  assign CLBLM_L_X70Y136_SLICE_X104Y136_B = CLBLM_L_X70Y136_SLICE_X104Y136_BO6;
  assign CLBLM_L_X70Y136_SLICE_X104Y136_C = CLBLM_L_X70Y136_SLICE_X104Y136_CO6;
  assign CLBLM_L_X70Y136_SLICE_X104Y136_D = CLBLM_L_X70Y136_SLICE_X104Y136_DO6;
  assign CLBLM_L_X70Y136_SLICE_X105Y136_A = CLBLM_L_X70Y136_SLICE_X105Y136_AO6;
  assign CLBLM_L_X70Y136_SLICE_X105Y136_B = CLBLM_L_X70Y136_SLICE_X105Y136_BO6;
  assign CLBLM_L_X70Y136_SLICE_X105Y136_C = CLBLM_L_X70Y136_SLICE_X105Y136_CO6;
  assign CLBLM_L_X70Y136_SLICE_X105Y136_D = CLBLM_L_X70Y136_SLICE_X105Y136_DO6;
  assign CLBLM_L_X70Y136_SLICE_X105Y136_AMUX = CLBLM_L_X70Y136_SLICE_X105Y136_A5Q;
  assign CLBLM_L_X70Y136_SLICE_X105Y136_BMUX = CLBLM_L_X70Y136_SLICE_X105Y136_BO5;
  assign CLBLM_L_X72Y98_SLICE_X108Y98_A = CLBLM_L_X72Y98_SLICE_X108Y98_AO6;
  assign CLBLM_L_X72Y98_SLICE_X108Y98_B = CLBLM_L_X72Y98_SLICE_X108Y98_BO6;
  assign CLBLM_L_X72Y98_SLICE_X108Y98_C = CLBLM_L_X72Y98_SLICE_X108Y98_CO6;
  assign CLBLM_L_X72Y98_SLICE_X108Y98_D = CLBLM_L_X72Y98_SLICE_X108Y98_DO6;
  assign CLBLM_L_X72Y98_SLICE_X108Y98_AMUX = CLBLM_L_X72Y98_SLICE_X108Y98_A5Q;
  assign CLBLM_L_X72Y98_SLICE_X108Y98_BMUX = CLBLM_L_X72Y98_SLICE_X108Y98_B5Q;
  assign CLBLM_L_X72Y98_SLICE_X109Y98_A = CLBLM_L_X72Y98_SLICE_X109Y98_AO6;
  assign CLBLM_L_X72Y98_SLICE_X109Y98_B = CLBLM_L_X72Y98_SLICE_X109Y98_BO6;
  assign CLBLM_L_X72Y98_SLICE_X109Y98_C = CLBLM_L_X72Y98_SLICE_X109Y98_CO6;
  assign CLBLM_L_X72Y98_SLICE_X109Y98_D = CLBLM_L_X72Y98_SLICE_X109Y98_DO6;
  assign CLBLM_L_X72Y103_SLICE_X108Y103_A = CLBLM_L_X72Y103_SLICE_X108Y103_AO6;
  assign CLBLM_L_X72Y103_SLICE_X108Y103_B = CLBLM_L_X72Y103_SLICE_X108Y103_BO6;
  assign CLBLM_L_X72Y103_SLICE_X108Y103_C = CLBLM_L_X72Y103_SLICE_X108Y103_CO6;
  assign CLBLM_L_X72Y103_SLICE_X108Y103_D = CLBLM_L_X72Y103_SLICE_X108Y103_DO6;
  assign CLBLM_L_X72Y103_SLICE_X108Y103_AMUX = CLBLM_L_X72Y103_SLICE_X108Y103_A5Q;
  assign CLBLM_L_X72Y103_SLICE_X108Y103_BMUX = CLBLM_L_X72Y103_SLICE_X108Y103_BO5;
  assign CLBLM_L_X72Y103_SLICE_X108Y103_CMUX = CLBLM_L_X72Y103_SLICE_X108Y103_CO5;
  assign CLBLM_L_X72Y103_SLICE_X108Y103_DMUX = CLBLM_L_X72Y103_SLICE_X108Y103_DO5;
  assign CLBLM_L_X72Y103_SLICE_X109Y103_A = CLBLM_L_X72Y103_SLICE_X109Y103_AO6;
  assign CLBLM_L_X72Y103_SLICE_X109Y103_B = CLBLM_L_X72Y103_SLICE_X109Y103_BO6;
  assign CLBLM_L_X72Y103_SLICE_X109Y103_C = CLBLM_L_X72Y103_SLICE_X109Y103_CO6;
  assign CLBLM_L_X72Y103_SLICE_X109Y103_D = CLBLM_L_X72Y103_SLICE_X109Y103_DO6;
  assign CLBLM_L_X72Y103_SLICE_X109Y103_AMUX = CLBLM_L_X72Y103_SLICE_X109Y103_AO5;
  assign CLBLM_L_X72Y104_SLICE_X108Y104_A = CLBLM_L_X72Y104_SLICE_X108Y104_AO6;
  assign CLBLM_L_X72Y104_SLICE_X108Y104_B = CLBLM_L_X72Y104_SLICE_X108Y104_BO6;
  assign CLBLM_L_X72Y104_SLICE_X108Y104_C = CLBLM_L_X72Y104_SLICE_X108Y104_CO6;
  assign CLBLM_L_X72Y104_SLICE_X108Y104_D = CLBLM_L_X72Y104_SLICE_X108Y104_DO6;
  assign CLBLM_L_X72Y104_SLICE_X109Y104_A = CLBLM_L_X72Y104_SLICE_X109Y104_AO6;
  assign CLBLM_L_X72Y104_SLICE_X109Y104_B = CLBLM_L_X72Y104_SLICE_X109Y104_BO6;
  assign CLBLM_L_X72Y104_SLICE_X109Y104_C = CLBLM_L_X72Y104_SLICE_X109Y104_CO6;
  assign CLBLM_L_X72Y104_SLICE_X109Y104_D = CLBLM_L_X72Y104_SLICE_X109Y104_DO6;
  assign CLBLM_L_X72Y104_SLICE_X109Y104_AMUX = CLBLM_L_X72Y104_SLICE_X109Y104_A5Q;
  assign CLBLM_L_X72Y104_SLICE_X109Y104_BMUX = CLBLM_L_X72Y104_SLICE_X109Y104_B5Q;
  assign CLBLM_L_X72Y104_SLICE_X109Y104_CMUX = CLBLM_L_X72Y104_SLICE_X109Y104_C5Q;
  assign CLBLM_L_X72Y105_SLICE_X108Y105_A = CLBLM_L_X72Y105_SLICE_X108Y105_AO6;
  assign CLBLM_L_X72Y105_SLICE_X108Y105_B = CLBLM_L_X72Y105_SLICE_X108Y105_BO6;
  assign CLBLM_L_X72Y105_SLICE_X108Y105_C = CLBLM_L_X72Y105_SLICE_X108Y105_CO6;
  assign CLBLM_L_X72Y105_SLICE_X108Y105_D = CLBLM_L_X72Y105_SLICE_X108Y105_DO6;
  assign CLBLM_L_X72Y105_SLICE_X108Y105_AMUX = CLBLM_L_X72Y105_SLICE_X108Y105_A5Q;
  assign CLBLM_L_X72Y105_SLICE_X109Y105_A = CLBLM_L_X72Y105_SLICE_X109Y105_AO6;
  assign CLBLM_L_X72Y105_SLICE_X109Y105_B = CLBLM_L_X72Y105_SLICE_X109Y105_BO6;
  assign CLBLM_L_X72Y105_SLICE_X109Y105_C = CLBLM_L_X72Y105_SLICE_X109Y105_CO6;
  assign CLBLM_L_X72Y105_SLICE_X109Y105_D = CLBLM_L_X72Y105_SLICE_X109Y105_DO6;
  assign CLBLM_L_X72Y105_SLICE_X109Y105_BMUX = CLBLM_L_X72Y105_SLICE_X109Y105_B5Q;
  assign CLBLM_L_X72Y106_SLICE_X108Y106_A = CLBLM_L_X72Y106_SLICE_X108Y106_AO6;
  assign CLBLM_L_X72Y106_SLICE_X108Y106_B = CLBLM_L_X72Y106_SLICE_X108Y106_BO6;
  assign CLBLM_L_X72Y106_SLICE_X108Y106_C = CLBLM_L_X72Y106_SLICE_X108Y106_CO6;
  assign CLBLM_L_X72Y106_SLICE_X108Y106_D = CLBLM_L_X72Y106_SLICE_X108Y106_DO6;
  assign CLBLM_L_X72Y106_SLICE_X108Y106_AMUX = CLBLM_L_X72Y106_SLICE_X108Y106_A5Q;
  assign CLBLM_L_X72Y106_SLICE_X108Y106_BMUX = CLBLM_L_X72Y106_SLICE_X108Y106_BO6;
  assign CLBLM_L_X72Y106_SLICE_X108Y106_DMUX = CLBLM_L_X72Y106_SLICE_X108Y106_DO6;
  assign CLBLM_L_X72Y106_SLICE_X109Y106_A = CLBLM_L_X72Y106_SLICE_X109Y106_AO6;
  assign CLBLM_L_X72Y106_SLICE_X109Y106_B = CLBLM_L_X72Y106_SLICE_X109Y106_BO6;
  assign CLBLM_L_X72Y106_SLICE_X109Y106_C = CLBLM_L_X72Y106_SLICE_X109Y106_CO6;
  assign CLBLM_L_X72Y106_SLICE_X109Y106_D = CLBLM_L_X72Y106_SLICE_X109Y106_DO6;
  assign CLBLM_L_X72Y107_SLICE_X108Y107_A = CLBLM_L_X72Y107_SLICE_X108Y107_AO6;
  assign CLBLM_L_X72Y107_SLICE_X108Y107_B = CLBLM_L_X72Y107_SLICE_X108Y107_BO6;
  assign CLBLM_L_X72Y107_SLICE_X108Y107_C = CLBLM_L_X72Y107_SLICE_X108Y107_CO6;
  assign CLBLM_L_X72Y107_SLICE_X108Y107_D = CLBLM_L_X72Y107_SLICE_X108Y107_DO6;
  assign CLBLM_L_X72Y107_SLICE_X108Y107_AMUX = CLBLM_L_X72Y107_SLICE_X108Y107_A5Q;
  assign CLBLM_L_X72Y107_SLICE_X108Y107_BMUX = CLBLM_L_X72Y107_SLICE_X108Y107_BO5;
  assign CLBLM_L_X72Y107_SLICE_X109Y107_A = CLBLM_L_X72Y107_SLICE_X109Y107_AO6;
  assign CLBLM_L_X72Y107_SLICE_X109Y107_B = CLBLM_L_X72Y107_SLICE_X109Y107_BO6;
  assign CLBLM_L_X72Y107_SLICE_X109Y107_C = CLBLM_L_X72Y107_SLICE_X109Y107_CO6;
  assign CLBLM_L_X72Y107_SLICE_X109Y107_D = CLBLM_L_X72Y107_SLICE_X109Y107_DO6;
  assign CLBLM_L_X72Y107_SLICE_X109Y107_AMUX = CLBLM_L_X72Y107_SLICE_X109Y107_A5Q;
  assign CLBLM_L_X72Y107_SLICE_X109Y107_BMUX = CLBLM_L_X72Y107_SLICE_X109Y107_BO5;
  assign CLBLM_L_X72Y108_SLICE_X108Y108_A = CLBLM_L_X72Y108_SLICE_X108Y108_AO6;
  assign CLBLM_L_X72Y108_SLICE_X108Y108_B = CLBLM_L_X72Y108_SLICE_X108Y108_BO6;
  assign CLBLM_L_X72Y108_SLICE_X108Y108_C = CLBLM_L_X72Y108_SLICE_X108Y108_CO6;
  assign CLBLM_L_X72Y108_SLICE_X108Y108_D = CLBLM_L_X72Y108_SLICE_X108Y108_DO6;
  assign CLBLM_L_X72Y108_SLICE_X108Y108_BMUX = CLBLM_L_X72Y108_SLICE_X108Y108_BO5;
  assign CLBLM_L_X72Y108_SLICE_X109Y108_A = CLBLM_L_X72Y108_SLICE_X109Y108_AO6;
  assign CLBLM_L_X72Y108_SLICE_X109Y108_B = CLBLM_L_X72Y108_SLICE_X109Y108_BO6;
  assign CLBLM_L_X72Y108_SLICE_X109Y108_C = CLBLM_L_X72Y108_SLICE_X109Y108_CO6;
  assign CLBLM_L_X72Y108_SLICE_X109Y108_D = CLBLM_L_X72Y108_SLICE_X109Y108_DO6;
  assign CLBLM_L_X72Y108_SLICE_X109Y108_AMUX = CLBLM_L_X72Y108_SLICE_X109Y108_A5Q;
  assign CLBLM_L_X72Y108_SLICE_X109Y108_BMUX = CLBLM_L_X72Y108_SLICE_X109Y108_BO5;
  assign CLBLM_L_X72Y108_SLICE_X109Y108_CMUX = CLBLM_L_X72Y108_SLICE_X109Y108_CO5;
  assign CLBLM_L_X72Y109_SLICE_X108Y109_A = CLBLM_L_X72Y109_SLICE_X108Y109_AO6;
  assign CLBLM_L_X72Y109_SLICE_X108Y109_B = CLBLM_L_X72Y109_SLICE_X108Y109_BO6;
  assign CLBLM_L_X72Y109_SLICE_X108Y109_C = CLBLM_L_X72Y109_SLICE_X108Y109_CO6;
  assign CLBLM_L_X72Y109_SLICE_X108Y109_D = CLBLM_L_X72Y109_SLICE_X108Y109_DO6;
  assign CLBLM_L_X72Y109_SLICE_X109Y109_A = CLBLM_L_X72Y109_SLICE_X109Y109_AO6;
  assign CLBLM_L_X72Y109_SLICE_X109Y109_B = CLBLM_L_X72Y109_SLICE_X109Y109_BO6;
  assign CLBLM_L_X72Y109_SLICE_X109Y109_C = CLBLM_L_X72Y109_SLICE_X109Y109_CO6;
  assign CLBLM_L_X72Y109_SLICE_X109Y109_D = CLBLM_L_X72Y109_SLICE_X109Y109_DO6;
  assign CLBLM_L_X72Y109_SLICE_X109Y109_AMUX = CLBLM_L_X72Y109_SLICE_X109Y109_A5Q;
  assign CLBLM_L_X72Y109_SLICE_X109Y109_BMUX = CLBLM_L_X72Y109_SLICE_X109Y109_B5Q;
  assign CLBLM_L_X72Y109_SLICE_X109Y109_CMUX = CLBLM_L_X72Y109_SLICE_X109Y109_C5Q;
  assign CLBLM_L_X72Y111_SLICE_X108Y111_A = CLBLM_L_X72Y111_SLICE_X108Y111_AO6;
  assign CLBLM_L_X72Y111_SLICE_X108Y111_B = CLBLM_L_X72Y111_SLICE_X108Y111_BO6;
  assign CLBLM_L_X72Y111_SLICE_X108Y111_C = CLBLM_L_X72Y111_SLICE_X108Y111_CO6;
  assign CLBLM_L_X72Y111_SLICE_X108Y111_D = CLBLM_L_X72Y111_SLICE_X108Y111_DO6;
  assign CLBLM_L_X72Y111_SLICE_X108Y111_AMUX = CLBLM_L_X72Y111_SLICE_X108Y111_AO5;
  assign CLBLM_L_X72Y111_SLICE_X108Y111_CMUX = CLBLM_L_X72Y111_SLICE_X108Y111_C5Q;
  assign CLBLM_L_X72Y111_SLICE_X109Y111_A = CLBLM_L_X72Y111_SLICE_X109Y111_AO6;
  assign CLBLM_L_X72Y111_SLICE_X109Y111_B = CLBLM_L_X72Y111_SLICE_X109Y111_BO6;
  assign CLBLM_L_X72Y111_SLICE_X109Y111_C = CLBLM_L_X72Y111_SLICE_X109Y111_CO6;
  assign CLBLM_L_X72Y111_SLICE_X109Y111_D = CLBLM_L_X72Y111_SLICE_X109Y111_DO6;
  assign CLBLM_L_X72Y111_SLICE_X109Y111_AMUX = CLBLM_L_X72Y111_SLICE_X109Y111_A5Q;
  assign CLBLM_L_X72Y113_SLICE_X108Y113_A = CLBLM_L_X72Y113_SLICE_X108Y113_AO6;
  assign CLBLM_L_X72Y113_SLICE_X108Y113_B = CLBLM_L_X72Y113_SLICE_X108Y113_BO6;
  assign CLBLM_L_X72Y113_SLICE_X108Y113_C = CLBLM_L_X72Y113_SLICE_X108Y113_CO6;
  assign CLBLM_L_X72Y113_SLICE_X108Y113_D = CLBLM_L_X72Y113_SLICE_X108Y113_DO6;
  assign CLBLM_L_X72Y113_SLICE_X109Y113_A = CLBLM_L_X72Y113_SLICE_X109Y113_AO6;
  assign CLBLM_L_X72Y113_SLICE_X109Y113_B = CLBLM_L_X72Y113_SLICE_X109Y113_BO6;
  assign CLBLM_L_X72Y113_SLICE_X109Y113_C = CLBLM_L_X72Y113_SLICE_X109Y113_CO6;
  assign CLBLM_L_X72Y113_SLICE_X109Y113_D = CLBLM_L_X72Y113_SLICE_X109Y113_DO6;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_A = CLBLM_L_X72Y116_SLICE_X108Y116_AO6;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_B = CLBLM_L_X72Y116_SLICE_X108Y116_BO6;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_C = CLBLM_L_X72Y116_SLICE_X108Y116_CO6;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_D = CLBLM_L_X72Y116_SLICE_X108Y116_DO6;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_A = CLBLM_L_X72Y116_SLICE_X109Y116_AO6;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_B = CLBLM_L_X72Y116_SLICE_X109Y116_BO6;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_C = CLBLM_L_X72Y116_SLICE_X109Y116_CO6;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_D = CLBLM_L_X72Y116_SLICE_X109Y116_DO6;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_A = CLBLM_L_X72Y117_SLICE_X108Y117_AO6;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_B = CLBLM_L_X72Y117_SLICE_X108Y117_BO6;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_C = CLBLM_L_X72Y117_SLICE_X108Y117_CO6;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_D = CLBLM_L_X72Y117_SLICE_X108Y117_DO6;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_A = CLBLM_L_X72Y117_SLICE_X109Y117_AO6;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_B = CLBLM_L_X72Y117_SLICE_X109Y117_BO6;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_C = CLBLM_L_X72Y117_SLICE_X109Y117_CO6;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_D = CLBLM_L_X72Y117_SLICE_X109Y117_DO6;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_A = CLBLM_L_X72Y118_SLICE_X108Y118_AO6;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_B = CLBLM_L_X72Y118_SLICE_X108Y118_BO6;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_C = CLBLM_L_X72Y118_SLICE_X108Y118_CO6;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_D = CLBLM_L_X72Y118_SLICE_X108Y118_DO6;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_AMUX = CLBLM_L_X72Y118_SLICE_X108Y118_A5Q;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_BMUX = CLBLM_L_X72Y118_SLICE_X108Y118_B5Q;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_CMUX = CLBLM_L_X72Y118_SLICE_X108Y118_C5Q;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_DMUX = CLBLM_L_X72Y118_SLICE_X108Y118_D5Q;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_A = CLBLM_L_X72Y118_SLICE_X109Y118_AO6;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_B = CLBLM_L_X72Y118_SLICE_X109Y118_BO6;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_C = CLBLM_L_X72Y118_SLICE_X109Y118_CO6;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_D = CLBLM_L_X72Y118_SLICE_X109Y118_DO6;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_AMUX = CLBLM_L_X72Y118_SLICE_X109Y118_A5Q;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_A = CLBLM_L_X72Y119_SLICE_X108Y119_AO6;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_B = CLBLM_L_X72Y119_SLICE_X108Y119_BO6;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_C = CLBLM_L_X72Y119_SLICE_X108Y119_CO6;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_D = CLBLM_L_X72Y119_SLICE_X108Y119_DO6;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_AMUX = CLBLM_L_X72Y119_SLICE_X108Y119_A5Q;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_CMUX = CLBLM_L_X72Y119_SLICE_X108Y119_C5Q;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_A = CLBLM_L_X72Y119_SLICE_X109Y119_AO6;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_B = CLBLM_L_X72Y119_SLICE_X109Y119_BO6;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_C = CLBLM_L_X72Y119_SLICE_X109Y119_CO6;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_D = CLBLM_L_X72Y119_SLICE_X109Y119_DO6;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_AMUX = CLBLM_L_X72Y119_SLICE_X109Y119_A5Q;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_BMUX = CLBLM_L_X72Y119_SLICE_X109Y119_B5Q;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_CMUX = CLBLM_L_X72Y119_SLICE_X109Y119_CO6;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_DMUX = CLBLM_L_X72Y119_SLICE_X109Y119_DO6;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_A = CLBLM_L_X72Y120_SLICE_X108Y120_AO6;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_B = CLBLM_L_X72Y120_SLICE_X108Y120_BO6;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_C = CLBLM_L_X72Y120_SLICE_X108Y120_CO6;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_D = CLBLM_L_X72Y120_SLICE_X108Y120_DO6;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_AMUX = CLBLM_L_X72Y120_SLICE_X108Y120_A5Q;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_A = CLBLM_L_X72Y120_SLICE_X109Y120_AO6;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_B = CLBLM_L_X72Y120_SLICE_X109Y120_BO6;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_C = CLBLM_L_X72Y120_SLICE_X109Y120_CO6;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_D = CLBLM_L_X72Y120_SLICE_X109Y120_DO6;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_A = CLBLM_L_X72Y121_SLICE_X108Y121_AO6;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_B = CLBLM_L_X72Y121_SLICE_X108Y121_BO6;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_C = CLBLM_L_X72Y121_SLICE_X108Y121_CO6;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_D = CLBLM_L_X72Y121_SLICE_X108Y121_DO6;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_AMUX = CLBLM_L_X72Y121_SLICE_X108Y121_A5Q;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_A = CLBLM_L_X72Y121_SLICE_X109Y121_AO6;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_B = CLBLM_L_X72Y121_SLICE_X109Y121_BO6;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_C = CLBLM_L_X72Y121_SLICE_X109Y121_CO6;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_D = CLBLM_L_X72Y121_SLICE_X109Y121_DO6;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_AMUX = CLBLM_L_X72Y121_SLICE_X109Y121_A5Q;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_A = CLBLM_L_X72Y122_SLICE_X108Y122_AO6;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_B = CLBLM_L_X72Y122_SLICE_X108Y122_BO6;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_C = CLBLM_L_X72Y122_SLICE_X108Y122_CO6;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_D = CLBLM_L_X72Y122_SLICE_X108Y122_DO6;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_A = CLBLM_L_X72Y122_SLICE_X109Y122_AO6;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_B = CLBLM_L_X72Y122_SLICE_X109Y122_BO6;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_C = CLBLM_L_X72Y122_SLICE_X109Y122_CO6;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_D = CLBLM_L_X72Y122_SLICE_X109Y122_DO6;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_AMUX = CLBLM_L_X72Y122_SLICE_X109Y122_A5Q;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_CMUX = CLBLM_L_X72Y122_SLICE_X109Y122_CO5;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_A = CLBLM_L_X72Y123_SLICE_X108Y123_AO6;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_B = CLBLM_L_X72Y123_SLICE_X108Y123_BO6;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_C = CLBLM_L_X72Y123_SLICE_X108Y123_CO6;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_D = CLBLM_L_X72Y123_SLICE_X108Y123_DO6;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_AMUX = CLBLM_L_X72Y123_SLICE_X108Y123_A5Q;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_BMUX = CLBLM_L_X72Y123_SLICE_X108Y123_BO5;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_CMUX = CLBLM_L_X72Y123_SLICE_X108Y123_CO5;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_A = CLBLM_L_X72Y123_SLICE_X109Y123_AO6;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_B = CLBLM_L_X72Y123_SLICE_X109Y123_BO6;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_C = CLBLM_L_X72Y123_SLICE_X109Y123_CO6;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_D = CLBLM_L_X72Y123_SLICE_X109Y123_DO6;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_A = CLBLM_L_X72Y124_SLICE_X108Y124_AO6;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_B = CLBLM_L_X72Y124_SLICE_X108Y124_BO6;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_C = CLBLM_L_X72Y124_SLICE_X108Y124_CO6;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_D = CLBLM_L_X72Y124_SLICE_X108Y124_DO6;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_A = CLBLM_L_X72Y124_SLICE_X109Y124_AO6;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_B = CLBLM_L_X72Y124_SLICE_X109Y124_BO6;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_C = CLBLM_L_X72Y124_SLICE_X109Y124_CO6;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_D = CLBLM_L_X72Y124_SLICE_X109Y124_DO6;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_A = CLBLM_L_X72Y125_SLICE_X108Y125_AO6;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_B = CLBLM_L_X72Y125_SLICE_X108Y125_BO6;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_C = CLBLM_L_X72Y125_SLICE_X108Y125_CO6;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_D = CLBLM_L_X72Y125_SLICE_X108Y125_DO6;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_A = CLBLM_L_X72Y125_SLICE_X109Y125_AO6;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_B = CLBLM_L_X72Y125_SLICE_X109Y125_BO6;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_C = CLBLM_L_X72Y125_SLICE_X109Y125_CO6;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_D = CLBLM_L_X72Y125_SLICE_X109Y125_DO6;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_A = CLBLM_L_X72Y126_SLICE_X108Y126_AO6;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_B = CLBLM_L_X72Y126_SLICE_X108Y126_BO6;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_C = CLBLM_L_X72Y126_SLICE_X108Y126_CO6;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_D = CLBLM_L_X72Y126_SLICE_X108Y126_DO6;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_A = CLBLM_L_X72Y126_SLICE_X109Y126_AO6;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_B = CLBLM_L_X72Y126_SLICE_X109Y126_BO6;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_C = CLBLM_L_X72Y126_SLICE_X109Y126_CO6;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_D = CLBLM_L_X72Y126_SLICE_X109Y126_DO6;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_A = CLBLM_L_X72Y127_SLICE_X108Y127_AO6;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_B = CLBLM_L_X72Y127_SLICE_X108Y127_BO6;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_C = CLBLM_L_X72Y127_SLICE_X108Y127_CO6;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_D = CLBLM_L_X72Y127_SLICE_X108Y127_DO6;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_AMUX = CLBLM_L_X72Y127_SLICE_X108Y127_A5Q;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_BMUX = CLBLM_L_X72Y127_SLICE_X108Y127_BO5;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_A = CLBLM_L_X72Y127_SLICE_X109Y127_AO6;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_B = CLBLM_L_X72Y127_SLICE_X109Y127_BO6;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_C = CLBLM_L_X72Y127_SLICE_X109Y127_CO6;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_D = CLBLM_L_X72Y127_SLICE_X109Y127_DO6;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_A = CLBLM_L_X72Y128_SLICE_X108Y128_AO6;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_B = CLBLM_L_X72Y128_SLICE_X108Y128_BO6;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_C = CLBLM_L_X72Y128_SLICE_X108Y128_CO6;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_D = CLBLM_L_X72Y128_SLICE_X108Y128_DO6;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_AMUX = CLBLM_L_X72Y128_SLICE_X108Y128_A5Q;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_BMUX = CLBLM_L_X72Y128_SLICE_X108Y128_BO5;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_A = CLBLM_L_X72Y128_SLICE_X109Y128_AO6;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_B = CLBLM_L_X72Y128_SLICE_X109Y128_BO6;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_C = CLBLM_L_X72Y128_SLICE_X109Y128_CO6;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_D = CLBLM_L_X72Y128_SLICE_X109Y128_DO6;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_A = CLBLM_L_X72Y129_SLICE_X108Y129_AO6;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_B = CLBLM_L_X72Y129_SLICE_X108Y129_BO6;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_C = CLBLM_L_X72Y129_SLICE_X108Y129_CO6;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_D = CLBLM_L_X72Y129_SLICE_X108Y129_DO6;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_AMUX = CLBLM_L_X72Y129_SLICE_X108Y129_AO5;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_A = CLBLM_L_X72Y129_SLICE_X109Y129_AO6;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_B = CLBLM_L_X72Y129_SLICE_X109Y129_BO6;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_C = CLBLM_L_X72Y129_SLICE_X109Y129_CO6;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_D = CLBLM_L_X72Y129_SLICE_X109Y129_DO6;
  assign CLBLM_L_X72Y130_SLICE_X108Y130_A = CLBLM_L_X72Y130_SLICE_X108Y130_AO6;
  assign CLBLM_L_X72Y130_SLICE_X108Y130_B = CLBLM_L_X72Y130_SLICE_X108Y130_BO6;
  assign CLBLM_L_X72Y130_SLICE_X108Y130_C = CLBLM_L_X72Y130_SLICE_X108Y130_CO6;
  assign CLBLM_L_X72Y130_SLICE_X108Y130_D = CLBLM_L_X72Y130_SLICE_X108Y130_DO6;
  assign CLBLM_L_X72Y130_SLICE_X109Y130_A = CLBLM_L_X72Y130_SLICE_X109Y130_AO6;
  assign CLBLM_L_X72Y130_SLICE_X109Y130_B = CLBLM_L_X72Y130_SLICE_X109Y130_BO6;
  assign CLBLM_L_X72Y130_SLICE_X109Y130_C = CLBLM_L_X72Y130_SLICE_X109Y130_CO6;
  assign CLBLM_L_X72Y130_SLICE_X109Y130_D = CLBLM_L_X72Y130_SLICE_X109Y130_DO6;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_A = CLBLM_L_X72Y131_SLICE_X108Y131_AO6;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_B = CLBLM_L_X72Y131_SLICE_X108Y131_BO6;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_C = CLBLM_L_X72Y131_SLICE_X108Y131_CO6;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_D = CLBLM_L_X72Y131_SLICE_X108Y131_DO6;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_AMUX = CLBLM_L_X72Y131_SLICE_X108Y131_A5Q;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_DMUX = CLBLM_L_X72Y131_SLICE_X108Y131_DO5;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_A = CLBLM_L_X72Y131_SLICE_X109Y131_AO6;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_B = CLBLM_L_X72Y131_SLICE_X109Y131_BO6;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_C = CLBLM_L_X72Y131_SLICE_X109Y131_CO6;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_D = CLBLM_L_X72Y131_SLICE_X109Y131_DO6;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_AMUX = CLBLM_L_X72Y131_SLICE_X109Y131_AO5;
  assign CLBLM_L_X72Y132_SLICE_X108Y132_A = CLBLM_L_X72Y132_SLICE_X108Y132_AO6;
  assign CLBLM_L_X72Y132_SLICE_X108Y132_B = CLBLM_L_X72Y132_SLICE_X108Y132_BO6;
  assign CLBLM_L_X72Y132_SLICE_X108Y132_C = CLBLM_L_X72Y132_SLICE_X108Y132_CO6;
  assign CLBLM_L_X72Y132_SLICE_X108Y132_D = CLBLM_L_X72Y132_SLICE_X108Y132_DO6;
  assign CLBLM_L_X72Y132_SLICE_X109Y132_A = CLBLM_L_X72Y132_SLICE_X109Y132_AO6;
  assign CLBLM_L_X72Y132_SLICE_X109Y132_B = CLBLM_L_X72Y132_SLICE_X109Y132_BO6;
  assign CLBLM_L_X72Y132_SLICE_X109Y132_C = CLBLM_L_X72Y132_SLICE_X109Y132_CO6;
  assign CLBLM_L_X72Y132_SLICE_X109Y132_D = CLBLM_L_X72Y132_SLICE_X109Y132_DO6;
  assign CLBLM_L_X72Y132_SLICE_X109Y132_CMUX = CLBLM_L_X72Y132_SLICE_X109Y132_CO6;
  assign CLBLM_L_X72Y133_SLICE_X108Y133_A = CLBLM_L_X72Y133_SLICE_X108Y133_AO6;
  assign CLBLM_L_X72Y133_SLICE_X108Y133_B = CLBLM_L_X72Y133_SLICE_X108Y133_BO6;
  assign CLBLM_L_X72Y133_SLICE_X108Y133_C = CLBLM_L_X72Y133_SLICE_X108Y133_CO6;
  assign CLBLM_L_X72Y133_SLICE_X108Y133_D = CLBLM_L_X72Y133_SLICE_X108Y133_DO6;
  assign CLBLM_L_X72Y133_SLICE_X108Y133_AMUX = CLBLM_L_X72Y133_SLICE_X108Y133_A5Q;
  assign CLBLM_L_X72Y133_SLICE_X108Y133_BMUX = CLBLM_L_X72Y133_SLICE_X108Y133_BO5;
  assign CLBLM_L_X72Y133_SLICE_X108Y133_DMUX = CLBLM_L_X72Y133_SLICE_X108Y133_DO5;
  assign CLBLM_L_X72Y133_SLICE_X109Y133_A = CLBLM_L_X72Y133_SLICE_X109Y133_AO6;
  assign CLBLM_L_X72Y133_SLICE_X109Y133_B = CLBLM_L_X72Y133_SLICE_X109Y133_BO6;
  assign CLBLM_L_X72Y133_SLICE_X109Y133_C = CLBLM_L_X72Y133_SLICE_X109Y133_CO6;
  assign CLBLM_L_X72Y133_SLICE_X109Y133_D = CLBLM_L_X72Y133_SLICE_X109Y133_DO6;
  assign CLBLM_L_X72Y133_SLICE_X109Y133_AMUX = CLBLM_L_X72Y133_SLICE_X109Y133_AO5;
  assign CLBLM_L_X72Y134_SLICE_X108Y134_A = CLBLM_L_X72Y134_SLICE_X108Y134_AO6;
  assign CLBLM_L_X72Y134_SLICE_X108Y134_B = CLBLM_L_X72Y134_SLICE_X108Y134_BO6;
  assign CLBLM_L_X72Y134_SLICE_X108Y134_C = CLBLM_L_X72Y134_SLICE_X108Y134_CO6;
  assign CLBLM_L_X72Y134_SLICE_X108Y134_D = CLBLM_L_X72Y134_SLICE_X108Y134_DO6;
  assign CLBLM_L_X72Y134_SLICE_X109Y134_A = CLBLM_L_X72Y134_SLICE_X109Y134_AO6;
  assign CLBLM_L_X72Y134_SLICE_X109Y134_B = CLBLM_L_X72Y134_SLICE_X109Y134_BO6;
  assign CLBLM_L_X72Y134_SLICE_X109Y134_C = CLBLM_L_X72Y134_SLICE_X109Y134_CO6;
  assign CLBLM_L_X72Y134_SLICE_X109Y134_D = CLBLM_L_X72Y134_SLICE_X109Y134_DO6;
  assign CLBLM_L_X72Y134_SLICE_X109Y134_AMUX = CLBLM_L_X72Y134_SLICE_X109Y134_AO5;
  assign CLBLM_L_X72Y134_SLICE_X109Y134_BMUX = CLBLM_L_X72Y134_SLICE_X109Y134_BO5;
  assign CLBLM_L_X74Y102_SLICE_X112Y102_A = CLBLM_L_X74Y102_SLICE_X112Y102_AO6;
  assign CLBLM_L_X74Y102_SLICE_X112Y102_B = CLBLM_L_X74Y102_SLICE_X112Y102_BO6;
  assign CLBLM_L_X74Y102_SLICE_X112Y102_C = CLBLM_L_X74Y102_SLICE_X112Y102_CO6;
  assign CLBLM_L_X74Y102_SLICE_X112Y102_D = CLBLM_L_X74Y102_SLICE_X112Y102_DO6;
  assign CLBLM_L_X74Y102_SLICE_X113Y102_A = CLBLM_L_X74Y102_SLICE_X113Y102_AO6;
  assign CLBLM_L_X74Y102_SLICE_X113Y102_B = CLBLM_L_X74Y102_SLICE_X113Y102_BO6;
  assign CLBLM_L_X74Y102_SLICE_X113Y102_C = CLBLM_L_X74Y102_SLICE_X113Y102_CO6;
  assign CLBLM_L_X74Y102_SLICE_X113Y102_D = CLBLM_L_X74Y102_SLICE_X113Y102_DO6;
  assign CLBLM_L_X74Y103_SLICE_X112Y103_A = CLBLM_L_X74Y103_SLICE_X112Y103_AO6;
  assign CLBLM_L_X74Y103_SLICE_X112Y103_B = CLBLM_L_X74Y103_SLICE_X112Y103_BO6;
  assign CLBLM_L_X74Y103_SLICE_X112Y103_C = CLBLM_L_X74Y103_SLICE_X112Y103_CO6;
  assign CLBLM_L_X74Y103_SLICE_X112Y103_D = CLBLM_L_X74Y103_SLICE_X112Y103_DO6;
  assign CLBLM_L_X74Y103_SLICE_X112Y103_DMUX = CLBLM_L_X74Y103_SLICE_X112Y103_DO6;
  assign CLBLM_L_X74Y103_SLICE_X113Y103_A = CLBLM_L_X74Y103_SLICE_X113Y103_AO6;
  assign CLBLM_L_X74Y103_SLICE_X113Y103_B = CLBLM_L_X74Y103_SLICE_X113Y103_BO6;
  assign CLBLM_L_X74Y103_SLICE_X113Y103_C = CLBLM_L_X74Y103_SLICE_X113Y103_CO6;
  assign CLBLM_L_X74Y103_SLICE_X113Y103_D = CLBLM_L_X74Y103_SLICE_X113Y103_DO6;
  assign CLBLM_L_X74Y104_SLICE_X112Y104_A = CLBLM_L_X74Y104_SLICE_X112Y104_AO6;
  assign CLBLM_L_X74Y104_SLICE_X112Y104_B = CLBLM_L_X74Y104_SLICE_X112Y104_BO6;
  assign CLBLM_L_X74Y104_SLICE_X112Y104_C = CLBLM_L_X74Y104_SLICE_X112Y104_CO6;
  assign CLBLM_L_X74Y104_SLICE_X112Y104_D = CLBLM_L_X74Y104_SLICE_X112Y104_DO6;
  assign CLBLM_L_X74Y104_SLICE_X113Y104_A = CLBLM_L_X74Y104_SLICE_X113Y104_AO6;
  assign CLBLM_L_X74Y104_SLICE_X113Y104_B = CLBLM_L_X74Y104_SLICE_X113Y104_BO6;
  assign CLBLM_L_X74Y104_SLICE_X113Y104_C = CLBLM_L_X74Y104_SLICE_X113Y104_CO6;
  assign CLBLM_L_X74Y104_SLICE_X113Y104_D = CLBLM_L_X74Y104_SLICE_X113Y104_DO6;
  assign CLBLM_L_X74Y107_SLICE_X112Y107_A = CLBLM_L_X74Y107_SLICE_X112Y107_AO6;
  assign CLBLM_L_X74Y107_SLICE_X112Y107_B = CLBLM_L_X74Y107_SLICE_X112Y107_BO6;
  assign CLBLM_L_X74Y107_SLICE_X112Y107_C = CLBLM_L_X74Y107_SLICE_X112Y107_CO6;
  assign CLBLM_L_X74Y107_SLICE_X112Y107_D = CLBLM_L_X74Y107_SLICE_X112Y107_DO6;
  assign CLBLM_L_X74Y107_SLICE_X113Y107_A = CLBLM_L_X74Y107_SLICE_X113Y107_AO6;
  assign CLBLM_L_X74Y107_SLICE_X113Y107_B = CLBLM_L_X74Y107_SLICE_X113Y107_BO6;
  assign CLBLM_L_X74Y107_SLICE_X113Y107_C = CLBLM_L_X74Y107_SLICE_X113Y107_CO6;
  assign CLBLM_L_X74Y107_SLICE_X113Y107_D = CLBLM_L_X74Y107_SLICE_X113Y107_DO6;
  assign CLBLM_L_X74Y109_SLICE_X112Y109_A = CLBLM_L_X74Y109_SLICE_X112Y109_AO6;
  assign CLBLM_L_X74Y109_SLICE_X112Y109_B = CLBLM_L_X74Y109_SLICE_X112Y109_BO6;
  assign CLBLM_L_X74Y109_SLICE_X112Y109_C = CLBLM_L_X74Y109_SLICE_X112Y109_CO6;
  assign CLBLM_L_X74Y109_SLICE_X112Y109_D = CLBLM_L_X74Y109_SLICE_X112Y109_DO6;
  assign CLBLM_L_X74Y109_SLICE_X113Y109_A = CLBLM_L_X74Y109_SLICE_X113Y109_AO6;
  assign CLBLM_L_X74Y109_SLICE_X113Y109_B = CLBLM_L_X74Y109_SLICE_X113Y109_BO6;
  assign CLBLM_L_X74Y109_SLICE_X113Y109_C = CLBLM_L_X74Y109_SLICE_X113Y109_CO6;
  assign CLBLM_L_X74Y109_SLICE_X113Y109_D = CLBLM_L_X74Y109_SLICE_X113Y109_DO6;
  assign CLBLM_L_X74Y109_SLICE_X113Y109_AMUX = CLBLM_L_X74Y109_SLICE_X113Y109_A5Q;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_A = CLBLM_L_X74Y117_SLICE_X112Y117_AO6;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_B = CLBLM_L_X74Y117_SLICE_X112Y117_BO6;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_C = CLBLM_L_X74Y117_SLICE_X112Y117_CO6;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_D = CLBLM_L_X74Y117_SLICE_X112Y117_DO6;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_A = CLBLM_L_X74Y117_SLICE_X113Y117_AO6;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_B = CLBLM_L_X74Y117_SLICE_X113Y117_BO6;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_C = CLBLM_L_X74Y117_SLICE_X113Y117_CO6;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_D = CLBLM_L_X74Y117_SLICE_X113Y117_DO6;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_A = CLBLM_L_X74Y118_SLICE_X112Y118_AO6;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_B = CLBLM_L_X74Y118_SLICE_X112Y118_BO6;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_C = CLBLM_L_X74Y118_SLICE_X112Y118_CO6;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_D = CLBLM_L_X74Y118_SLICE_X112Y118_DO6;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_BMUX = CLBLM_L_X74Y118_SLICE_X112Y118_BO5;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_A = CLBLM_L_X74Y118_SLICE_X113Y118_AO6;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_B = CLBLM_L_X74Y118_SLICE_X113Y118_BO6;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_C = CLBLM_L_X74Y118_SLICE_X113Y118_CO6;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_D = CLBLM_L_X74Y118_SLICE_X113Y118_DO6;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_A = CLBLM_L_X74Y119_SLICE_X112Y119_AO6;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_B = CLBLM_L_X74Y119_SLICE_X112Y119_BO6;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_C = CLBLM_L_X74Y119_SLICE_X112Y119_CO6;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_D = CLBLM_L_X74Y119_SLICE_X112Y119_DO6;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_BMUX = CLBLM_L_X74Y119_SLICE_X112Y119_BO5;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_A = CLBLM_L_X74Y119_SLICE_X113Y119_AO6;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_B = CLBLM_L_X74Y119_SLICE_X113Y119_BO6;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_C = CLBLM_L_X74Y119_SLICE_X113Y119_CO6;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_D = CLBLM_L_X74Y119_SLICE_X113Y119_DO6;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_AMUX = CLBLM_L_X74Y119_SLICE_X113Y119_AO6;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_A = CLBLM_L_X74Y120_SLICE_X112Y120_AO6;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_B = CLBLM_L_X74Y120_SLICE_X112Y120_BO6;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_C = CLBLM_L_X74Y120_SLICE_X112Y120_CO6;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_D = CLBLM_L_X74Y120_SLICE_X112Y120_DO6;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_A = CLBLM_L_X74Y120_SLICE_X113Y120_AO6;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_B = CLBLM_L_X74Y120_SLICE_X113Y120_BO6;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_C = CLBLM_L_X74Y120_SLICE_X113Y120_CO6;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_D = CLBLM_L_X74Y120_SLICE_X113Y120_DO6;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_A = CLBLM_L_X74Y121_SLICE_X112Y121_AO6;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_B = CLBLM_L_X74Y121_SLICE_X112Y121_BO6;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_C = CLBLM_L_X74Y121_SLICE_X112Y121_CO6;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_D = CLBLM_L_X74Y121_SLICE_X112Y121_DO6;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_A = CLBLM_L_X74Y121_SLICE_X113Y121_AO6;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_B = CLBLM_L_X74Y121_SLICE_X113Y121_BO6;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_C = CLBLM_L_X74Y121_SLICE_X113Y121_CO6;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_D = CLBLM_L_X74Y121_SLICE_X113Y121_DO6;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_AMUX = CLBLM_L_X74Y121_SLICE_X113Y121_A5Q;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_BMUX = CLBLM_L_X74Y121_SLICE_X113Y121_B5Q;
  assign CLBLM_L_X74Y122_SLICE_X112Y122_A = CLBLM_L_X74Y122_SLICE_X112Y122_AO6;
  assign CLBLM_L_X74Y122_SLICE_X112Y122_B = CLBLM_L_X74Y122_SLICE_X112Y122_BO6;
  assign CLBLM_L_X74Y122_SLICE_X112Y122_C = CLBLM_L_X74Y122_SLICE_X112Y122_CO6;
  assign CLBLM_L_X74Y122_SLICE_X112Y122_D = CLBLM_L_X74Y122_SLICE_X112Y122_DO6;
  assign CLBLM_L_X74Y122_SLICE_X112Y122_AMUX = CLBLM_L_X74Y122_SLICE_X112Y122_A5Q;
  assign CLBLM_L_X74Y122_SLICE_X113Y122_A = CLBLM_L_X74Y122_SLICE_X113Y122_AO6;
  assign CLBLM_L_X74Y122_SLICE_X113Y122_B = CLBLM_L_X74Y122_SLICE_X113Y122_BO6;
  assign CLBLM_L_X74Y122_SLICE_X113Y122_C = CLBLM_L_X74Y122_SLICE_X113Y122_CO6;
  assign CLBLM_L_X74Y122_SLICE_X113Y122_D = CLBLM_L_X74Y122_SLICE_X113Y122_DO6;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_A = CLBLM_L_X74Y123_SLICE_X112Y123_AO6;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_B = CLBLM_L_X74Y123_SLICE_X112Y123_BO6;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_C = CLBLM_L_X74Y123_SLICE_X112Y123_CO6;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_D = CLBLM_L_X74Y123_SLICE_X112Y123_DO6;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_BMUX = CLBLM_L_X74Y123_SLICE_X112Y123_B5Q;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_A = CLBLM_L_X74Y123_SLICE_X113Y123_AO6;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_B = CLBLM_L_X74Y123_SLICE_X113Y123_BO6;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_C = CLBLM_L_X74Y123_SLICE_X113Y123_CO6;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_D = CLBLM_L_X74Y123_SLICE_X113Y123_DO6;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_AMUX = CLBLM_L_X74Y123_SLICE_X113Y123_A5Q;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_CMUX = CLBLM_L_X74Y123_SLICE_X113Y123_CO5;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_A = CLBLM_L_X74Y125_SLICE_X112Y125_AO6;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_B = CLBLM_L_X74Y125_SLICE_X112Y125_BO6;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_C = CLBLM_L_X74Y125_SLICE_X112Y125_CO6;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_D = CLBLM_L_X74Y125_SLICE_X112Y125_DO6;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_A = CLBLM_L_X74Y125_SLICE_X113Y125_AO6;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_B = CLBLM_L_X74Y125_SLICE_X113Y125_BO6;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_C = CLBLM_L_X74Y125_SLICE_X113Y125_CO6;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_D = CLBLM_L_X74Y125_SLICE_X113Y125_DO6;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_A = CLBLM_L_X74Y126_SLICE_X112Y126_AO6;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_B = CLBLM_L_X74Y126_SLICE_X112Y126_BO6;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_C = CLBLM_L_X74Y126_SLICE_X112Y126_CO6;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_D = CLBLM_L_X74Y126_SLICE_X112Y126_DO6;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_AMUX = CLBLM_L_X74Y126_SLICE_X112Y126_A5Q;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_BMUX = CLBLM_L_X74Y126_SLICE_X112Y126_BO5;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_CMUX = CLBLM_L_X74Y126_SLICE_X112Y126_CO5;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_A = CLBLM_L_X74Y126_SLICE_X113Y126_AO6;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_B = CLBLM_L_X74Y126_SLICE_X113Y126_BO6;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_C = CLBLM_L_X74Y126_SLICE_X113Y126_CO6;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_D = CLBLM_L_X74Y126_SLICE_X113Y126_DO6;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_AMUX = CLBLM_L_X74Y126_SLICE_X113Y126_A5Q;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_A = CLBLM_L_X74Y127_SLICE_X112Y127_AO6;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_B = CLBLM_L_X74Y127_SLICE_X112Y127_BO6;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_C = CLBLM_L_X74Y127_SLICE_X112Y127_CO6;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_D = CLBLM_L_X74Y127_SLICE_X112Y127_DO6;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_AMUX = CLBLM_L_X74Y127_SLICE_X112Y127_AO5;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_CMUX = CLBLM_L_X74Y127_SLICE_X112Y127_CO6;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_A = CLBLM_L_X74Y127_SLICE_X113Y127_AO6;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_B = CLBLM_L_X74Y127_SLICE_X113Y127_BO6;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_C = CLBLM_L_X74Y127_SLICE_X113Y127_CO6;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_D = CLBLM_L_X74Y127_SLICE_X113Y127_DO6;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_AMUX = CLBLM_L_X74Y127_SLICE_X113Y127_A5Q;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_BMUX = CLBLM_L_X74Y127_SLICE_X113Y127_BO5;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_A = CLBLM_L_X74Y128_SLICE_X112Y128_AO6;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_B = CLBLM_L_X74Y128_SLICE_X112Y128_BO6;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_C = CLBLM_L_X74Y128_SLICE_X112Y128_CO6;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_D = CLBLM_L_X74Y128_SLICE_X112Y128_DO6;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_A = CLBLM_L_X74Y128_SLICE_X113Y128_AO6;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_B = CLBLM_L_X74Y128_SLICE_X113Y128_BO6;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_C = CLBLM_L_X74Y128_SLICE_X113Y128_CO6;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_D = CLBLM_L_X74Y128_SLICE_X113Y128_DO6;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_AMUX = CLBLM_L_X74Y128_SLICE_X113Y128_AO5;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_BMUX = CLBLM_L_X74Y128_SLICE_X113Y128_BO5;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_A = CLBLM_L_X74Y129_SLICE_X112Y129_AO6;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_B = CLBLM_L_X74Y129_SLICE_X112Y129_BO6;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_C = CLBLM_L_X74Y129_SLICE_X112Y129_CO6;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_D = CLBLM_L_X74Y129_SLICE_X112Y129_DO6;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_AMUX = CLBLM_L_X74Y129_SLICE_X112Y129_A5Q;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_A = CLBLM_L_X74Y129_SLICE_X113Y129_AO6;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_B = CLBLM_L_X74Y129_SLICE_X113Y129_BO6;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_C = CLBLM_L_X74Y129_SLICE_X113Y129_CO6;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_D = CLBLM_L_X74Y129_SLICE_X113Y129_DO6;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_BMUX = CLBLM_L_X74Y129_SLICE_X113Y129_BO5;
  assign CLBLM_L_X74Y131_SLICE_X112Y131_A = CLBLM_L_X74Y131_SLICE_X112Y131_AO6;
  assign CLBLM_L_X74Y131_SLICE_X112Y131_B = CLBLM_L_X74Y131_SLICE_X112Y131_BO6;
  assign CLBLM_L_X74Y131_SLICE_X112Y131_C = CLBLM_L_X74Y131_SLICE_X112Y131_CO6;
  assign CLBLM_L_X74Y131_SLICE_X112Y131_D = CLBLM_L_X74Y131_SLICE_X112Y131_DO6;
  assign CLBLM_L_X74Y131_SLICE_X113Y131_A = CLBLM_L_X74Y131_SLICE_X113Y131_AO6;
  assign CLBLM_L_X74Y131_SLICE_X113Y131_B = CLBLM_L_X74Y131_SLICE_X113Y131_BO6;
  assign CLBLM_L_X74Y131_SLICE_X113Y131_C = CLBLM_L_X74Y131_SLICE_X113Y131_CO6;
  assign CLBLM_L_X74Y131_SLICE_X113Y131_D = CLBLM_L_X74Y131_SLICE_X113Y131_DO6;
  assign CLBLM_L_X74Y132_SLICE_X112Y132_A = CLBLM_L_X74Y132_SLICE_X112Y132_AO6;
  assign CLBLM_L_X74Y132_SLICE_X112Y132_B = CLBLM_L_X74Y132_SLICE_X112Y132_BO6;
  assign CLBLM_L_X74Y132_SLICE_X112Y132_C = CLBLM_L_X74Y132_SLICE_X112Y132_CO6;
  assign CLBLM_L_X74Y132_SLICE_X112Y132_D = CLBLM_L_X74Y132_SLICE_X112Y132_DO6;
  assign CLBLM_L_X74Y132_SLICE_X112Y132_AMUX = CLBLM_L_X74Y132_SLICE_X112Y132_A5Q;
  assign CLBLM_L_X74Y132_SLICE_X112Y132_BMUX = CLBLM_L_X74Y132_SLICE_X112Y132_BO5;
  assign CLBLM_L_X74Y132_SLICE_X112Y132_CMUX = CLBLM_L_X74Y132_SLICE_X112Y132_C5Q;
  assign CLBLM_L_X74Y132_SLICE_X113Y132_A = CLBLM_L_X74Y132_SLICE_X113Y132_AO6;
  assign CLBLM_L_X74Y132_SLICE_X113Y132_B = CLBLM_L_X74Y132_SLICE_X113Y132_BO6;
  assign CLBLM_L_X74Y132_SLICE_X113Y132_C = CLBLM_L_X74Y132_SLICE_X113Y132_CO6;
  assign CLBLM_L_X74Y132_SLICE_X113Y132_D = CLBLM_L_X74Y132_SLICE_X113Y132_DO6;
  assign CLBLM_L_X74Y133_SLICE_X112Y133_A = CLBLM_L_X74Y133_SLICE_X112Y133_AO6;
  assign CLBLM_L_X74Y133_SLICE_X112Y133_B = CLBLM_L_X74Y133_SLICE_X112Y133_BO6;
  assign CLBLM_L_X74Y133_SLICE_X112Y133_C = CLBLM_L_X74Y133_SLICE_X112Y133_CO6;
  assign CLBLM_L_X74Y133_SLICE_X112Y133_D = CLBLM_L_X74Y133_SLICE_X112Y133_DO6;
  assign CLBLM_L_X74Y133_SLICE_X112Y133_DMUX = CLBLM_L_X74Y133_SLICE_X112Y133_DO5;
  assign CLBLM_L_X74Y133_SLICE_X113Y133_A = CLBLM_L_X74Y133_SLICE_X113Y133_AO6;
  assign CLBLM_L_X74Y133_SLICE_X113Y133_B = CLBLM_L_X74Y133_SLICE_X113Y133_BO6;
  assign CLBLM_L_X74Y133_SLICE_X113Y133_C = CLBLM_L_X74Y133_SLICE_X113Y133_CO6;
  assign CLBLM_L_X74Y133_SLICE_X113Y133_D = CLBLM_L_X74Y133_SLICE_X113Y133_DO6;
  assign CLBLM_L_X74Y133_SLICE_X113Y133_AMUX = CLBLM_L_X74Y133_SLICE_X113Y133_AO5;
  assign CLBLM_L_X74Y134_SLICE_X112Y134_A = CLBLM_L_X74Y134_SLICE_X112Y134_AO6;
  assign CLBLM_L_X74Y134_SLICE_X112Y134_B = CLBLM_L_X74Y134_SLICE_X112Y134_BO6;
  assign CLBLM_L_X74Y134_SLICE_X112Y134_C = CLBLM_L_X74Y134_SLICE_X112Y134_CO6;
  assign CLBLM_L_X74Y134_SLICE_X112Y134_D = CLBLM_L_X74Y134_SLICE_X112Y134_DO6;
  assign CLBLM_L_X74Y134_SLICE_X112Y134_AMUX = CLBLM_L_X74Y134_SLICE_X112Y134_AO5;
  assign CLBLM_L_X74Y134_SLICE_X113Y134_A = CLBLM_L_X74Y134_SLICE_X113Y134_AO6;
  assign CLBLM_L_X74Y134_SLICE_X113Y134_B = CLBLM_L_X74Y134_SLICE_X113Y134_BO6;
  assign CLBLM_L_X74Y134_SLICE_X113Y134_C = CLBLM_L_X74Y134_SLICE_X113Y134_CO6;
  assign CLBLM_L_X74Y134_SLICE_X113Y134_D = CLBLM_L_X74Y134_SLICE_X113Y134_DO6;
  assign CLBLM_L_X74Y134_SLICE_X113Y134_AMUX = CLBLM_L_X74Y134_SLICE_X113Y134_A5Q;
  assign CLBLM_L_X74Y134_SLICE_X113Y134_DMUX = CLBLM_L_X74Y134_SLICE_X113Y134_DO5;
  assign CLBLM_L_X74Y135_SLICE_X112Y135_A = CLBLM_L_X74Y135_SLICE_X112Y135_AO6;
  assign CLBLM_L_X74Y135_SLICE_X112Y135_B = CLBLM_L_X74Y135_SLICE_X112Y135_BO6;
  assign CLBLM_L_X74Y135_SLICE_X112Y135_C = CLBLM_L_X74Y135_SLICE_X112Y135_CO6;
  assign CLBLM_L_X74Y135_SLICE_X112Y135_D = CLBLM_L_X74Y135_SLICE_X112Y135_DO6;
  assign CLBLM_L_X74Y135_SLICE_X113Y135_A = CLBLM_L_X74Y135_SLICE_X113Y135_AO6;
  assign CLBLM_L_X74Y135_SLICE_X113Y135_B = CLBLM_L_X74Y135_SLICE_X113Y135_BO6;
  assign CLBLM_L_X74Y135_SLICE_X113Y135_C = CLBLM_L_X74Y135_SLICE_X113Y135_CO6;
  assign CLBLM_L_X74Y135_SLICE_X113Y135_D = CLBLM_L_X74Y135_SLICE_X113Y135_DO6;
  assign CLBLM_L_X76Y109_SLICE_X116Y109_A = CLBLM_L_X76Y109_SLICE_X116Y109_AO6;
  assign CLBLM_L_X76Y109_SLICE_X116Y109_B = CLBLM_L_X76Y109_SLICE_X116Y109_BO6;
  assign CLBLM_L_X76Y109_SLICE_X116Y109_C = CLBLM_L_X76Y109_SLICE_X116Y109_CO6;
  assign CLBLM_L_X76Y109_SLICE_X116Y109_D = CLBLM_L_X76Y109_SLICE_X116Y109_DO6;
  assign CLBLM_L_X76Y109_SLICE_X117Y109_A = CLBLM_L_X76Y109_SLICE_X117Y109_AO6;
  assign CLBLM_L_X76Y109_SLICE_X117Y109_B = CLBLM_L_X76Y109_SLICE_X117Y109_BO6;
  assign CLBLM_L_X76Y109_SLICE_X117Y109_C = CLBLM_L_X76Y109_SLICE_X117Y109_CO6;
  assign CLBLM_L_X76Y109_SLICE_X117Y109_D = CLBLM_L_X76Y109_SLICE_X117Y109_DO6;
  assign CLBLM_L_X76Y111_SLICE_X116Y111_A = CLBLM_L_X76Y111_SLICE_X116Y111_AO6;
  assign CLBLM_L_X76Y111_SLICE_X116Y111_B = CLBLM_L_X76Y111_SLICE_X116Y111_BO6;
  assign CLBLM_L_X76Y111_SLICE_X116Y111_C = CLBLM_L_X76Y111_SLICE_X116Y111_CO6;
  assign CLBLM_L_X76Y111_SLICE_X116Y111_D = CLBLM_L_X76Y111_SLICE_X116Y111_DO6;
  assign CLBLM_L_X76Y111_SLICE_X117Y111_A = CLBLM_L_X76Y111_SLICE_X117Y111_AO6;
  assign CLBLM_L_X76Y111_SLICE_X117Y111_B = CLBLM_L_X76Y111_SLICE_X117Y111_BO6;
  assign CLBLM_L_X76Y111_SLICE_X117Y111_C = CLBLM_L_X76Y111_SLICE_X117Y111_CO6;
  assign CLBLM_L_X76Y111_SLICE_X117Y111_D = CLBLM_L_X76Y111_SLICE_X117Y111_DO6;
  assign CLBLM_L_X76Y118_SLICE_X116Y118_A = CLBLM_L_X76Y118_SLICE_X116Y118_AO6;
  assign CLBLM_L_X76Y118_SLICE_X116Y118_B = CLBLM_L_X76Y118_SLICE_X116Y118_BO6;
  assign CLBLM_L_X76Y118_SLICE_X116Y118_C = CLBLM_L_X76Y118_SLICE_X116Y118_CO6;
  assign CLBLM_L_X76Y118_SLICE_X116Y118_D = CLBLM_L_X76Y118_SLICE_X116Y118_DO6;
  assign CLBLM_L_X76Y118_SLICE_X116Y118_AMUX = CLBLM_L_X76Y118_SLICE_X116Y118_A5Q;
  assign CLBLM_L_X76Y118_SLICE_X117Y118_A = CLBLM_L_X76Y118_SLICE_X117Y118_AO6;
  assign CLBLM_L_X76Y118_SLICE_X117Y118_B = CLBLM_L_X76Y118_SLICE_X117Y118_BO6;
  assign CLBLM_L_X76Y118_SLICE_X117Y118_C = CLBLM_L_X76Y118_SLICE_X117Y118_CO6;
  assign CLBLM_L_X76Y118_SLICE_X117Y118_D = CLBLM_L_X76Y118_SLICE_X117Y118_DO6;
  assign CLBLM_L_X76Y119_SLICE_X116Y119_A = CLBLM_L_X76Y119_SLICE_X116Y119_AO6;
  assign CLBLM_L_X76Y119_SLICE_X116Y119_B = CLBLM_L_X76Y119_SLICE_X116Y119_BO6;
  assign CLBLM_L_X76Y119_SLICE_X116Y119_C = CLBLM_L_X76Y119_SLICE_X116Y119_CO6;
  assign CLBLM_L_X76Y119_SLICE_X116Y119_D = CLBLM_L_X76Y119_SLICE_X116Y119_DO6;
  assign CLBLM_L_X76Y119_SLICE_X116Y119_AMUX = CLBLM_L_X76Y119_SLICE_X116Y119_A5Q;
  assign CLBLM_L_X76Y119_SLICE_X117Y119_A = CLBLM_L_X76Y119_SLICE_X117Y119_AO6;
  assign CLBLM_L_X76Y119_SLICE_X117Y119_B = CLBLM_L_X76Y119_SLICE_X117Y119_BO6;
  assign CLBLM_L_X76Y119_SLICE_X117Y119_C = CLBLM_L_X76Y119_SLICE_X117Y119_CO6;
  assign CLBLM_L_X76Y119_SLICE_X117Y119_D = CLBLM_L_X76Y119_SLICE_X117Y119_DO6;
  assign CLBLM_L_X76Y122_SLICE_X116Y122_A = CLBLM_L_X76Y122_SLICE_X116Y122_AO6;
  assign CLBLM_L_X76Y122_SLICE_X116Y122_B = CLBLM_L_X76Y122_SLICE_X116Y122_BO6;
  assign CLBLM_L_X76Y122_SLICE_X116Y122_C = CLBLM_L_X76Y122_SLICE_X116Y122_CO6;
  assign CLBLM_L_X76Y122_SLICE_X116Y122_D = CLBLM_L_X76Y122_SLICE_X116Y122_DO6;
  assign CLBLM_L_X76Y122_SLICE_X116Y122_AMUX = CLBLM_L_X76Y122_SLICE_X116Y122_A5Q;
  assign CLBLM_L_X76Y122_SLICE_X116Y122_CMUX = CLBLM_L_X76Y122_SLICE_X116Y122_C5Q;
  assign CLBLM_L_X76Y122_SLICE_X117Y122_A = CLBLM_L_X76Y122_SLICE_X117Y122_AO6;
  assign CLBLM_L_X76Y122_SLICE_X117Y122_B = CLBLM_L_X76Y122_SLICE_X117Y122_BO6;
  assign CLBLM_L_X76Y122_SLICE_X117Y122_C = CLBLM_L_X76Y122_SLICE_X117Y122_CO6;
  assign CLBLM_L_X76Y122_SLICE_X117Y122_D = CLBLM_L_X76Y122_SLICE_X117Y122_DO6;
  assign CLBLM_L_X76Y123_SLICE_X116Y123_A = CLBLM_L_X76Y123_SLICE_X116Y123_AO6;
  assign CLBLM_L_X76Y123_SLICE_X116Y123_B = CLBLM_L_X76Y123_SLICE_X116Y123_BO6;
  assign CLBLM_L_X76Y123_SLICE_X116Y123_C = CLBLM_L_X76Y123_SLICE_X116Y123_CO6;
  assign CLBLM_L_X76Y123_SLICE_X116Y123_D = CLBLM_L_X76Y123_SLICE_X116Y123_DO6;
  assign CLBLM_L_X76Y123_SLICE_X116Y123_AMUX = CLBLM_L_X76Y123_SLICE_X116Y123_A5Q;
  assign CLBLM_L_X76Y123_SLICE_X117Y123_A = CLBLM_L_X76Y123_SLICE_X117Y123_AO6;
  assign CLBLM_L_X76Y123_SLICE_X117Y123_B = CLBLM_L_X76Y123_SLICE_X117Y123_BO6;
  assign CLBLM_L_X76Y123_SLICE_X117Y123_C = CLBLM_L_X76Y123_SLICE_X117Y123_CO6;
  assign CLBLM_L_X76Y123_SLICE_X117Y123_D = CLBLM_L_X76Y123_SLICE_X117Y123_DO6;
  assign CLBLM_L_X76Y123_SLICE_X117Y123_AMUX = CLBLM_L_X76Y123_SLICE_X117Y123_AO5;
  assign CLBLM_L_X76Y123_SLICE_X117Y123_BMUX = CLBLM_L_X76Y123_SLICE_X117Y123_B5Q;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_A = CLBLM_L_X76Y124_SLICE_X116Y124_AO6;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_B = CLBLM_L_X76Y124_SLICE_X116Y124_BO6;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_C = CLBLM_L_X76Y124_SLICE_X116Y124_CO6;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_D = CLBLM_L_X76Y124_SLICE_X116Y124_DO6;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_AMUX = CLBLM_L_X76Y124_SLICE_X116Y124_A5Q;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_BMUX = CLBLM_L_X76Y124_SLICE_X116Y124_B5Q;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_A = CLBLM_L_X76Y124_SLICE_X117Y124_AO6;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_B = CLBLM_L_X76Y124_SLICE_X117Y124_BO6;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_C = CLBLM_L_X76Y124_SLICE_X117Y124_CO6;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_D = CLBLM_L_X76Y124_SLICE_X117Y124_DO6;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_A = CLBLM_L_X76Y125_SLICE_X116Y125_AO6;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_B = CLBLM_L_X76Y125_SLICE_X116Y125_BO6;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_C = CLBLM_L_X76Y125_SLICE_X116Y125_CO6;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_D = CLBLM_L_X76Y125_SLICE_X116Y125_DO6;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_AMUX = CLBLM_L_X76Y125_SLICE_X116Y125_A5Q;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_CMUX = CLBLM_L_X76Y125_SLICE_X116Y125_C5Q;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_A = CLBLM_L_X76Y125_SLICE_X117Y125_AO6;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_B = CLBLM_L_X76Y125_SLICE_X117Y125_BO6;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_C = CLBLM_L_X76Y125_SLICE_X117Y125_CO6;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_D = CLBLM_L_X76Y125_SLICE_X117Y125_DO6;
  assign CLBLM_L_X76Y126_SLICE_X116Y126_A = CLBLM_L_X76Y126_SLICE_X116Y126_AO6;
  assign CLBLM_L_X76Y126_SLICE_X116Y126_B = CLBLM_L_X76Y126_SLICE_X116Y126_BO6;
  assign CLBLM_L_X76Y126_SLICE_X116Y126_C = CLBLM_L_X76Y126_SLICE_X116Y126_CO6;
  assign CLBLM_L_X76Y126_SLICE_X116Y126_D = CLBLM_L_X76Y126_SLICE_X116Y126_DO6;
  assign CLBLM_L_X76Y126_SLICE_X116Y126_AMUX = CLBLM_L_X76Y126_SLICE_X116Y126_AO5;
  assign CLBLM_L_X76Y126_SLICE_X116Y126_BMUX = CLBLM_L_X76Y126_SLICE_X116Y126_B5Q;
  assign CLBLM_L_X76Y126_SLICE_X117Y126_A = CLBLM_L_X76Y126_SLICE_X117Y126_AO6;
  assign CLBLM_L_X76Y126_SLICE_X117Y126_B = CLBLM_L_X76Y126_SLICE_X117Y126_BO6;
  assign CLBLM_L_X76Y126_SLICE_X117Y126_C = CLBLM_L_X76Y126_SLICE_X117Y126_CO6;
  assign CLBLM_L_X76Y126_SLICE_X117Y126_D = CLBLM_L_X76Y126_SLICE_X117Y126_DO6;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_A = CLBLM_L_X76Y127_SLICE_X116Y127_AO6;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_B = CLBLM_L_X76Y127_SLICE_X116Y127_BO6;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_C = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_D = CLBLM_L_X76Y127_SLICE_X116Y127_DO6;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_A = CLBLM_L_X76Y127_SLICE_X117Y127_AO6;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_B = CLBLM_L_X76Y127_SLICE_X117Y127_BO6;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_C = CLBLM_L_X76Y127_SLICE_X117Y127_CO6;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_D = CLBLM_L_X76Y127_SLICE_X117Y127_DO6;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_A = CLBLM_L_X76Y128_SLICE_X116Y128_AO6;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_B = CLBLM_L_X76Y128_SLICE_X116Y128_BO6;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_C = CLBLM_L_X76Y128_SLICE_X116Y128_CO6;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_D = CLBLM_L_X76Y128_SLICE_X116Y128_DO6;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_AMUX = CLBLM_L_X76Y128_SLICE_X116Y128_A5Q;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_CMUX = CLBLM_L_X76Y128_SLICE_X116Y128_C5Q;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_A = CLBLM_L_X76Y128_SLICE_X117Y128_AO6;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_B = CLBLM_L_X76Y128_SLICE_X117Y128_BO6;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_C = CLBLM_L_X76Y128_SLICE_X117Y128_CO6;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_D = CLBLM_L_X76Y128_SLICE_X117Y128_DO6;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_AMUX = CLBLM_L_X76Y128_SLICE_X117Y128_A5Q;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_BMUX = CLBLM_L_X76Y128_SLICE_X117Y128_B5Q;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_CMUX = CLBLM_L_X76Y128_SLICE_X117Y128_CO5;
  assign CLBLM_L_X76Y129_SLICE_X116Y129_A = CLBLM_L_X76Y129_SLICE_X116Y129_AO6;
  assign CLBLM_L_X76Y129_SLICE_X116Y129_B = CLBLM_L_X76Y129_SLICE_X116Y129_BO6;
  assign CLBLM_L_X76Y129_SLICE_X116Y129_C = CLBLM_L_X76Y129_SLICE_X116Y129_CO6;
  assign CLBLM_L_X76Y129_SLICE_X116Y129_D = CLBLM_L_X76Y129_SLICE_X116Y129_DO6;
  assign CLBLM_L_X76Y129_SLICE_X116Y129_AMUX = CLBLM_L_X76Y129_SLICE_X116Y129_AO5;
  assign CLBLM_L_X76Y129_SLICE_X116Y129_BMUX = CLBLM_L_X76Y129_SLICE_X116Y129_B5Q;
  assign CLBLM_L_X76Y129_SLICE_X116Y129_DMUX = CLBLM_L_X76Y129_SLICE_X116Y129_DO6;
  assign CLBLM_L_X76Y129_SLICE_X117Y129_A = CLBLM_L_X76Y129_SLICE_X117Y129_AO6;
  assign CLBLM_L_X76Y129_SLICE_X117Y129_B = CLBLM_L_X76Y129_SLICE_X117Y129_BO6;
  assign CLBLM_L_X76Y129_SLICE_X117Y129_C = CLBLM_L_X76Y129_SLICE_X117Y129_CO6;
  assign CLBLM_L_X76Y129_SLICE_X117Y129_D = CLBLM_L_X76Y129_SLICE_X117Y129_DO6;
  assign CLBLM_L_X76Y130_SLICE_X116Y130_A = CLBLM_L_X76Y130_SLICE_X116Y130_AO6;
  assign CLBLM_L_X76Y130_SLICE_X116Y130_B = CLBLM_L_X76Y130_SLICE_X116Y130_BO6;
  assign CLBLM_L_X76Y130_SLICE_X116Y130_C = CLBLM_L_X76Y130_SLICE_X116Y130_CO6;
  assign CLBLM_L_X76Y130_SLICE_X116Y130_D = CLBLM_L_X76Y130_SLICE_X116Y130_DO6;
  assign CLBLM_L_X76Y130_SLICE_X116Y130_AMUX = CLBLM_L_X76Y130_SLICE_X116Y130_A5Q;
  assign CLBLM_L_X76Y130_SLICE_X116Y130_CMUX = CLBLM_L_X76Y130_SLICE_X116Y130_CO5;
  assign CLBLM_L_X76Y130_SLICE_X117Y130_A = CLBLM_L_X76Y130_SLICE_X117Y130_AO6;
  assign CLBLM_L_X76Y130_SLICE_X117Y130_B = CLBLM_L_X76Y130_SLICE_X117Y130_BO6;
  assign CLBLM_L_X76Y130_SLICE_X117Y130_C = CLBLM_L_X76Y130_SLICE_X117Y130_CO6;
  assign CLBLM_L_X76Y130_SLICE_X117Y130_D = CLBLM_L_X76Y130_SLICE_X117Y130_DO6;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_A = CLBLM_L_X76Y133_SLICE_X116Y133_AO6;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_B = CLBLM_L_X76Y133_SLICE_X116Y133_BO6;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_C = CLBLM_L_X76Y133_SLICE_X116Y133_CO6;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_D = CLBLM_L_X76Y133_SLICE_X116Y133_DO6;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_A = CLBLM_L_X76Y133_SLICE_X117Y133_AO6;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_B = CLBLM_L_X76Y133_SLICE_X117Y133_BO6;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_C = CLBLM_L_X76Y133_SLICE_X117Y133_CO6;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_D = CLBLM_L_X76Y133_SLICE_X117Y133_DO6;
  assign CLBLM_L_X76Y134_SLICE_X116Y134_A = CLBLM_L_X76Y134_SLICE_X116Y134_AO6;
  assign CLBLM_L_X76Y134_SLICE_X116Y134_B = CLBLM_L_X76Y134_SLICE_X116Y134_BO6;
  assign CLBLM_L_X76Y134_SLICE_X116Y134_C = CLBLM_L_X76Y134_SLICE_X116Y134_CO6;
  assign CLBLM_L_X76Y134_SLICE_X116Y134_D = CLBLM_L_X76Y134_SLICE_X116Y134_DO6;
  assign CLBLM_L_X76Y134_SLICE_X117Y134_A = CLBLM_L_X76Y134_SLICE_X117Y134_AO6;
  assign CLBLM_L_X76Y134_SLICE_X117Y134_B = CLBLM_L_X76Y134_SLICE_X117Y134_BO6;
  assign CLBLM_L_X76Y134_SLICE_X117Y134_C = CLBLM_L_X76Y134_SLICE_X117Y134_CO6;
  assign CLBLM_L_X76Y134_SLICE_X117Y134_D = CLBLM_L_X76Y134_SLICE_X117Y134_DO6;
  assign CLBLM_L_X76Y134_SLICE_X117Y134_CMUX = CLBLM_L_X76Y134_SLICE_X117Y134_CO6;
  assign CLBLM_L_X78Y104_SLICE_X120Y104_A = CLBLM_L_X78Y104_SLICE_X120Y104_AO6;
  assign CLBLM_L_X78Y104_SLICE_X120Y104_B = CLBLM_L_X78Y104_SLICE_X120Y104_BO6;
  assign CLBLM_L_X78Y104_SLICE_X120Y104_C = CLBLM_L_X78Y104_SLICE_X120Y104_CO6;
  assign CLBLM_L_X78Y104_SLICE_X120Y104_D = CLBLM_L_X78Y104_SLICE_X120Y104_DO6;
  assign CLBLM_L_X78Y104_SLICE_X120Y104_AMUX = CLBLM_L_X78Y104_SLICE_X120Y104_A5Q;
  assign CLBLM_L_X78Y104_SLICE_X121Y104_A = CLBLM_L_X78Y104_SLICE_X121Y104_AO6;
  assign CLBLM_L_X78Y104_SLICE_X121Y104_B = CLBLM_L_X78Y104_SLICE_X121Y104_BO6;
  assign CLBLM_L_X78Y104_SLICE_X121Y104_C = CLBLM_L_X78Y104_SLICE_X121Y104_CO6;
  assign CLBLM_L_X78Y104_SLICE_X121Y104_D = CLBLM_L_X78Y104_SLICE_X121Y104_DO6;
  assign CLBLM_L_X78Y106_SLICE_X120Y106_A = CLBLM_L_X78Y106_SLICE_X120Y106_AO6;
  assign CLBLM_L_X78Y106_SLICE_X120Y106_B = CLBLM_L_X78Y106_SLICE_X120Y106_BO6;
  assign CLBLM_L_X78Y106_SLICE_X120Y106_C = CLBLM_L_X78Y106_SLICE_X120Y106_CO6;
  assign CLBLM_L_X78Y106_SLICE_X120Y106_D = CLBLM_L_X78Y106_SLICE_X120Y106_DO6;
  assign CLBLM_L_X78Y106_SLICE_X121Y106_A = CLBLM_L_X78Y106_SLICE_X121Y106_AO6;
  assign CLBLM_L_X78Y106_SLICE_X121Y106_B = CLBLM_L_X78Y106_SLICE_X121Y106_BO6;
  assign CLBLM_L_X78Y106_SLICE_X121Y106_C = CLBLM_L_X78Y106_SLICE_X121Y106_CO6;
  assign CLBLM_L_X78Y106_SLICE_X121Y106_D = CLBLM_L_X78Y106_SLICE_X121Y106_DO6;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_A = CLBLM_L_X78Y120_SLICE_X120Y120_AO6;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_B = CLBLM_L_X78Y120_SLICE_X120Y120_BO6;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_C = CLBLM_L_X78Y120_SLICE_X120Y120_CO6;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_D = CLBLM_L_X78Y120_SLICE_X120Y120_DO6;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_A = CLBLM_L_X78Y120_SLICE_X121Y120_AO6;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_B = CLBLM_L_X78Y120_SLICE_X121Y120_BO6;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_C = CLBLM_L_X78Y120_SLICE_X121Y120_CO6;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_D = CLBLM_L_X78Y120_SLICE_X121Y120_DO6;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_A = CLBLM_L_X78Y121_SLICE_X120Y121_AO6;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_B = CLBLM_L_X78Y121_SLICE_X120Y121_BO6;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_C = CLBLM_L_X78Y121_SLICE_X120Y121_CO6;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_D = CLBLM_L_X78Y121_SLICE_X120Y121_DO6;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_CMUX = CLBLM_L_X78Y121_SLICE_X120Y121_CO5;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_A = CLBLM_L_X78Y121_SLICE_X121Y121_AO6;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_B = CLBLM_L_X78Y121_SLICE_X121Y121_BO6;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_C = CLBLM_L_X78Y121_SLICE_X121Y121_CO6;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_D = CLBLM_L_X78Y121_SLICE_X121Y121_DO6;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_A = CLBLM_L_X78Y122_SLICE_X120Y122_AO6;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_B = CLBLM_L_X78Y122_SLICE_X120Y122_BO6;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_C = CLBLM_L_X78Y122_SLICE_X120Y122_CO6;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_D = CLBLM_L_X78Y122_SLICE_X120Y122_DO6;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_AMUX = CLBLM_L_X78Y122_SLICE_X120Y122_AO5;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_A = CLBLM_L_X78Y122_SLICE_X121Y122_AO6;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_B = CLBLM_L_X78Y122_SLICE_X121Y122_BO6;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_C = CLBLM_L_X78Y122_SLICE_X121Y122_CO6;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_D = CLBLM_L_X78Y122_SLICE_X121Y122_DO6;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_A = CLBLM_L_X78Y123_SLICE_X120Y123_AO6;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_B = CLBLM_L_X78Y123_SLICE_X120Y123_BO6;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_C = CLBLM_L_X78Y123_SLICE_X120Y123_CO6;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_D = CLBLM_L_X78Y123_SLICE_X120Y123_DO6;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_AMUX = CLBLM_L_X78Y123_SLICE_X120Y123_AO6;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_A = CLBLM_L_X78Y123_SLICE_X121Y123_AO6;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_B = CLBLM_L_X78Y123_SLICE_X121Y123_BO6;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_C = CLBLM_L_X78Y123_SLICE_X121Y123_CO6;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_D = CLBLM_L_X78Y123_SLICE_X121Y123_DO6;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_AMUX = CLBLM_L_X78Y123_SLICE_X121Y123_A5Q;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_CMUX = CLBLM_L_X78Y123_SLICE_X121Y123_CO5;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_A = CLBLM_L_X78Y124_SLICE_X120Y124_AO6;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_B = CLBLM_L_X78Y124_SLICE_X120Y124_BO6;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_C = CLBLM_L_X78Y124_SLICE_X120Y124_CO6;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_D = CLBLM_L_X78Y124_SLICE_X120Y124_DO6;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_A = CLBLM_L_X78Y124_SLICE_X121Y124_AO6;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_B = CLBLM_L_X78Y124_SLICE_X121Y124_BO6;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_C = CLBLM_L_X78Y124_SLICE_X121Y124_CO6;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_D = CLBLM_L_X78Y124_SLICE_X121Y124_DO6;
  assign CLBLM_L_X78Y127_SLICE_X120Y127_A = CLBLM_L_X78Y127_SLICE_X120Y127_AO6;
  assign CLBLM_L_X78Y127_SLICE_X120Y127_B = CLBLM_L_X78Y127_SLICE_X120Y127_BO6;
  assign CLBLM_L_X78Y127_SLICE_X120Y127_C = CLBLM_L_X78Y127_SLICE_X120Y127_CO6;
  assign CLBLM_L_X78Y127_SLICE_X120Y127_D = CLBLM_L_X78Y127_SLICE_X120Y127_DO6;
  assign CLBLM_L_X78Y127_SLICE_X121Y127_A = CLBLM_L_X78Y127_SLICE_X121Y127_AO6;
  assign CLBLM_L_X78Y127_SLICE_X121Y127_B = CLBLM_L_X78Y127_SLICE_X121Y127_BO6;
  assign CLBLM_L_X78Y127_SLICE_X121Y127_C = CLBLM_L_X78Y127_SLICE_X121Y127_CO6;
  assign CLBLM_L_X78Y127_SLICE_X121Y127_D = CLBLM_L_X78Y127_SLICE_X121Y127_DO6;
  assign CLBLM_L_X78Y127_SLICE_X121Y127_AMUX = CLBLM_L_X78Y127_SLICE_X121Y127_AO5;
  assign CLBLM_L_X78Y128_SLICE_X120Y128_A = CLBLM_L_X78Y128_SLICE_X120Y128_AO6;
  assign CLBLM_L_X78Y128_SLICE_X120Y128_B = CLBLM_L_X78Y128_SLICE_X120Y128_BO6;
  assign CLBLM_L_X78Y128_SLICE_X120Y128_C = CLBLM_L_X78Y128_SLICE_X120Y128_CO6;
  assign CLBLM_L_X78Y128_SLICE_X120Y128_D = CLBLM_L_X78Y128_SLICE_X120Y128_DO6;
  assign CLBLM_L_X78Y128_SLICE_X121Y128_A = CLBLM_L_X78Y128_SLICE_X121Y128_AO6;
  assign CLBLM_L_X78Y128_SLICE_X121Y128_B = CLBLM_L_X78Y128_SLICE_X121Y128_BO6;
  assign CLBLM_L_X78Y128_SLICE_X121Y128_C = CLBLM_L_X78Y128_SLICE_X121Y128_CO6;
  assign CLBLM_L_X78Y128_SLICE_X121Y128_D = CLBLM_L_X78Y128_SLICE_X121Y128_DO6;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_A = CLBLM_L_X78Y129_SLICE_X120Y129_AO6;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_B = CLBLM_L_X78Y129_SLICE_X120Y129_BO6;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_C = CLBLM_L_X78Y129_SLICE_X120Y129_CO6;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_D = CLBLM_L_X78Y129_SLICE_X120Y129_DO6;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_A = CLBLM_L_X78Y129_SLICE_X121Y129_AO6;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_B = CLBLM_L_X78Y129_SLICE_X121Y129_BO6;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_C = CLBLM_L_X78Y129_SLICE_X121Y129_CO6;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_D = CLBLM_L_X78Y129_SLICE_X121Y129_DO6;
  assign CLBLM_L_X78Y130_SLICE_X120Y130_A = CLBLM_L_X78Y130_SLICE_X120Y130_AO6;
  assign CLBLM_L_X78Y130_SLICE_X120Y130_B = CLBLM_L_X78Y130_SLICE_X120Y130_BO6;
  assign CLBLM_L_X78Y130_SLICE_X120Y130_C = CLBLM_L_X78Y130_SLICE_X120Y130_CO6;
  assign CLBLM_L_X78Y130_SLICE_X120Y130_D = CLBLM_L_X78Y130_SLICE_X120Y130_DO6;
  assign CLBLM_L_X78Y130_SLICE_X121Y130_A = CLBLM_L_X78Y130_SLICE_X121Y130_AO6;
  assign CLBLM_L_X78Y130_SLICE_X121Y130_B = CLBLM_L_X78Y130_SLICE_X121Y130_BO6;
  assign CLBLM_L_X78Y130_SLICE_X121Y130_C = CLBLM_L_X78Y130_SLICE_X121Y130_CO6;
  assign CLBLM_L_X78Y130_SLICE_X121Y130_D = CLBLM_L_X78Y130_SLICE_X121Y130_DO6;
  assign CLBLM_L_X78Y131_SLICE_X120Y131_A = CLBLM_L_X78Y131_SLICE_X120Y131_AO6;
  assign CLBLM_L_X78Y131_SLICE_X120Y131_B = CLBLM_L_X78Y131_SLICE_X120Y131_BO6;
  assign CLBLM_L_X78Y131_SLICE_X120Y131_C = CLBLM_L_X78Y131_SLICE_X120Y131_CO6;
  assign CLBLM_L_X78Y131_SLICE_X120Y131_D = CLBLM_L_X78Y131_SLICE_X120Y131_DO6;
  assign CLBLM_L_X78Y131_SLICE_X121Y131_A = CLBLM_L_X78Y131_SLICE_X121Y131_AO6;
  assign CLBLM_L_X78Y131_SLICE_X121Y131_B = CLBLM_L_X78Y131_SLICE_X121Y131_BO6;
  assign CLBLM_L_X78Y131_SLICE_X121Y131_C = CLBLM_L_X78Y131_SLICE_X121Y131_CO6;
  assign CLBLM_L_X78Y131_SLICE_X121Y131_D = CLBLM_L_X78Y131_SLICE_X121Y131_DO6;
  assign CLBLM_L_X80Y132_SLICE_X124Y132_A = CLBLM_L_X80Y132_SLICE_X124Y132_AO6;
  assign CLBLM_L_X80Y132_SLICE_X124Y132_B = CLBLM_L_X80Y132_SLICE_X124Y132_BO6;
  assign CLBLM_L_X80Y132_SLICE_X124Y132_C = CLBLM_L_X80Y132_SLICE_X124Y132_CO6;
  assign CLBLM_L_X80Y132_SLICE_X124Y132_D = CLBLM_L_X80Y132_SLICE_X124Y132_DO6;
  assign CLBLM_L_X80Y132_SLICE_X125Y132_A = CLBLM_L_X80Y132_SLICE_X125Y132_AO6;
  assign CLBLM_L_X80Y132_SLICE_X125Y132_B = CLBLM_L_X80Y132_SLICE_X125Y132_BO6;
  assign CLBLM_L_X80Y132_SLICE_X125Y132_C = CLBLM_L_X80Y132_SLICE_X125Y132_CO6;
  assign CLBLM_L_X80Y132_SLICE_X125Y132_D = CLBLM_L_X80Y132_SLICE_X125Y132_DO6;
  assign CLBLM_L_X82Y98_SLICE_X128Y98_A = CLBLM_L_X82Y98_SLICE_X128Y98_AO6;
  assign CLBLM_L_X82Y98_SLICE_X128Y98_B = CLBLM_L_X82Y98_SLICE_X128Y98_BO6;
  assign CLBLM_L_X82Y98_SLICE_X128Y98_C = CLBLM_L_X82Y98_SLICE_X128Y98_CO6;
  assign CLBLM_L_X82Y98_SLICE_X128Y98_D = CLBLM_L_X82Y98_SLICE_X128Y98_DO6;
  assign CLBLM_L_X82Y98_SLICE_X128Y98_AMUX = CLBLM_L_X82Y98_SLICE_X128Y98_A5Q;
  assign CLBLM_L_X82Y98_SLICE_X129Y98_A = CLBLM_L_X82Y98_SLICE_X129Y98_AO6;
  assign CLBLM_L_X82Y98_SLICE_X129Y98_B = CLBLM_L_X82Y98_SLICE_X129Y98_BO6;
  assign CLBLM_L_X82Y98_SLICE_X129Y98_C = CLBLM_L_X82Y98_SLICE_X129Y98_CO6;
  assign CLBLM_L_X82Y98_SLICE_X129Y98_D = CLBLM_L_X82Y98_SLICE_X129Y98_DO6;
  assign CLBLM_L_X82Y130_SLICE_X128Y130_A = CLBLM_L_X82Y130_SLICE_X128Y130_AO6;
  assign CLBLM_L_X82Y130_SLICE_X128Y130_B = CLBLM_L_X82Y130_SLICE_X128Y130_BO6;
  assign CLBLM_L_X82Y130_SLICE_X128Y130_C = CLBLM_L_X82Y130_SLICE_X128Y130_CO6;
  assign CLBLM_L_X82Y130_SLICE_X128Y130_D = CLBLM_L_X82Y130_SLICE_X128Y130_DO6;
  assign CLBLM_L_X82Y130_SLICE_X129Y130_A = CLBLM_L_X82Y130_SLICE_X129Y130_AO6;
  assign CLBLM_L_X82Y130_SLICE_X129Y130_B = CLBLM_L_X82Y130_SLICE_X129Y130_BO6;
  assign CLBLM_L_X82Y130_SLICE_X129Y130_C = CLBLM_L_X82Y130_SLICE_X129Y130_CO6;
  assign CLBLM_L_X82Y130_SLICE_X129Y130_D = CLBLM_L_X82Y130_SLICE_X129Y130_DO6;
  assign CLBLM_R_X53Y122_SLICE_X80Y122_A = CLBLM_R_X53Y122_SLICE_X80Y122_AO6;
  assign CLBLM_R_X53Y122_SLICE_X80Y122_B = CLBLM_R_X53Y122_SLICE_X80Y122_BO6;
  assign CLBLM_R_X53Y122_SLICE_X80Y122_C = CLBLM_R_X53Y122_SLICE_X80Y122_CO6;
  assign CLBLM_R_X53Y122_SLICE_X80Y122_D = CLBLM_R_X53Y122_SLICE_X80Y122_DO6;
  assign CLBLM_R_X53Y122_SLICE_X81Y122_A = CLBLM_R_X53Y122_SLICE_X81Y122_AO6;
  assign CLBLM_R_X53Y122_SLICE_X81Y122_B = CLBLM_R_X53Y122_SLICE_X81Y122_BO6;
  assign CLBLM_R_X53Y122_SLICE_X81Y122_C = CLBLM_R_X53Y122_SLICE_X81Y122_CO6;
  assign CLBLM_R_X53Y122_SLICE_X81Y122_D = CLBLM_R_X53Y122_SLICE_X81Y122_DO6;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_A = CLBLM_R_X63Y96_SLICE_X94Y96_AO6;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_B = CLBLM_R_X63Y96_SLICE_X94Y96_BO6;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_C = CLBLM_R_X63Y96_SLICE_X94Y96_CO6;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_D = CLBLM_R_X63Y96_SLICE_X94Y96_DO6;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_A = CLBLM_R_X63Y96_SLICE_X95Y96_AO6;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_B = CLBLM_R_X63Y96_SLICE_X95Y96_BO6;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_C = CLBLM_R_X63Y96_SLICE_X95Y96_CO6;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_D = CLBLM_R_X63Y96_SLICE_X95Y96_DO6;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_A = CLBLM_R_X63Y97_SLICE_X94Y97_AO6;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_B = CLBLM_R_X63Y97_SLICE_X94Y97_BO6;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_C = CLBLM_R_X63Y97_SLICE_X94Y97_CO6;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_D = CLBLM_R_X63Y97_SLICE_X94Y97_DO6;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_AMUX = CLBLM_R_X63Y97_SLICE_X94Y97_AO5;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_BMUX = CLBLM_R_X63Y97_SLICE_X94Y97_B5Q;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_A = CLBLM_R_X63Y97_SLICE_X95Y97_AO6;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_B = CLBLM_R_X63Y97_SLICE_X95Y97_BO6;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_C = CLBLM_R_X63Y97_SLICE_X95Y97_CO6;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_D = CLBLM_R_X63Y97_SLICE_X95Y97_DO6;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_BMUX = CLBLM_R_X63Y97_SLICE_X95Y97_BO6;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_A = CLBLM_R_X63Y98_SLICE_X94Y98_AO6;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_B = CLBLM_R_X63Y98_SLICE_X94Y98_BO6;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_C = CLBLM_R_X63Y98_SLICE_X94Y98_CO6;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_D = CLBLM_R_X63Y98_SLICE_X94Y98_DO6;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_AMUX = CLBLM_R_X63Y98_SLICE_X94Y98_AO5;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_BMUX = CLBLM_R_X63Y98_SLICE_X94Y98_BO5;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_CMUX = CLBLM_R_X63Y98_SLICE_X94Y98_CO6;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_DMUX = CLBLM_R_X63Y98_SLICE_X94Y98_DO6;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_A = CLBLM_R_X63Y98_SLICE_X95Y98_AO6;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_B = CLBLM_R_X63Y98_SLICE_X95Y98_BO6;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_C = CLBLM_R_X63Y98_SLICE_X95Y98_CO6;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_D = CLBLM_R_X63Y98_SLICE_X95Y98_DO6;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_A = CLBLM_R_X63Y99_SLICE_X94Y99_AO6;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_B = CLBLM_R_X63Y99_SLICE_X94Y99_BO6;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_C = CLBLM_R_X63Y99_SLICE_X94Y99_CO6;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_D = CLBLM_R_X63Y99_SLICE_X94Y99_DO6;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_AMUX = CLBLM_R_X63Y99_SLICE_X94Y99_A5Q;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_BMUX = CLBLM_R_X63Y99_SLICE_X94Y99_BO5;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_CMUX = CLBLM_R_X63Y99_SLICE_X94Y99_CO5;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_DMUX = CLBLM_R_X63Y99_SLICE_X94Y99_D5Q;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_A = CLBLM_R_X63Y99_SLICE_X95Y99_AO6;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_B = CLBLM_R_X63Y99_SLICE_X95Y99_BO6;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_C = CLBLM_R_X63Y99_SLICE_X95Y99_CO6;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_D = CLBLM_R_X63Y99_SLICE_X95Y99_DO6;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_AMUX = CLBLM_R_X63Y99_SLICE_X95Y99_AO5;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_BMUX = CLBLM_R_X63Y99_SLICE_X95Y99_B5Q;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_CMUX = CLBLM_R_X63Y99_SLICE_X95Y99_CO6;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_A = CLBLM_R_X63Y101_SLICE_X94Y101_AO6;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_B = CLBLM_R_X63Y101_SLICE_X94Y101_BO6;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_C = CLBLM_R_X63Y101_SLICE_X94Y101_CO6;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_D = CLBLM_R_X63Y101_SLICE_X94Y101_DO6;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_AMUX = CLBLM_R_X63Y101_SLICE_X94Y101_AO5;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_BMUX = CLBLM_R_X63Y101_SLICE_X94Y101_BO5;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_A = CLBLM_R_X63Y101_SLICE_X95Y101_AO6;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_B = CLBLM_R_X63Y101_SLICE_X95Y101_BO6;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_C = CLBLM_R_X63Y101_SLICE_X95Y101_CO6;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_D = CLBLM_R_X63Y101_SLICE_X95Y101_DO6;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_A = CLBLM_R_X63Y102_SLICE_X94Y102_AO6;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_B = CLBLM_R_X63Y102_SLICE_X94Y102_BO6;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_C = CLBLM_R_X63Y102_SLICE_X94Y102_CO6;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_D = CLBLM_R_X63Y102_SLICE_X94Y102_DO6;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_DMUX = CLBLM_R_X63Y102_SLICE_X94Y102_DO5;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_A = CLBLM_R_X63Y102_SLICE_X95Y102_AO6;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_B = CLBLM_R_X63Y102_SLICE_X95Y102_BO6;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_C = CLBLM_R_X63Y102_SLICE_X95Y102_CO6;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_D = CLBLM_R_X63Y102_SLICE_X95Y102_DO6;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_AMUX = CLBLM_R_X63Y102_SLICE_X95Y102_AO5;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_A = CLBLM_R_X63Y103_SLICE_X94Y103_AO6;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_B = CLBLM_R_X63Y103_SLICE_X94Y103_BO6;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_C = CLBLM_R_X63Y103_SLICE_X94Y103_CO6;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_D = CLBLM_R_X63Y103_SLICE_X94Y103_DO6;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_AMUX = CLBLM_R_X63Y103_SLICE_X94Y103_AO5;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_A = CLBLM_R_X63Y103_SLICE_X95Y103_AO6;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_B = CLBLM_R_X63Y103_SLICE_X95Y103_BO6;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_C = CLBLM_R_X63Y103_SLICE_X95Y103_CO6;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_D = CLBLM_R_X63Y103_SLICE_X95Y103_DO6;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_BMUX = CLBLM_R_X63Y103_SLICE_X95Y103_BO5;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_A = CLBLM_R_X63Y105_SLICE_X94Y105_AO6;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_B = CLBLM_R_X63Y105_SLICE_X94Y105_BO6;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_C = CLBLM_R_X63Y105_SLICE_X94Y105_CO6;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_D = CLBLM_R_X63Y105_SLICE_X94Y105_DO6;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_CMUX = CLBLM_R_X63Y105_SLICE_X94Y105_C5Q;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_A = CLBLM_R_X63Y105_SLICE_X95Y105_AO6;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_B = CLBLM_R_X63Y105_SLICE_X95Y105_BO6;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_C = CLBLM_R_X63Y105_SLICE_X95Y105_CO6;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_D = CLBLM_R_X63Y105_SLICE_X95Y105_DO6;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_AMUX = CLBLM_R_X63Y105_SLICE_X95Y105_A5Q;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_CMUX = CLBLM_R_X63Y105_SLICE_X95Y105_C5Q;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_A = CLBLM_R_X63Y106_SLICE_X94Y106_AO6;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_B = CLBLM_R_X63Y106_SLICE_X94Y106_BO6;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_C = CLBLM_R_X63Y106_SLICE_X94Y106_CO6;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_D = CLBLM_R_X63Y106_SLICE_X94Y106_DO6;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_AMUX = CLBLM_R_X63Y106_SLICE_X94Y106_AO5;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_A = CLBLM_R_X63Y106_SLICE_X95Y106_AO6;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_B = CLBLM_R_X63Y106_SLICE_X95Y106_BO6;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_C = CLBLM_R_X63Y106_SLICE_X95Y106_CO6;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_D = CLBLM_R_X63Y106_SLICE_X95Y106_DO6;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_DMUX = CLBLM_R_X63Y106_SLICE_X95Y106_DO6;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_A = CLBLM_R_X63Y107_SLICE_X94Y107_AO6;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_B = CLBLM_R_X63Y107_SLICE_X94Y107_BO6;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_C = CLBLM_R_X63Y107_SLICE_X94Y107_CO6;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_D = CLBLM_R_X63Y107_SLICE_X94Y107_DO6;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_CMUX = CLBLM_R_X63Y107_SLICE_X94Y107_CO6;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_A = CLBLM_R_X63Y107_SLICE_X95Y107_AO6;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_B = CLBLM_R_X63Y107_SLICE_X95Y107_BO6;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_C = CLBLM_R_X63Y107_SLICE_X95Y107_CO6;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_D = CLBLM_R_X63Y107_SLICE_X95Y107_DO6;
  assign CLBLM_R_X63Y122_SLICE_X94Y122_A = CLBLM_R_X63Y122_SLICE_X94Y122_AO6;
  assign CLBLM_R_X63Y122_SLICE_X94Y122_B = CLBLM_R_X63Y122_SLICE_X94Y122_BO6;
  assign CLBLM_R_X63Y122_SLICE_X94Y122_C = CLBLM_R_X63Y122_SLICE_X94Y122_CO6;
  assign CLBLM_R_X63Y122_SLICE_X94Y122_D = CLBLM_R_X63Y122_SLICE_X94Y122_DO6;
  assign CLBLM_R_X63Y122_SLICE_X95Y122_A = CLBLM_R_X63Y122_SLICE_X95Y122_AO6;
  assign CLBLM_R_X63Y122_SLICE_X95Y122_B = CLBLM_R_X63Y122_SLICE_X95Y122_BO6;
  assign CLBLM_R_X63Y122_SLICE_X95Y122_C = CLBLM_R_X63Y122_SLICE_X95Y122_CO6;
  assign CLBLM_R_X63Y122_SLICE_X95Y122_D = CLBLM_R_X63Y122_SLICE_X95Y122_DO6;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_A = CLBLM_R_X65Y99_SLICE_X98Y99_AO6;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_B = CLBLM_R_X65Y99_SLICE_X98Y99_BO6;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_C = CLBLM_R_X65Y99_SLICE_X98Y99_CO6;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_D = CLBLM_R_X65Y99_SLICE_X98Y99_DO6;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_A = CLBLM_R_X65Y99_SLICE_X99Y99_AO6;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_B = CLBLM_R_X65Y99_SLICE_X99Y99_BO6;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_C = CLBLM_R_X65Y99_SLICE_X99Y99_CO6;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_D = CLBLM_R_X65Y99_SLICE_X99Y99_DO6;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_CMUX = CLBLM_R_X65Y99_SLICE_X99Y99_C5Q;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_A = CLBLM_R_X65Y100_SLICE_X98Y100_AO6;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_B = CLBLM_R_X65Y100_SLICE_X98Y100_BO6;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_C = CLBLM_R_X65Y100_SLICE_X98Y100_CO6;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_D = CLBLM_R_X65Y100_SLICE_X98Y100_DO6;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_A = CLBLM_R_X65Y100_SLICE_X99Y100_AO6;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_B = CLBLM_R_X65Y100_SLICE_X99Y100_BO6;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_C = CLBLM_R_X65Y100_SLICE_X99Y100_CO6;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_D = CLBLM_R_X65Y100_SLICE_X99Y100_DO6;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_AMUX = CLBLM_R_X65Y100_SLICE_X99Y100_A5Q;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_A = CLBLM_R_X65Y101_SLICE_X98Y101_AO6;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_B = CLBLM_R_X65Y101_SLICE_X98Y101_BO6;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_C = CLBLM_R_X65Y101_SLICE_X98Y101_CO6;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_D = CLBLM_R_X65Y101_SLICE_X98Y101_DO6;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_A = CLBLM_R_X65Y101_SLICE_X99Y101_AO6;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_B = CLBLM_R_X65Y101_SLICE_X99Y101_BO6;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_C = CLBLM_R_X65Y101_SLICE_X99Y101_CO6;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_D = CLBLM_R_X65Y101_SLICE_X99Y101_DO6;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_A = CLBLM_R_X65Y102_SLICE_X98Y102_AO6;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_B = CLBLM_R_X65Y102_SLICE_X98Y102_BO6;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_C = CLBLM_R_X65Y102_SLICE_X98Y102_CO6;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_D = CLBLM_R_X65Y102_SLICE_X98Y102_DO6;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_A = CLBLM_R_X65Y102_SLICE_X99Y102_AO6;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_B = CLBLM_R_X65Y102_SLICE_X99Y102_BO6;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_C = CLBLM_R_X65Y102_SLICE_X99Y102_CO6;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_D = CLBLM_R_X65Y102_SLICE_X99Y102_DO6;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_A = CLBLM_R_X65Y103_SLICE_X98Y103_AO6;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_B = CLBLM_R_X65Y103_SLICE_X98Y103_BO6;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_C = CLBLM_R_X65Y103_SLICE_X98Y103_CO6;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_D = CLBLM_R_X65Y103_SLICE_X98Y103_DO6;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_AMUX = CLBLM_R_X65Y103_SLICE_X98Y103_A5Q;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_A = CLBLM_R_X65Y103_SLICE_X99Y103_AO6;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_B = CLBLM_R_X65Y103_SLICE_X99Y103_BO6;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_C = CLBLM_R_X65Y103_SLICE_X99Y103_CO6;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_D = CLBLM_R_X65Y103_SLICE_X99Y103_DO6;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_DMUX = CLBLM_R_X65Y103_SLICE_X99Y103_DO6;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_A = CLBLM_R_X65Y104_SLICE_X98Y104_AO6;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_B = CLBLM_R_X65Y104_SLICE_X98Y104_BO6;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_C = CLBLM_R_X65Y104_SLICE_X98Y104_CO6;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_D = CLBLM_R_X65Y104_SLICE_X98Y104_DO6;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_AMUX = CLBLM_R_X65Y104_SLICE_X98Y104_AO5;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_BMUX = CLBLM_R_X65Y104_SLICE_X98Y104_B5Q;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_CMUX = CLBLM_R_X65Y104_SLICE_X98Y104_C5Q;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_A = CLBLM_R_X65Y104_SLICE_X99Y104_AO6;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_B = CLBLM_R_X65Y104_SLICE_X99Y104_BO6;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_C = CLBLM_R_X65Y104_SLICE_X99Y104_CO6;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_D = CLBLM_R_X65Y104_SLICE_X99Y104_DO6;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_AMUX = CLBLM_R_X65Y104_SLICE_X99Y104_A5Q;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_BMUX = CLBLM_R_X65Y104_SLICE_X99Y104_B5Q;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_A = CLBLM_R_X65Y105_SLICE_X98Y105_AO6;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_B = CLBLM_R_X65Y105_SLICE_X98Y105_BO6;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_C = CLBLM_R_X65Y105_SLICE_X98Y105_CO6;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_D = CLBLM_R_X65Y105_SLICE_X98Y105_DO6;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_BMUX = CLBLM_R_X65Y105_SLICE_X98Y105_B5Q;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_A = CLBLM_R_X65Y105_SLICE_X99Y105_AO6;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_B = CLBLM_R_X65Y105_SLICE_X99Y105_BO6;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_C = CLBLM_R_X65Y105_SLICE_X99Y105_CO6;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_D = CLBLM_R_X65Y105_SLICE_X99Y105_DO6;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_BMUX = CLBLM_R_X65Y105_SLICE_X99Y105_BO5;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_CMUX = CLBLM_R_X65Y105_SLICE_X99Y105_C5Q;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_DMUX = CLBLM_R_X65Y105_SLICE_X99Y105_D5Q;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_A = CLBLM_R_X65Y106_SLICE_X98Y106_AO6;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_B = CLBLM_R_X65Y106_SLICE_X98Y106_BO6;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_C = CLBLM_R_X65Y106_SLICE_X98Y106_CO6;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_D = CLBLM_R_X65Y106_SLICE_X98Y106_DO6;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_A = CLBLM_R_X65Y106_SLICE_X99Y106_AO6;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_B = CLBLM_R_X65Y106_SLICE_X99Y106_BO6;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_C = CLBLM_R_X65Y106_SLICE_X99Y106_CO6;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_D = CLBLM_R_X65Y106_SLICE_X99Y106_DO6;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_CMUX = CLBLM_R_X65Y106_SLICE_X99Y106_C5Q;
  assign CLBLM_R_X65Y108_SLICE_X98Y108_A = CLBLM_R_X65Y108_SLICE_X98Y108_AO6;
  assign CLBLM_R_X65Y108_SLICE_X98Y108_B = CLBLM_R_X65Y108_SLICE_X98Y108_BO6;
  assign CLBLM_R_X65Y108_SLICE_X98Y108_C = CLBLM_R_X65Y108_SLICE_X98Y108_CO6;
  assign CLBLM_R_X65Y108_SLICE_X98Y108_D = CLBLM_R_X65Y108_SLICE_X98Y108_DO6;
  assign CLBLM_R_X65Y108_SLICE_X99Y108_A = CLBLM_R_X65Y108_SLICE_X99Y108_AO6;
  assign CLBLM_R_X65Y108_SLICE_X99Y108_B = CLBLM_R_X65Y108_SLICE_X99Y108_BO6;
  assign CLBLM_R_X65Y108_SLICE_X99Y108_C = CLBLM_R_X65Y108_SLICE_X99Y108_CO6;
  assign CLBLM_R_X65Y108_SLICE_X99Y108_D = CLBLM_R_X65Y108_SLICE_X99Y108_DO6;
  assign CLBLM_R_X65Y108_SLICE_X99Y108_CMUX = CLBLM_R_X65Y108_SLICE_X99Y108_CO6;
  assign CLBLM_R_X65Y109_SLICE_X98Y109_A = CLBLM_R_X65Y109_SLICE_X98Y109_AO6;
  assign CLBLM_R_X65Y109_SLICE_X98Y109_B = CLBLM_R_X65Y109_SLICE_X98Y109_BO6;
  assign CLBLM_R_X65Y109_SLICE_X98Y109_C = CLBLM_R_X65Y109_SLICE_X98Y109_CO6;
  assign CLBLM_R_X65Y109_SLICE_X98Y109_D = CLBLM_R_X65Y109_SLICE_X98Y109_DO6;
  assign CLBLM_R_X65Y109_SLICE_X98Y109_AMUX = CLBLM_R_X65Y109_SLICE_X98Y109_A5Q;
  assign CLBLM_R_X65Y109_SLICE_X99Y109_A = CLBLM_R_X65Y109_SLICE_X99Y109_AO6;
  assign CLBLM_R_X65Y109_SLICE_X99Y109_B = CLBLM_R_X65Y109_SLICE_X99Y109_BO6;
  assign CLBLM_R_X65Y109_SLICE_X99Y109_C = CLBLM_R_X65Y109_SLICE_X99Y109_CO6;
  assign CLBLM_R_X65Y109_SLICE_X99Y109_D = CLBLM_R_X65Y109_SLICE_X99Y109_DO6;
  assign CLBLM_R_X65Y109_SLICE_X99Y109_AMUX = CLBLM_R_X65Y109_SLICE_X99Y109_A5Q;
  assign CLBLM_R_X65Y109_SLICE_X99Y109_DMUX = CLBLM_R_X65Y109_SLICE_X99Y109_DO5;
  assign CLBLM_R_X65Y110_SLICE_X98Y110_A = CLBLM_R_X65Y110_SLICE_X98Y110_AO6;
  assign CLBLM_R_X65Y110_SLICE_X98Y110_B = CLBLM_R_X65Y110_SLICE_X98Y110_BO6;
  assign CLBLM_R_X65Y110_SLICE_X98Y110_C = CLBLM_R_X65Y110_SLICE_X98Y110_CO6;
  assign CLBLM_R_X65Y110_SLICE_X98Y110_D = CLBLM_R_X65Y110_SLICE_X98Y110_DO6;
  assign CLBLM_R_X65Y110_SLICE_X98Y110_AMUX = CLBLM_R_X65Y110_SLICE_X98Y110_A5Q;
  assign CLBLM_R_X65Y110_SLICE_X99Y110_A = CLBLM_R_X65Y110_SLICE_X99Y110_AO6;
  assign CLBLM_R_X65Y110_SLICE_X99Y110_B = CLBLM_R_X65Y110_SLICE_X99Y110_BO6;
  assign CLBLM_R_X65Y110_SLICE_X99Y110_C = CLBLM_R_X65Y110_SLICE_X99Y110_CO6;
  assign CLBLM_R_X65Y110_SLICE_X99Y110_D = CLBLM_R_X65Y110_SLICE_X99Y110_DO6;
  assign CLBLM_R_X65Y110_SLICE_X99Y110_AMUX = CLBLM_R_X65Y110_SLICE_X99Y110_AO5;
  assign CLBLM_R_X65Y110_SLICE_X99Y110_BMUX = CLBLM_R_X65Y110_SLICE_X99Y110_B5Q;
  assign CLBLM_R_X65Y111_SLICE_X98Y111_A = CLBLM_R_X65Y111_SLICE_X98Y111_AO6;
  assign CLBLM_R_X65Y111_SLICE_X98Y111_B = CLBLM_R_X65Y111_SLICE_X98Y111_BO6;
  assign CLBLM_R_X65Y111_SLICE_X98Y111_C = CLBLM_R_X65Y111_SLICE_X98Y111_CO6;
  assign CLBLM_R_X65Y111_SLICE_X98Y111_D = CLBLM_R_X65Y111_SLICE_X98Y111_DO6;
  assign CLBLM_R_X65Y111_SLICE_X99Y111_A = CLBLM_R_X65Y111_SLICE_X99Y111_AO6;
  assign CLBLM_R_X65Y111_SLICE_X99Y111_B = CLBLM_R_X65Y111_SLICE_X99Y111_BO6;
  assign CLBLM_R_X65Y111_SLICE_X99Y111_C = CLBLM_R_X65Y111_SLICE_X99Y111_CO6;
  assign CLBLM_R_X65Y111_SLICE_X99Y111_D = CLBLM_R_X65Y111_SLICE_X99Y111_DO6;
  assign CLBLM_R_X65Y111_SLICE_X99Y111_AMUX = CLBLM_R_X65Y111_SLICE_X99Y111_AO5;
  assign CLBLM_R_X67Y96_SLICE_X100Y96_A = CLBLM_R_X67Y96_SLICE_X100Y96_AO6;
  assign CLBLM_R_X67Y96_SLICE_X100Y96_B = CLBLM_R_X67Y96_SLICE_X100Y96_BO6;
  assign CLBLM_R_X67Y96_SLICE_X100Y96_C = CLBLM_R_X67Y96_SLICE_X100Y96_CO6;
  assign CLBLM_R_X67Y96_SLICE_X100Y96_D = CLBLM_R_X67Y96_SLICE_X100Y96_DO6;
  assign CLBLM_R_X67Y96_SLICE_X101Y96_A = CLBLM_R_X67Y96_SLICE_X101Y96_AO6;
  assign CLBLM_R_X67Y96_SLICE_X101Y96_B = CLBLM_R_X67Y96_SLICE_X101Y96_BO6;
  assign CLBLM_R_X67Y96_SLICE_X101Y96_C = CLBLM_R_X67Y96_SLICE_X101Y96_CO6;
  assign CLBLM_R_X67Y96_SLICE_X101Y96_D = CLBLM_R_X67Y96_SLICE_X101Y96_DO6;
  assign CLBLM_R_X67Y97_SLICE_X100Y97_A = CLBLM_R_X67Y97_SLICE_X100Y97_AO6;
  assign CLBLM_R_X67Y97_SLICE_X100Y97_B = CLBLM_R_X67Y97_SLICE_X100Y97_BO6;
  assign CLBLM_R_X67Y97_SLICE_X100Y97_C = CLBLM_R_X67Y97_SLICE_X100Y97_CO6;
  assign CLBLM_R_X67Y97_SLICE_X100Y97_D = CLBLM_R_X67Y97_SLICE_X100Y97_DO6;
  assign CLBLM_R_X67Y97_SLICE_X101Y97_A = CLBLM_R_X67Y97_SLICE_X101Y97_AO6;
  assign CLBLM_R_X67Y97_SLICE_X101Y97_B = CLBLM_R_X67Y97_SLICE_X101Y97_BO6;
  assign CLBLM_R_X67Y97_SLICE_X101Y97_C = CLBLM_R_X67Y97_SLICE_X101Y97_CO6;
  assign CLBLM_R_X67Y97_SLICE_X101Y97_D = CLBLM_R_X67Y97_SLICE_X101Y97_DO6;
  assign CLBLM_R_X67Y98_SLICE_X100Y98_A = CLBLM_R_X67Y98_SLICE_X100Y98_AO6;
  assign CLBLM_R_X67Y98_SLICE_X100Y98_B = CLBLM_R_X67Y98_SLICE_X100Y98_BO6;
  assign CLBLM_R_X67Y98_SLICE_X100Y98_C = CLBLM_R_X67Y98_SLICE_X100Y98_CO6;
  assign CLBLM_R_X67Y98_SLICE_X100Y98_D = CLBLM_R_X67Y98_SLICE_X100Y98_DO6;
  assign CLBLM_R_X67Y98_SLICE_X100Y98_AMUX = CLBLM_R_X67Y98_SLICE_X100Y98_A5Q;
  assign CLBLM_R_X67Y98_SLICE_X100Y98_BMUX = CLBLM_R_X67Y98_SLICE_X100Y98_B5Q;
  assign CLBLM_R_X67Y98_SLICE_X100Y98_CMUX = CLBLM_R_X67Y98_SLICE_X100Y98_CO5;
  assign CLBLM_R_X67Y98_SLICE_X101Y98_A = CLBLM_R_X67Y98_SLICE_X101Y98_AO6;
  assign CLBLM_R_X67Y98_SLICE_X101Y98_B = CLBLM_R_X67Y98_SLICE_X101Y98_BO6;
  assign CLBLM_R_X67Y98_SLICE_X101Y98_C = CLBLM_R_X67Y98_SLICE_X101Y98_CO6;
  assign CLBLM_R_X67Y98_SLICE_X101Y98_D = CLBLM_R_X67Y98_SLICE_X101Y98_DO6;
  assign CLBLM_R_X67Y98_SLICE_X101Y98_AMUX = CLBLM_R_X67Y98_SLICE_X101Y98_AO5;
  assign CLBLM_R_X67Y98_SLICE_X101Y98_BMUX = CLBLM_R_X67Y98_SLICE_X101Y98_BO5;
  assign CLBLM_R_X67Y98_SLICE_X101Y98_CMUX = CLBLM_R_X67Y98_SLICE_X101Y98_CO5;
  assign CLBLM_R_X67Y99_SLICE_X100Y99_A = CLBLM_R_X67Y99_SLICE_X100Y99_AO6;
  assign CLBLM_R_X67Y99_SLICE_X100Y99_B = CLBLM_R_X67Y99_SLICE_X100Y99_BO6;
  assign CLBLM_R_X67Y99_SLICE_X100Y99_C = CLBLM_R_X67Y99_SLICE_X100Y99_CO6;
  assign CLBLM_R_X67Y99_SLICE_X100Y99_D = CLBLM_R_X67Y99_SLICE_X100Y99_DO6;
  assign CLBLM_R_X67Y99_SLICE_X101Y99_A = CLBLM_R_X67Y99_SLICE_X101Y99_AO6;
  assign CLBLM_R_X67Y99_SLICE_X101Y99_B = CLBLM_R_X67Y99_SLICE_X101Y99_BO6;
  assign CLBLM_R_X67Y99_SLICE_X101Y99_C = CLBLM_R_X67Y99_SLICE_X101Y99_CO6;
  assign CLBLM_R_X67Y99_SLICE_X101Y99_D = CLBLM_R_X67Y99_SLICE_X101Y99_DO6;
  assign CLBLM_R_X67Y100_SLICE_X100Y100_A = CLBLM_R_X67Y100_SLICE_X100Y100_AO6;
  assign CLBLM_R_X67Y100_SLICE_X100Y100_B = CLBLM_R_X67Y100_SLICE_X100Y100_BO6;
  assign CLBLM_R_X67Y100_SLICE_X100Y100_C = CLBLM_R_X67Y100_SLICE_X100Y100_CO6;
  assign CLBLM_R_X67Y100_SLICE_X100Y100_D = CLBLM_R_X67Y100_SLICE_X100Y100_DO6;
  assign CLBLM_R_X67Y100_SLICE_X100Y100_AMUX = CLBLM_R_X67Y100_SLICE_X100Y100_A5Q;
  assign CLBLM_R_X67Y100_SLICE_X101Y100_A = CLBLM_R_X67Y100_SLICE_X101Y100_AO6;
  assign CLBLM_R_X67Y100_SLICE_X101Y100_B = CLBLM_R_X67Y100_SLICE_X101Y100_BO6;
  assign CLBLM_R_X67Y100_SLICE_X101Y100_C = CLBLM_R_X67Y100_SLICE_X101Y100_CO6;
  assign CLBLM_R_X67Y100_SLICE_X101Y100_D = CLBLM_R_X67Y100_SLICE_X101Y100_DO6;
  assign CLBLM_R_X67Y101_SLICE_X100Y101_A = CLBLM_R_X67Y101_SLICE_X100Y101_AO6;
  assign CLBLM_R_X67Y101_SLICE_X100Y101_B = CLBLM_R_X67Y101_SLICE_X100Y101_BO6;
  assign CLBLM_R_X67Y101_SLICE_X100Y101_C = CLBLM_R_X67Y101_SLICE_X100Y101_CO6;
  assign CLBLM_R_X67Y101_SLICE_X100Y101_D = CLBLM_R_X67Y101_SLICE_X100Y101_DO6;
  assign CLBLM_R_X67Y101_SLICE_X100Y101_BMUX = CLBLM_R_X67Y101_SLICE_X100Y101_BO5;
  assign CLBLM_R_X67Y101_SLICE_X101Y101_A = CLBLM_R_X67Y101_SLICE_X101Y101_AO6;
  assign CLBLM_R_X67Y101_SLICE_X101Y101_B = CLBLM_R_X67Y101_SLICE_X101Y101_BO6;
  assign CLBLM_R_X67Y101_SLICE_X101Y101_C = CLBLM_R_X67Y101_SLICE_X101Y101_CO6;
  assign CLBLM_R_X67Y101_SLICE_X101Y101_D = CLBLM_R_X67Y101_SLICE_X101Y101_DO6;
  assign CLBLM_R_X67Y101_SLICE_X101Y101_CMUX = CLBLM_R_X67Y101_SLICE_X101Y101_CO6;
  assign CLBLM_R_X67Y103_SLICE_X100Y103_A = CLBLM_R_X67Y103_SLICE_X100Y103_AO6;
  assign CLBLM_R_X67Y103_SLICE_X100Y103_B = CLBLM_R_X67Y103_SLICE_X100Y103_BO6;
  assign CLBLM_R_X67Y103_SLICE_X100Y103_C = CLBLM_R_X67Y103_SLICE_X100Y103_CO6;
  assign CLBLM_R_X67Y103_SLICE_X100Y103_D = CLBLM_R_X67Y103_SLICE_X100Y103_DO6;
  assign CLBLM_R_X67Y103_SLICE_X100Y103_AMUX = CLBLM_R_X67Y103_SLICE_X100Y103_AO5;
  assign CLBLM_R_X67Y103_SLICE_X100Y103_BMUX = CLBLM_R_X67Y103_SLICE_X100Y103_B5Q;
  assign CLBLM_R_X67Y103_SLICE_X101Y103_A = CLBLM_R_X67Y103_SLICE_X101Y103_AO6;
  assign CLBLM_R_X67Y103_SLICE_X101Y103_B = CLBLM_R_X67Y103_SLICE_X101Y103_BO6;
  assign CLBLM_R_X67Y103_SLICE_X101Y103_C = CLBLM_R_X67Y103_SLICE_X101Y103_CO6;
  assign CLBLM_R_X67Y103_SLICE_X101Y103_D = CLBLM_R_X67Y103_SLICE_X101Y103_DO6;
  assign CLBLM_R_X67Y105_SLICE_X100Y105_A = CLBLM_R_X67Y105_SLICE_X100Y105_AO6;
  assign CLBLM_R_X67Y105_SLICE_X100Y105_B = CLBLM_R_X67Y105_SLICE_X100Y105_BO6;
  assign CLBLM_R_X67Y105_SLICE_X100Y105_C = CLBLM_R_X67Y105_SLICE_X100Y105_CO6;
  assign CLBLM_R_X67Y105_SLICE_X100Y105_D = CLBLM_R_X67Y105_SLICE_X100Y105_DO6;
  assign CLBLM_R_X67Y105_SLICE_X100Y105_AMUX = CLBLM_R_X67Y105_SLICE_X100Y105_AO6;
  assign CLBLM_R_X67Y105_SLICE_X100Y105_CMUX = CLBLM_R_X67Y105_SLICE_X100Y105_CO5;
  assign CLBLM_R_X67Y105_SLICE_X100Y105_DMUX = CLBLM_R_X67Y105_SLICE_X100Y105_DO5;
  assign CLBLM_R_X67Y105_SLICE_X101Y105_A = CLBLM_R_X67Y105_SLICE_X101Y105_AO6;
  assign CLBLM_R_X67Y105_SLICE_X101Y105_B = CLBLM_R_X67Y105_SLICE_X101Y105_BO6;
  assign CLBLM_R_X67Y105_SLICE_X101Y105_C = CLBLM_R_X67Y105_SLICE_X101Y105_CO6;
  assign CLBLM_R_X67Y105_SLICE_X101Y105_D = CLBLM_R_X67Y105_SLICE_X101Y105_DO6;
  assign CLBLM_R_X67Y105_SLICE_X101Y105_DMUX = CLBLM_R_X67Y105_SLICE_X101Y105_DO6;
  assign CLBLM_R_X67Y108_SLICE_X100Y108_A = CLBLM_R_X67Y108_SLICE_X100Y108_AO6;
  assign CLBLM_R_X67Y108_SLICE_X100Y108_B = CLBLM_R_X67Y108_SLICE_X100Y108_BO6;
  assign CLBLM_R_X67Y108_SLICE_X100Y108_C = CLBLM_R_X67Y108_SLICE_X100Y108_CO6;
  assign CLBLM_R_X67Y108_SLICE_X100Y108_D = CLBLM_R_X67Y108_SLICE_X100Y108_DO6;
  assign CLBLM_R_X67Y108_SLICE_X100Y108_BMUX = CLBLM_R_X67Y108_SLICE_X100Y108_BO5;
  assign CLBLM_R_X67Y108_SLICE_X100Y108_CMUX = CLBLM_R_X67Y108_SLICE_X100Y108_C5Q;
  assign CLBLM_R_X67Y108_SLICE_X101Y108_A = CLBLM_R_X67Y108_SLICE_X101Y108_AO6;
  assign CLBLM_R_X67Y108_SLICE_X101Y108_B = CLBLM_R_X67Y108_SLICE_X101Y108_BO6;
  assign CLBLM_R_X67Y108_SLICE_X101Y108_C = CLBLM_R_X67Y108_SLICE_X101Y108_CO6;
  assign CLBLM_R_X67Y108_SLICE_X101Y108_D = CLBLM_R_X67Y108_SLICE_X101Y108_DO6;
  assign CLBLM_R_X67Y108_SLICE_X101Y108_AMUX = CLBLM_R_X67Y108_SLICE_X101Y108_AO5;
  assign CLBLM_R_X67Y109_SLICE_X100Y109_A = CLBLM_R_X67Y109_SLICE_X100Y109_AO6;
  assign CLBLM_R_X67Y109_SLICE_X100Y109_B = CLBLM_R_X67Y109_SLICE_X100Y109_BO6;
  assign CLBLM_R_X67Y109_SLICE_X100Y109_C = CLBLM_R_X67Y109_SLICE_X100Y109_CO6;
  assign CLBLM_R_X67Y109_SLICE_X100Y109_D = CLBLM_R_X67Y109_SLICE_X100Y109_DO6;
  assign CLBLM_R_X67Y109_SLICE_X100Y109_DMUX = CLBLM_R_X67Y109_SLICE_X100Y109_DO5;
  assign CLBLM_R_X67Y109_SLICE_X101Y109_A = CLBLM_R_X67Y109_SLICE_X101Y109_AO6;
  assign CLBLM_R_X67Y109_SLICE_X101Y109_B = CLBLM_R_X67Y109_SLICE_X101Y109_BO6;
  assign CLBLM_R_X67Y109_SLICE_X101Y109_C = CLBLM_R_X67Y109_SLICE_X101Y109_CO6;
  assign CLBLM_R_X67Y109_SLICE_X101Y109_D = CLBLM_R_X67Y109_SLICE_X101Y109_DO6;
  assign CLBLM_R_X67Y110_SLICE_X100Y110_A = CLBLM_R_X67Y110_SLICE_X100Y110_AO6;
  assign CLBLM_R_X67Y110_SLICE_X100Y110_B = CLBLM_R_X67Y110_SLICE_X100Y110_BO6;
  assign CLBLM_R_X67Y110_SLICE_X100Y110_C = CLBLM_R_X67Y110_SLICE_X100Y110_CO6;
  assign CLBLM_R_X67Y110_SLICE_X100Y110_D = CLBLM_R_X67Y110_SLICE_X100Y110_DO6;
  assign CLBLM_R_X67Y110_SLICE_X101Y110_A = CLBLM_R_X67Y110_SLICE_X101Y110_AO6;
  assign CLBLM_R_X67Y110_SLICE_X101Y110_B = CLBLM_R_X67Y110_SLICE_X101Y110_BO6;
  assign CLBLM_R_X67Y110_SLICE_X101Y110_C = CLBLM_R_X67Y110_SLICE_X101Y110_CO6;
  assign CLBLM_R_X67Y110_SLICE_X101Y110_D = CLBLM_R_X67Y110_SLICE_X101Y110_DO6;
  assign CLBLM_R_X67Y111_SLICE_X100Y111_A = CLBLM_R_X67Y111_SLICE_X100Y111_AO6;
  assign CLBLM_R_X67Y111_SLICE_X100Y111_B = CLBLM_R_X67Y111_SLICE_X100Y111_BO6;
  assign CLBLM_R_X67Y111_SLICE_X100Y111_C = CLBLM_R_X67Y111_SLICE_X100Y111_CO6;
  assign CLBLM_R_X67Y111_SLICE_X100Y111_D = CLBLM_R_X67Y111_SLICE_X100Y111_DO6;
  assign CLBLM_R_X67Y111_SLICE_X100Y111_AMUX = CLBLM_R_X67Y111_SLICE_X100Y111_A5Q;
  assign CLBLM_R_X67Y111_SLICE_X100Y111_CMUX = CLBLM_R_X67Y111_SLICE_X100Y111_CO5;
  assign CLBLM_R_X67Y111_SLICE_X101Y111_A = CLBLM_R_X67Y111_SLICE_X101Y111_AO6;
  assign CLBLM_R_X67Y111_SLICE_X101Y111_B = CLBLM_R_X67Y111_SLICE_X101Y111_BO6;
  assign CLBLM_R_X67Y111_SLICE_X101Y111_C = CLBLM_R_X67Y111_SLICE_X101Y111_CO6;
  assign CLBLM_R_X67Y111_SLICE_X101Y111_D = CLBLM_R_X67Y111_SLICE_X101Y111_DO6;
  assign CLBLM_R_X67Y111_SLICE_X101Y111_AMUX = CLBLM_R_X67Y111_SLICE_X101Y111_A5Q;
  assign CLBLM_R_X67Y111_SLICE_X101Y111_BMUX = CLBLM_R_X67Y111_SLICE_X101Y111_B5Q;
  assign CLBLM_R_X67Y111_SLICE_X101Y111_CMUX = CLBLM_R_X67Y111_SLICE_X101Y111_CO5;
  assign CLBLM_R_X67Y111_SLICE_X101Y111_DMUX = CLBLM_R_X67Y111_SLICE_X101Y111_DO5;
  assign CLBLM_R_X67Y115_SLICE_X100Y115_A = CLBLM_R_X67Y115_SLICE_X100Y115_AO6;
  assign CLBLM_R_X67Y115_SLICE_X100Y115_B = CLBLM_R_X67Y115_SLICE_X100Y115_BO6;
  assign CLBLM_R_X67Y115_SLICE_X100Y115_C = CLBLM_R_X67Y115_SLICE_X100Y115_CO6;
  assign CLBLM_R_X67Y115_SLICE_X100Y115_D = CLBLM_R_X67Y115_SLICE_X100Y115_DO6;
  assign CLBLM_R_X67Y115_SLICE_X100Y115_AMUX = CLBLM_R_X67Y115_SLICE_X100Y115_A5Q;
  assign CLBLM_R_X67Y115_SLICE_X101Y115_A = CLBLM_R_X67Y115_SLICE_X101Y115_AO6;
  assign CLBLM_R_X67Y115_SLICE_X101Y115_B = CLBLM_R_X67Y115_SLICE_X101Y115_BO6;
  assign CLBLM_R_X67Y115_SLICE_X101Y115_C = CLBLM_R_X67Y115_SLICE_X101Y115_CO6;
  assign CLBLM_R_X67Y115_SLICE_X101Y115_D = CLBLM_R_X67Y115_SLICE_X101Y115_DO6;
  assign CLBLM_R_X67Y116_SLICE_X100Y116_A = CLBLM_R_X67Y116_SLICE_X100Y116_AO6;
  assign CLBLM_R_X67Y116_SLICE_X100Y116_B = CLBLM_R_X67Y116_SLICE_X100Y116_BO6;
  assign CLBLM_R_X67Y116_SLICE_X100Y116_C = CLBLM_R_X67Y116_SLICE_X100Y116_CO6;
  assign CLBLM_R_X67Y116_SLICE_X100Y116_D = CLBLM_R_X67Y116_SLICE_X100Y116_DO6;
  assign CLBLM_R_X67Y116_SLICE_X100Y116_BMUX = CLBLM_R_X67Y116_SLICE_X100Y116_B5Q;
  assign CLBLM_R_X67Y116_SLICE_X100Y116_CMUX = CLBLM_R_X67Y116_SLICE_X100Y116_C5Q;
  assign CLBLM_R_X67Y116_SLICE_X101Y116_A = CLBLM_R_X67Y116_SLICE_X101Y116_AO6;
  assign CLBLM_R_X67Y116_SLICE_X101Y116_B = CLBLM_R_X67Y116_SLICE_X101Y116_BO6;
  assign CLBLM_R_X67Y116_SLICE_X101Y116_C = CLBLM_R_X67Y116_SLICE_X101Y116_CO6;
  assign CLBLM_R_X67Y116_SLICE_X101Y116_D = CLBLM_R_X67Y116_SLICE_X101Y116_DO6;
  assign CLBLM_R_X67Y116_SLICE_X101Y116_AMUX = CLBLM_R_X67Y116_SLICE_X101Y116_A5Q;
  assign CLBLM_R_X67Y118_SLICE_X100Y118_A = CLBLM_R_X67Y118_SLICE_X100Y118_AO6;
  assign CLBLM_R_X67Y118_SLICE_X100Y118_B = CLBLM_R_X67Y118_SLICE_X100Y118_BO6;
  assign CLBLM_R_X67Y118_SLICE_X100Y118_C = CLBLM_R_X67Y118_SLICE_X100Y118_CO6;
  assign CLBLM_R_X67Y118_SLICE_X100Y118_D = CLBLM_R_X67Y118_SLICE_X100Y118_DO6;
  assign CLBLM_R_X67Y118_SLICE_X100Y118_AMUX = CLBLM_R_X67Y118_SLICE_X100Y118_A5Q;
  assign CLBLM_R_X67Y118_SLICE_X101Y118_A = CLBLM_R_X67Y118_SLICE_X101Y118_AO6;
  assign CLBLM_R_X67Y118_SLICE_X101Y118_B = CLBLM_R_X67Y118_SLICE_X101Y118_BO6;
  assign CLBLM_R_X67Y118_SLICE_X101Y118_C = CLBLM_R_X67Y118_SLICE_X101Y118_CO6;
  assign CLBLM_R_X67Y118_SLICE_X101Y118_D = CLBLM_R_X67Y118_SLICE_X101Y118_DO6;
  assign CLBLM_R_X67Y118_SLICE_X101Y118_AMUX = CLBLM_R_X67Y118_SLICE_X101Y118_A5Q;
  assign CLBLM_R_X103Y67_SLICE_X162Y67_A = CLBLM_R_X103Y67_SLICE_X162Y67_AO6;
  assign CLBLM_R_X103Y67_SLICE_X162Y67_B = CLBLM_R_X103Y67_SLICE_X162Y67_BO6;
  assign CLBLM_R_X103Y67_SLICE_X162Y67_C = CLBLM_R_X103Y67_SLICE_X162Y67_CO6;
  assign CLBLM_R_X103Y67_SLICE_X162Y67_D = CLBLM_R_X103Y67_SLICE_X162Y67_DO6;
  assign CLBLM_R_X103Y67_SLICE_X163Y67_A = CLBLM_R_X103Y67_SLICE_X163Y67_AO6;
  assign CLBLM_R_X103Y67_SLICE_X163Y67_B = CLBLM_R_X103Y67_SLICE_X163Y67_BO6;
  assign CLBLM_R_X103Y67_SLICE_X163Y67_C = CLBLM_R_X103Y67_SLICE_X163Y67_CO6;
  assign CLBLM_R_X103Y67_SLICE_X163Y67_D = CLBLM_R_X103Y67_SLICE_X163Y67_DO6;
  assign CLBLM_R_X103Y69_SLICE_X162Y69_A = CLBLM_R_X103Y69_SLICE_X162Y69_AO6;
  assign CLBLM_R_X103Y69_SLICE_X162Y69_B = CLBLM_R_X103Y69_SLICE_X162Y69_BO6;
  assign CLBLM_R_X103Y69_SLICE_X162Y69_C = CLBLM_R_X103Y69_SLICE_X162Y69_CO6;
  assign CLBLM_R_X103Y69_SLICE_X162Y69_D = CLBLM_R_X103Y69_SLICE_X162Y69_DO6;
  assign CLBLM_R_X103Y69_SLICE_X162Y69_AMUX = CLBLM_R_X103Y69_SLICE_X162Y69_A5Q;
  assign CLBLM_R_X103Y69_SLICE_X163Y69_A = CLBLM_R_X103Y69_SLICE_X163Y69_AO6;
  assign CLBLM_R_X103Y69_SLICE_X163Y69_B = CLBLM_R_X103Y69_SLICE_X163Y69_BO6;
  assign CLBLM_R_X103Y69_SLICE_X163Y69_C = CLBLM_R_X103Y69_SLICE_X163Y69_CO6;
  assign CLBLM_R_X103Y69_SLICE_X163Y69_D = CLBLM_R_X103Y69_SLICE_X163Y69_DO6;
  assign CLBLM_R_X103Y75_SLICE_X162Y75_A = CLBLM_R_X103Y75_SLICE_X162Y75_AO6;
  assign CLBLM_R_X103Y75_SLICE_X162Y75_B = CLBLM_R_X103Y75_SLICE_X162Y75_BO6;
  assign CLBLM_R_X103Y75_SLICE_X162Y75_C = CLBLM_R_X103Y75_SLICE_X162Y75_CO6;
  assign CLBLM_R_X103Y75_SLICE_X162Y75_D = CLBLM_R_X103Y75_SLICE_X162Y75_DO6;
  assign CLBLM_R_X103Y75_SLICE_X163Y75_A = CLBLM_R_X103Y75_SLICE_X163Y75_AO6;
  assign CLBLM_R_X103Y75_SLICE_X163Y75_B = CLBLM_R_X103Y75_SLICE_X163Y75_BO6;
  assign CLBLM_R_X103Y75_SLICE_X163Y75_C = CLBLM_R_X103Y75_SLICE_X163Y75_CO6;
  assign CLBLM_R_X103Y75_SLICE_X163Y75_D = CLBLM_R_X103Y75_SLICE_X163Y75_DO6;
  assign CLBLM_R_X103Y76_SLICE_X162Y76_A = CLBLM_R_X103Y76_SLICE_X162Y76_AO6;
  assign CLBLM_R_X103Y76_SLICE_X162Y76_B = CLBLM_R_X103Y76_SLICE_X162Y76_BO6;
  assign CLBLM_R_X103Y76_SLICE_X162Y76_C = CLBLM_R_X103Y76_SLICE_X162Y76_CO6;
  assign CLBLM_R_X103Y76_SLICE_X162Y76_D = CLBLM_R_X103Y76_SLICE_X162Y76_DO6;
  assign CLBLM_R_X103Y76_SLICE_X163Y76_A = CLBLM_R_X103Y76_SLICE_X163Y76_AO6;
  assign CLBLM_R_X103Y76_SLICE_X163Y76_B = CLBLM_R_X103Y76_SLICE_X163Y76_BO6;
  assign CLBLM_R_X103Y76_SLICE_X163Y76_C = CLBLM_R_X103Y76_SLICE_X163Y76_CO6;
  assign CLBLM_R_X103Y76_SLICE_X163Y76_D = CLBLM_R_X103Y76_SLICE_X163Y76_DO6;
  assign LIOI3_X0Y51_OLOGIC_X0Y52_OQ = CLBLM_L_X68Y95_SLICE_X102Y95_A5Q;
  assign LIOI3_X0Y51_OLOGIC_X0Y52_TQ = 1'b1;
  assign LIOI3_X0Y51_OLOGIC_X0Y51_OQ = CLBLM_L_X62Y101_SLICE_X92Y101_AQ;
  assign LIOI3_X0Y51_OLOGIC_X0Y51_TQ = 1'b1;
  assign LIOI3_X0Y53_OLOGIC_X0Y54_OQ = CLBLM_L_X62Y92_SLICE_X92Y92_AQ;
  assign LIOI3_X0Y53_OLOGIC_X0Y54_TQ = 1'b1;
  assign LIOI3_X0Y53_OLOGIC_X0Y53_OQ = CLBLM_L_X62Y90_SLICE_X92Y90_AQ;
  assign LIOI3_X0Y53_OLOGIC_X0Y53_TQ = 1'b1;
  assign LIOI3_X0Y55_OLOGIC_X0Y56_OQ = CLBLM_L_X62Y92_SLICE_X92Y92_BQ;
  assign LIOI3_X0Y55_OLOGIC_X0Y56_TQ = 1'b1;
  assign LIOI3_X0Y55_OLOGIC_X0Y55_OQ = CLBLM_L_X60Y97_SLICE_X91Y97_AQ;
  assign LIOI3_X0Y55_OLOGIC_X0Y55_TQ = 1'b1;
  assign LIOI3_X0Y59_OLOGIC_X0Y60_OQ = CLBLM_L_X72Y106_SLICE_X108Y106_A5Q;
  assign LIOI3_X0Y59_OLOGIC_X0Y60_TQ = 1'b1;
  assign LIOI3_X0Y59_OLOGIC_X0Y59_OQ = CLBLM_L_X60Y101_SLICE_X90Y101_AQ;
  assign LIOI3_X0Y59_OLOGIC_X0Y59_TQ = 1'b1;
  assign LIOI3_X0Y61_OLOGIC_X0Y62_OQ = CLBLM_R_X65Y110_SLICE_X99Y110_B5Q;
  assign LIOI3_X0Y61_OLOGIC_X0Y62_TQ = 1'b1;
  assign LIOI3_X0Y61_OLOGIC_X0Y61_OQ = CLBLM_R_X65Y109_SLICE_X98Y109_A5Q;
  assign LIOI3_X0Y61_OLOGIC_X0Y61_TQ = 1'b1;
  assign LIOI3_X0Y65_OLOGIC_X0Y66_OQ = CLBLM_R_X65Y110_SLICE_X98Y110_A5Q;
  assign LIOI3_X0Y65_OLOGIC_X0Y66_TQ = 1'b1;
  assign LIOI3_X0Y65_OLOGIC_X0Y65_OQ = CLBLM_L_X72Y107_SLICE_X109Y107_BQ;
  assign LIOI3_X0Y65_OLOGIC_X0Y65_TQ = 1'b1;
  assign LIOI3_X0Y67_OLOGIC_X0Y68_OQ = CLBLL_R_X71Y134_SLICE_X106Y134_AQ;
  assign LIOI3_X0Y67_OLOGIC_X0Y68_TQ = 1'b1;
  assign LIOI3_X0Y67_OLOGIC_X0Y67_OQ = CLBLM_L_X72Y103_SLICE_X109Y103_AQ;
  assign LIOI3_X0Y67_OLOGIC_X0Y67_TQ = 1'b1;
  assign LIOI3_X0Y71_OLOGIC_X0Y72_OQ = CLBLM_L_X60Y104_SLICE_X90Y104_AQ;
  assign LIOI3_X0Y71_OLOGIC_X0Y72_TQ = 1'b1;
  assign LIOI3_X0Y71_OLOGIC_X0Y71_OQ = CLBLM_L_X60Y94_SLICE_X90Y94_AQ;
  assign LIOI3_X0Y71_OLOGIC_X0Y71_TQ = 1'b1;
  assign LIOI3_X0Y73_OLOGIC_X0Y74_OQ = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign LIOI3_X0Y73_OLOGIC_X0Y74_TQ = 1'b1;
  assign LIOI3_X0Y73_OLOGIC_X0Y73_OQ = CLBLM_L_X62Y105_SLICE_X93Y105_A5Q;
  assign LIOI3_X0Y73_OLOGIC_X0Y73_TQ = 1'b1;
  assign LIOI3_X0Y75_OLOGIC_X0Y76_OQ = CLBLM_L_X60Y99_SLICE_X90Y99_AQ;
  assign LIOI3_X0Y75_OLOGIC_X0Y76_TQ = 1'b1;
  assign LIOI3_X0Y75_OLOGIC_X0Y75_OQ = CLBLM_L_X60Y101_SLICE_X90Y101_BQ;
  assign LIOI3_X0Y75_OLOGIC_X0Y75_TQ = 1'b1;
  assign LIOI3_X0Y77_OLOGIC_X0Y78_OQ = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign LIOI3_X0Y77_OLOGIC_X0Y78_TQ = 1'b1;
  assign LIOI3_X0Y77_OLOGIC_X0Y77_OQ = CLBLM_L_X60Y97_SLICE_X90Y97_BQ;
  assign LIOI3_X0Y77_OLOGIC_X0Y77_TQ = 1'b1;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_OQ = CLBLM_L_X60Y92_SLICE_X90Y92_BQ;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_TQ = 1'b1;
  assign LIOI3_X0Y79_OLOGIC_X0Y79_OQ = CLBLM_L_X64Y106_SLICE_X96Y106_A5Q;
  assign LIOI3_X0Y79_OLOGIC_X0Y79_TQ = 1'b1;
  assign LIOI3_X0Y83_OLOGIC_X0Y84_OQ = CLBLM_L_X60Y99_SLICE_X90Y99_CQ;
  assign LIOI3_X0Y83_OLOGIC_X0Y84_TQ = 1'b1;
  assign LIOI3_X0Y83_OLOGIC_X0Y83_OQ = CLBLM_L_X70Y99_SLICE_X104Y99_AQ;
  assign LIOI3_X0Y83_OLOGIC_X0Y83_TQ = 1'b1;
  assign LIOI3_X0Y85_OLOGIC_X0Y86_OQ = CLBLM_L_X70Y100_SLICE_X105Y100_CQ;
  assign LIOI3_X0Y85_OLOGIC_X0Y86_TQ = 1'b1;
  assign LIOI3_X0Y85_OLOGIC_X0Y85_OQ = CLBLM_L_X60Y94_SLICE_X90Y94_BQ;
  assign LIOI3_X0Y85_OLOGIC_X0Y85_TQ = 1'b1;
  assign LIOI3_X0Y89_OLOGIC_X0Y90_OQ = CLBLM_R_X63Y103_SLICE_X94Y103_AQ;
  assign LIOI3_X0Y89_OLOGIC_X0Y90_TQ = 1'b1;
  assign LIOI3_X0Y89_OLOGIC_X0Y89_OQ = CLBLM_R_X63Y98_SLICE_X94Y98_BQ;
  assign LIOI3_X0Y89_OLOGIC_X0Y89_TQ = 1'b1;
  assign LIOI3_X0Y91_OLOGIC_X0Y92_OQ = CLBLM_L_X62Y95_SLICE_X92Y95_CQ;
  assign LIOI3_X0Y91_OLOGIC_X0Y92_TQ = 1'b1;
  assign LIOI3_X0Y91_OLOGIC_X0Y91_OQ = CLBLM_L_X60Y99_SLICE_X90Y99_DQ;
  assign LIOI3_X0Y91_OLOGIC_X0Y91_TQ = 1'b1;
  assign LIOI3_X0Y95_OLOGIC_X0Y96_OQ = CLBLM_R_X63Y97_SLICE_X95Y97_AQ;
  assign LIOI3_X0Y95_OLOGIC_X0Y96_TQ = 1'b1;
  assign LIOI3_X0Y95_OLOGIC_X0Y95_OQ = CLBLM_L_X70Y101_SLICE_X104Y101_AQ;
  assign LIOI3_X0Y95_OLOGIC_X0Y95_TQ = 1'b1;
  assign LIOI3_X0Y97_OLOGIC_X0Y98_OQ = CLBLM_L_X68Y97_SLICE_X103Y97_AQ;
  assign LIOI3_X0Y97_OLOGIC_X0Y98_TQ = 1'b1;
  assign LIOI3_X0Y97_OLOGIC_X0Y97_OQ = CLBLM_L_X62Y103_SLICE_X92Y103_A5Q;
  assign LIOI3_X0Y97_OLOGIC_X0Y97_TQ = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_OQ = RIOB33_X105Y59_IOB_X1Y59_I;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_TQ = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_OQ = RIOB33_X105Y57_IOB_X1Y58_I;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_OQ = RIOB33_X105Y53_IOB_X1Y53_I;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_OQ = RIOB33_X105Y55_IOB_X1Y56_I;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_OQ = RIOB33_X105Y59_IOB_X1Y60_I;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_OQ = RIOB33_X105Y53_IOB_X1Y54_I;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_OQ = CLBLL_R_X77Y129_SLICE_X118Y129_AQ;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_OQ = CLBLL_R_X75Y133_SLICE_X114Y133_AQ;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_OQ = CLBLM_L_X64Y99_SLICE_X97Y99_B5Q;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_OQ = CLBLM_R_X65Y106_SLICE_X99Y106_DQ;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_OQ = CLBLM_L_X76Y118_SLICE_X117Y118_CQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_OQ = CLBLM_R_X67Y118_SLICE_X100Y118_A5Q;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_OQ = CLBLM_R_X67Y116_SLICE_X100Y116_AQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_OQ = CLBLM_L_X76Y125_SLICE_X116Y125_AQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_OQ = RIOB33_X105Y51_IOB_X1Y52_I;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_OQ = CLBLL_R_X73Y123_SLICE_X110Y123_AQ;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_OQ = CLBLL_L_X34Y123_SLICE_X50Y123_AO6;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_OQ = CLBLM_R_X67Y108_SLICE_X100Y108_AO6;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_OQ = CLBLL_L_X2Y131_SLICE_X0Y131_AO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_OQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_OQ = CLBLL_R_X73Y131_SLICE_X110Y131_AQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_OQ = CLBLL_L_X34Y126_SLICE_X50Y126_AO6;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_OQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_OQ = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_OQ = CLBLM_L_X70Y135_SLICE_X104Y135_CO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_OQ = CLBLM_R_X63Y105_SLICE_X95Y105_A5Q;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_OQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_OQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_OQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_OQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_OQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_OQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_OQ = CLBLM_L_X72Y123_SLICE_X108Y123_BO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_OQ = CLBLL_R_X71Y130_SLICE_X106Y130_DO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_OQ = CLBLL_R_X73Y134_SLICE_X110Y134_AO5;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_OQ = CLBLL_R_X71Y124_SLICE_X106Y124_BO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_OQ = CLBLM_L_X64Y105_SLICE_X97Y105_DO6;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_OQ = CLBLM_L_X72Y128_SLICE_X109Y128_AO6;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_TQ = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_OQ = CLBLM_R_X67Y118_SLICE_X100Y118_A5Q;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_TQ = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_OQ = CLBLM_R_X65Y106_SLICE_X99Y106_DQ;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_TQ = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_OQ = CLBLM_L_X64Y99_SLICE_X97Y99_B5Q;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_TQ = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_OQ = CLBLM_L_X76Y118_SLICE_X117Y118_CQ;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_TQ = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_OQ = CLBLL_R_X71Y119_SLICE_X106Y119_AQ;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_TQ = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_OQ = CLBLM_R_X67Y116_SLICE_X100Y116_AQ;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_TQ = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_OQ = CLBLL_R_X71Y124_SLICE_X106Y124_AQ;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_TQ = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_OQ = CLBLM_L_X70Y110_SLICE_X104Y110_CQ;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_TQ = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_OQ = CLBLL_L_X2Y131_SLICE_X0Y131_AO6;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_TQ = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_OQ = CLBLL_L_X34Y123_SLICE_X50Y123_AO6;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_TQ = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_OQ = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_TQ = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_OQ = CLBLL_L_X34Y126_SLICE_X50Y126_AO6;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_TQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_OQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_TQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_OQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_TQ = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_OQ = CLBLM_L_X62Y107_SLICE_X92Y107_AO5;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_TQ = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_OQ = CLBLM_L_X68Y107_SLICE_X102Y107_BO6;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_TQ = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_OQ = CLBLM_L_X70Y135_SLICE_X104Y135_CO6;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_TQ = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_OQ = CLBLM_R_X63Y105_SLICE_X95Y105_A5Q;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_TQ = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_OQ = CLBLM_L_X72Y122_SLICE_X108Y122_AO6;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_TQ = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_OQ = CLBLM_L_X70Y134_SLICE_X104Y134_CO5;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_OQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_OQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_OQ = CLBLL_R_X73Y134_SLICE_X110Y134_AO5;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_OQ = CLBLM_L_X70Y125_SLICE_X104Y125_DO6;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_OQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_OQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_OQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_OQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_OQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_OQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_OQ = CLBLM_L_X64Y105_SLICE_X97Y105_DO6;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_OQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_OQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_OQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_TQ = 1'b1;
  assign LIOI3_SING_X0Y50_OLOGIC_X0Y50_OQ = CLBLM_L_X60Y97_SLICE_X90Y97_DQ;
  assign LIOI3_SING_X0Y50_OLOGIC_X0Y50_TQ = 1'b1;
  assign LIOI3_SING_X0Y99_OLOGIC_X0Y99_OQ = RIOB33_X105Y61_IOB_X1Y62_I;
  assign LIOI3_SING_X0Y99_OLOGIC_X0Y99_TQ = 1'b1;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ = RIOB33_X105Y57_IOB_X1Y57_I;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ = 1'b1;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ = CLBLM_R_X67Y105_SLICE_X101Y105_AO6;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ = 1'b1;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ = CLBLM_L_X74Y129_SLICE_X113Y129_BO6;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ = 1'b1;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ = 1'b1;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y58_OQ = CLBLM_L_X72Y107_SLICE_X108Y107_BQ;
  assign LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y58_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y57_OQ = CLBLM_L_X62Y95_SLICE_X92Y95_AQ;
  assign LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y57_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y69_OLOGIC_X0Y70_OQ = CLBLL_R_X75Y127_SLICE_X115Y127_AQ;
  assign LIOI3_TBYTESRC_X0Y69_OLOGIC_X0Y70_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y69_OLOGIC_X0Y69_OQ = CLBLM_L_X60Y92_SLICE_X90Y92_AQ;
  assign LIOI3_TBYTESRC_X0Y69_OLOGIC_X0Y69_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y81_OLOGIC_X0Y82_OQ = CLBLM_L_X62Y107_SLICE_X93Y107_A5Q;
  assign LIOI3_TBYTESRC_X0Y81_OLOGIC_X0Y82_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y81_OLOGIC_X0Y81_OQ = CLBLM_L_X60Y99_SLICE_X90Y99_BQ;
  assign LIOI3_TBYTESRC_X0Y81_OLOGIC_X0Y81_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y94_OQ = CLBLM_L_X62Y106_SLICE_X92Y106_AQ;
  assign LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y94_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y93_OQ = CLBLM_L_X62Y95_SLICE_X92Y95_BQ;
  assign LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y93_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ = CLBLM_L_X70Y110_SLICE_X104Y110_CQ;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ = RIOB33_X105Y55_IOB_X1Y55_I;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ = CLBLL_R_X71Y119_SLICE_X106Y119_AQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ = CLBLM_R_X63Y106_SLICE_X95Y106_AQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ = CLBLM_L_X70Y134_SLICE_X104Y134_CO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ = CLBLM_L_X62Y107_SLICE_X92Y107_AO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ = CLBLM_L_X64Y106_SLICE_X97Y106_AO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_OQ = CLBLM_L_X76Y125_SLICE_X116Y125_AQ;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_OQ = CLBLM_R_X63Y122_SLICE_X95Y122_CQ;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_OQ = CLBLM_L_X74Y120_SLICE_X112Y120_AO6;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_OQ = CLBLL_R_X73Y131_SLICE_X110Y131_AQ;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ = CLBLM_L_X70Y126_SLICE_X104Y126_DO6;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ = CLBLM_L_X64Y106_SLICE_X97Y106_AO6;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_OQ = CLBLL_R_X73Y103_SLICE_X111Y103_A5Q;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y63_OQ = CLBLL_R_X73Y102_SLICE_X111Y102_A5Q;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y63_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y88_OQ = CLBLM_L_X60Y94_SLICE_X90Y94_CQ;
  assign LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y88_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y87_OQ = CLBLM_R_X63Y97_SLICE_X94Y97_B5Q;
  assign LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y87_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ = CLBLL_R_X71Y124_SLICE_X106Y124_AQ;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ = CLBLM_R_X63Y122_SLICE_X95Y122_CQ;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_OQ = CLBLL_R_X73Y123_SLICE_X110Y123_AQ;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_OQ = CLBLM_R_X63Y106_SLICE_X95Y106_AQ;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ = CLBLL_R_X77Y124_SLICE_X118Y124_AO6;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ = 1'b1;
  assign RIOI3_X105Y51_ILOGIC_X1Y52_O = RIOB33_X105Y51_IOB_X1Y52_I;
  assign RIOI3_X105Y51_ILOGIC_X1Y51_O = RIOB33_X105Y51_IOB_X1Y51_I;
  assign RIOI3_X105Y53_ILOGIC_X1Y54_O = RIOB33_X105Y53_IOB_X1Y54_I;
  assign RIOI3_X105Y53_ILOGIC_X1Y53_O = RIOB33_X105Y53_IOB_X1Y53_I;
  assign RIOI3_X105Y55_ILOGIC_X1Y56_O = RIOB33_X105Y55_IOB_X1Y56_I;
  assign RIOI3_X105Y55_ILOGIC_X1Y55_O = RIOB33_X105Y55_IOB_X1Y55_I;
  assign RIOI3_X105Y59_ILOGIC_X1Y60_O = RIOB33_X105Y59_IOB_X1Y60_I;
  assign RIOI3_X105Y59_ILOGIC_X1Y59_O = RIOB33_X105Y59_IOB_X1Y59_I;
  assign RIOI3_X105Y61_ILOGIC_X1Y62_O = RIOB33_X105Y61_IOB_X1Y62_I;
  assign RIOI3_X105Y65_OLOGIC_X1Y66_OQ = CLBLM_R_X103Y67_SLICE_X162Y67_CQ;
  assign RIOI3_X105Y65_OLOGIC_X1Y66_TQ = 1'b1;
  assign RIOI3_X105Y65_OLOGIC_X1Y65_OQ = CLBLM_R_X103Y67_SLICE_X162Y67_BQ;
  assign RIOI3_X105Y65_OLOGIC_X1Y65_TQ = 1'b1;
  assign RIOI3_X105Y67_OLOGIC_X1Y68_OQ = CLBLM_R_X103Y67_SLICE_X163Y67_CQ;
  assign RIOI3_X105Y67_OLOGIC_X1Y68_TQ = 1'b1;
  assign RIOI3_X105Y67_OLOGIC_X1Y67_OQ = CLBLM_R_X103Y67_SLICE_X163Y67_BQ;
  assign RIOI3_X105Y67_OLOGIC_X1Y67_TQ = 1'b1;
  assign RIOI3_X105Y71_OLOGIC_X1Y72_OQ = CLBLM_R_X103Y76_SLICE_X162Y76_AQ;
  assign RIOI3_X105Y71_OLOGIC_X1Y72_TQ = 1'b1;
  assign RIOI3_X105Y71_OLOGIC_X1Y71_OQ = CLBLM_R_X103Y75_SLICE_X162Y75_BQ;
  assign RIOI3_X105Y71_OLOGIC_X1Y71_TQ = 1'b1;
  assign RIOI3_X105Y73_OLOGIC_X1Y74_OQ = CLBLM_R_X103Y75_SLICE_X162Y75_AQ;
  assign RIOI3_X105Y73_OLOGIC_X1Y74_TQ = 1'b1;
  assign RIOI3_X105Y73_OLOGIC_X1Y73_OQ = CLBLM_R_X103Y75_SLICE_X163Y75_AQ;
  assign RIOI3_X105Y73_OLOGIC_X1Y73_TQ = 1'b1;
  assign RIOI3_X105Y75_OLOGIC_X1Y76_OQ = CLBLM_R_X103Y75_SLICE_X163Y75_BQ;
  assign RIOI3_X105Y75_OLOGIC_X1Y76_TQ = 1'b1;
  assign RIOI3_X105Y75_OLOGIC_X1Y75_OQ = CLBLM_R_X103Y75_SLICE_X162Y75_CQ;
  assign RIOI3_X105Y75_OLOGIC_X1Y75_TQ = 1'b1;
  assign RIOI3_X105Y77_ILOGIC_X1Y78_O = RIOB33_X105Y77_IOB_X1Y78_I;
  assign RIOI3_X105Y77_OLOGIC_X1Y77_OQ = CLBLM_R_X103Y76_SLICE_X163Y76_AQ;
  assign RIOI3_X105Y77_OLOGIC_X1Y77_TQ = 1'b1;
  assign RIOI3_X105Y79_OLOGIC_X1Y80_OQ = 1'b0;
  assign RIOI3_X105Y79_OLOGIC_X1Y80_TQ = 1'b1;
  assign RIOI3_X105Y79_OLOGIC_X1Y79_OQ = CLBLL_R_X83Y94_SLICE_X130Y94_A5Q;
  assign RIOI3_X105Y79_OLOGIC_X1Y79_TQ = 1'b1;
  assign RIOI3_X105Y83_OLOGIC_X1Y84_OQ = CLBLM_L_X72Y118_SLICE_X108Y118_D5Q;
  assign RIOI3_X105Y83_OLOGIC_X1Y84_TQ = 1'b1;
  assign RIOI3_X105Y83_OLOGIC_X1Y83_OQ = CLBLM_R_X63Y105_SLICE_X95Y105_AQ;
  assign RIOI3_X105Y83_OLOGIC_X1Y83_TQ = 1'b1;
  assign RIOI3_X105Y85_OLOGIC_X1Y86_OQ = CLBLM_L_X64Y99_SLICE_X97Y99_A5Q;
  assign RIOI3_X105Y85_OLOGIC_X1Y86_TQ = 1'b1;
  assign RIOI3_X105Y85_OLOGIC_X1Y85_OQ = CLBLL_R_X71Y98_SLICE_X106Y98_AQ;
  assign RIOI3_X105Y85_OLOGIC_X1Y85_TQ = 1'b1;
  assign RIOI3_X105Y89_OLOGIC_X1Y90_OQ = CLBLM_L_X72Y119_SLICE_X108Y119_C5Q;
  assign RIOI3_X105Y89_OLOGIC_X1Y90_TQ = 1'b1;
  assign RIOI3_X105Y89_OLOGIC_X1Y89_OQ = CLBLM_L_X64Y101_SLICE_X96Y101_AQ;
  assign RIOI3_X105Y89_OLOGIC_X1Y89_TQ = 1'b1;
  assign RIOI3_X105Y91_OLOGIC_X1Y91_OQ = CLBLM_L_X68Y98_SLICE_X103Y98_AQ;
  assign RIOI3_X105Y91_OLOGIC_X1Y91_TQ = 1'b1;
  assign RIOI3_X105Y101_OLOGIC_X1Y102_OQ = CLBLL_R_X73Y131_SLICE_X111Y131_AQ;
  assign RIOI3_X105Y101_OLOGIC_X1Y102_TQ = 1'b1;
  assign RIOI3_X105Y101_OLOGIC_X1Y101_OQ = CLBLM_L_X72Y109_SLICE_X109Y109_DQ;
  assign RIOI3_X105Y101_OLOGIC_X1Y101_TQ = 1'b1;
  assign RIOI3_X105Y103_OLOGIC_X1Y104_OQ = CLBLM_L_X72Y106_SLICE_X108Y106_AQ;
  assign RIOI3_X105Y103_OLOGIC_X1Y104_TQ = 1'b1;
  assign RIOI3_X105Y103_OLOGIC_X1Y103_OQ = CLBLL_R_X77Y128_SLICE_X119Y128_DQ;
  assign RIOI3_X105Y103_OLOGIC_X1Y103_TQ = 1'b1;
  assign RIOI3_X105Y105_OLOGIC_X1Y106_OQ = CLBLL_R_X75Y103_SLICE_X115Y103_AQ;
  assign RIOI3_X105Y105_OLOGIC_X1Y106_TQ = 1'b1;
  assign RIOI3_X105Y105_OLOGIC_X1Y105_OQ = CLBLM_R_X65Y111_SLICE_X98Y111_AQ;
  assign RIOI3_X105Y105_OLOGIC_X1Y105_TQ = 1'b1;
  assign RIOI3_X105Y109_OLOGIC_X1Y110_OQ = CLBLM_L_X72Y111_SLICE_X108Y111_C5Q;
  assign RIOI3_X105Y109_OLOGIC_X1Y110_TQ = 1'b1;
  assign RIOI3_X105Y109_OLOGIC_X1Y109_OQ = CLBLL_R_X79Y104_SLICE_X122Y104_AQ;
  assign RIOI3_X105Y109_OLOGIC_X1Y109_TQ = 1'b1;
  assign RIOI3_X105Y111_OLOGIC_X1Y112_OQ = CLBLL_R_X71Y100_SLICE_X106Y100_BQ;
  assign RIOI3_X105Y111_OLOGIC_X1Y112_TQ = 1'b1;
  assign RIOI3_X105Y111_OLOGIC_X1Y111_OQ = CLBLM_L_X62Y107_SLICE_X93Y107_BQ;
  assign RIOI3_X105Y111_OLOGIC_X1Y111_TQ = 1'b1;
  assign RIOI3_X105Y115_OLOGIC_X1Y116_OQ = CLBLM_L_X68Y95_SLICE_X102Y95_AQ;
  assign RIOI3_X105Y115_OLOGIC_X1Y116_TQ = 1'b1;
  assign RIOI3_X105Y115_OLOGIC_X1Y115_OQ = CLBLM_L_X62Y100_SLICE_X92Y100_AQ;
  assign RIOI3_X105Y115_OLOGIC_X1Y115_TQ = 1'b1;
  assign RIOI3_X105Y117_OLOGIC_X1Y118_OQ = CLBLM_L_X70Y136_SLICE_X105Y136_A5Q;
  assign RIOI3_X105Y117_OLOGIC_X1Y118_TQ = 1'b1;
  assign RIOI3_X105Y117_OLOGIC_X1Y117_OQ = CLBLL_R_X73Y118_SLICE_X111Y118_AQ;
  assign RIOI3_X105Y117_OLOGIC_X1Y117_TQ = 1'b1;
  assign RIOI3_X105Y121_OLOGIC_X1Y122_OQ = CLBLM_R_X63Y98_SLICE_X94Y98_AQ;
  assign RIOI3_X105Y121_OLOGIC_X1Y122_TQ = 1'b1;
  assign RIOI3_X105Y121_OLOGIC_X1Y121_OQ = CLBLM_L_X70Y100_SLICE_X104Y100_A5Q;
  assign RIOI3_X105Y121_OLOGIC_X1Y121_TQ = 1'b1;
  assign RIOI3_X105Y123_OLOGIC_X1Y124_OQ = CLBLM_L_X68Y99_SLICE_X102Y99_AQ;
  assign RIOI3_X105Y123_OLOGIC_X1Y124_TQ = 1'b1;
  assign RIOI3_X105Y123_OLOGIC_X1Y123_OQ = CLBLM_R_X63Y101_SLICE_X94Y101_AQ;
  assign RIOI3_X105Y123_OLOGIC_X1Y123_TQ = 1'b1;
  assign RIOI3_X105Y125_OLOGIC_X1Y126_OQ = CLBLM_L_X76Y127_SLICE_X116Y127_AQ;
  assign RIOI3_X105Y125_OLOGIC_X1Y126_TQ = 1'b1;
  assign RIOI3_X105Y125_OLOGIC_X1Y125_OQ = CLBLM_L_X74Y129_SLICE_X112Y129_BQ;
  assign RIOI3_X105Y125_OLOGIC_X1Y125_TQ = 1'b1;
  assign RIOI3_X105Y127_OLOGIC_X1Y128_OQ = CLBLM_R_X65Y110_SLICE_X99Y110_CQ;
  assign RIOI3_X105Y127_OLOGIC_X1Y128_TQ = 1'b1;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_OQ = CLBLM_L_X72Y107_SLICE_X108Y107_A5Q;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_TQ = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_OQ = CLBLL_R_X73Y103_SLICE_X110Y103_B5Q;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_TQ = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_OQ = CLBLM_L_X78Y106_SLICE_X120Y106_AQ;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_TQ = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_OQ = CLBLL_R_X83Y130_SLICE_X130Y130_BQ;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_TQ = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_OQ = CLBLL_R_X83Y130_SLICE_X130Y130_AQ;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_TQ = 1'b1;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_OQ = CLBLL_R_X83Y130_SLICE_X130Y130_DQ;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_TQ = 1'b1;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_OQ = CLBLL_R_X83Y130_SLICE_X130Y130_CQ;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_TQ = 1'b1;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_OQ = CLBLM_L_X72Y107_SLICE_X109Y107_A5Q;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_TQ = 1'b1;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_OQ = CLBLL_R_X83Y132_SLICE_X130Y132_AQ;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_TQ = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_OQ = CLBLL_R_X73Y103_SLICE_X110Y103_A5Q;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_TQ = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_OQ = CLBLM_R_X65Y110_SLICE_X99Y110_AQ;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_TQ = 1'b1;
  assign RIOI3_X105Y145_OLOGIC_X1Y146_OQ = CLBLM_R_X63Y97_SLICE_X94Y97_AQ;
  assign RIOI3_X105Y145_OLOGIC_X1Y146_TQ = 1'b1;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_OQ = CLBLL_R_X75Y107_SLICE_X114Y107_AQ;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_TQ = 1'b1;
  assign RIOI3_X105Y147_OLOGIC_X1Y148_OQ = CLBLM_L_X62Y103_SLICE_X92Y103_B5Q;
  assign RIOI3_X105Y147_OLOGIC_X1Y148_TQ = 1'b1;
  assign RIOI3_X105Y147_OLOGIC_X1Y147_OQ = CLBLL_R_X77Y108_SLICE_X118Y108_AQ;
  assign RIOI3_X105Y147_OLOGIC_X1Y147_TQ = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_OQ = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_TQ = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_OQ = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_OQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_OQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_OQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_OQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_OQ = CLBLM_L_X74Y120_SLICE_X112Y120_AO6;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_OQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_OQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_OQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_OQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_OQ = CLBLM_L_X70Y111_SLICE_X105Y111_DO6;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_OQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_OQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_OQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_OQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_OQ = CLBLM_L_X70Y111_SLICE_X105Y111_DO6;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_OQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_OQ = CLBLL_R_X73Y119_SLICE_X110Y119_AQ;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_OQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_OQ = CLBLL_R_X73Y119_SLICE_X110Y119_BQ;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_OQ = CLBLM_L_X72Y119_SLICE_X109Y119_BQ;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_OQ = CLBLM_R_X67Y118_SLICE_X101Y118_AQ;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_OQ = CLBLM_L_X72Y119_SLICE_X108Y119_CQ;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_OQ = 1'b0;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_OQ = 1'b0;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_OQ = 1'b0;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_OQ = CLBLL_R_X71Y117_SLICE_X106Y117_A5Q;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_OQ = CLBLM_L_X76Y128_SLICE_X116Y128_C5Q;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_OQ = 1'b0;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_OQ = CLBLM_L_X72Y118_SLICE_X109Y118_A5Q;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_OQ = CLBLM_L_X68Y109_SLICE_X102Y109_AQ;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_OQ = 1'b0;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_OQ = CLBLL_R_X73Y104_SLICE_X110Y104_AQ;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_OQ = CLBLM_L_X80Y132_SLICE_X124Y132_AQ;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_OQ = CLBLL_R_X79Y135_SLICE_X122Y135_AQ;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_TQ = 1'b1;
  assign RIOI3_SING_X105Y50_ILOGIC_X1Y50_O = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign RIOI3_SING_X105Y100_OLOGIC_X1Y100_OQ = CLBLM_L_X78Y104_SLICE_X120Y104_A5Q;
  assign RIOI3_SING_X105Y100_OLOGIC_X1Y100_TQ = 1'b1;
  assign RIOI3_SING_X105Y149_OLOGIC_X1Y149_OQ = CLBLM_L_X76Y111_SLICE_X116Y111_BQ;
  assign RIOI3_SING_X105Y149_OLOGIC_X1Y149_TQ = 1'b1;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ = 1'b1;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ = 1'b1;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ = CLBLM_L_X74Y109_SLICE_X113Y109_AQ;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y57_ILOGIC_X1Y58_O = RIOB33_X105Y57_IOB_X1Y58_I;
  assign RIOI3_TBYTESRC_X105Y57_ILOGIC_X1Y57_O = RIOB33_X105Y57_IOB_X1Y57_I;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_OQ = CLBLM_L_X82Y98_SLICE_X128Y98_AQ;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_OQ = CLBLM_R_X103Y69_SLICE_X163Y69_AQ;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_OQ = CLBLL_R_X77Y104_SLICE_X119Y104_A5Q;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_OQ = CLBLL_R_X71Y110_SLICE_X106Y110_A5Q;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_OQ = CLBLL_R_X77Y113_SLICE_X118Y113_AQ;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_OQ = CLBLM_R_X103Y69_SLICE_X162Y69_AQ;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_OQ = CLBLM_L_X62Y106_SLICE_X93Y106_AQ;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_OQ = CLBLM_L_X76Y128_SLICE_X116Y128_CQ;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_OQ = CLBLL_R_X79Y104_SLICE_X122Y104_A5Q;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_OQ = CLBLM_L_X76Y111_SLICE_X116Y111_AQ;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_OQ = CLBLM_L_X70Y101_SLICE_X105Y101_AQ;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_OQ = CLBLM_L_X62Y106_SLICE_X92Y106_BQ;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ = CLBLL_R_X77Y128_SLICE_X119Y128_BQ;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ = CLBLL_R_X75Y133_SLICE_X114Y133_BQ;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ = CLBLM_L_X76Y129_SLICE_X116Y129_CQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ = 1'b0;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_OQ = CLBLM_R_X103Y67_SLICE_X163Y67_AQ;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_OQ = CLBLM_R_X103Y67_SLICE_X162Y67_AQ;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_OQ = CLBLM_L_X68Y105_SLICE_X102Y105_AQ;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_OQ = CLBLM_L_X64Y97_SLICE_X97Y97_AQ;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_OQ = 1'b0;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_OQ = CLBLM_L_X62Y99_SLICE_X93Y99_AQ;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_OQ = CLBLM_L_X82Y130_SLICE_X128Y130_AQ;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_OQ = CLBLL_R_X77Y125_SLICE_X118Y125_AQ;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ = CLBLL_R_X77Y124_SLICE_X118Y124_AO6;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ = 1'b0;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ = CLBLL_R_X71Y117_SLICE_X106Y117_B5Q;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ = CLBLL_R_X73Y108_SLICE_X110Y108_AQ;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ = 1'b1;
  assign CLBLM_R_X65Y110_SLICE_X98Y110_AX = CLBLM_R_X65Y110_SLICE_X99Y110_AQ;
  assign CLBLM_L_X76Y122_SLICE_X117Y122_A1 = 1'b1;
  assign CLBLM_L_X76Y122_SLICE_X117Y122_A2 = 1'b1;
  assign CLBLM_L_X76Y122_SLICE_X117Y122_A3 = 1'b1;
  assign CLBLM_L_X76Y122_SLICE_X117Y122_A4 = 1'b1;
  assign CLBLM_L_X76Y122_SLICE_X117Y122_A5 = 1'b1;
  assign CLBLM_L_X76Y122_SLICE_X117Y122_A6 = 1'b1;
  assign CLBLM_L_X76Y122_SLICE_X117Y122_AX = CLBLL_R_X77Y113_SLICE_X118Y113_AQ;
  assign CLBLM_L_X76Y122_SLICE_X117Y122_B1 = 1'b1;
  assign CLBLM_L_X76Y122_SLICE_X117Y122_B2 = 1'b1;
  assign CLBLM_L_X76Y122_SLICE_X117Y122_B3 = 1'b1;
  assign CLBLM_L_X76Y122_SLICE_X117Y122_B4 = 1'b1;
  assign CLBLM_L_X76Y122_SLICE_X117Y122_B5 = 1'b1;
  assign CLBLM_L_X76Y122_SLICE_X117Y122_B6 = 1'b1;
  assign CLBLM_R_X65Y110_SLICE_X98Y110_B2 = CLBLM_R_X65Y110_SLICE_X98Y110_BQ;
  assign CLBLM_R_X65Y110_SLICE_X98Y110_B3 = CLBLM_R_X67Y111_SLICE_X101Y111_CO6;
  assign LIOB33_X0Y79_IOB_X0Y79_O = CLBLM_L_X64Y106_SLICE_X96Y106_A5Q;
  assign CLBLM_L_X74Y135_SLICE_X112Y135_D1 = 1'b1;
  assign CLBLM_L_X76Y122_SLICE_X117Y122_C1 = 1'b1;
  assign CLBLM_L_X76Y122_SLICE_X117Y122_C2 = 1'b1;
  assign CLBLM_L_X76Y122_SLICE_X117Y122_C3 = 1'b1;
  assign CLBLM_L_X76Y122_SLICE_X117Y122_C4 = 1'b1;
  assign CLBLM_L_X74Y135_SLICE_X112Y135_D2 = 1'b1;
  assign CLBLM_L_X76Y122_SLICE_X117Y122_C5 = 1'b1;
  assign CLBLM_L_X76Y122_SLICE_X117Y122_C6 = 1'b1;
  assign CLBLM_L_X76Y122_SLICE_X117Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X65Y110_SLICE_X98Y110_B4 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X74Y135_SLICE_X112Y135_D3 = 1'b1;
  assign CLBLM_R_X65Y110_SLICE_X98Y110_B5 = CLBLM_R_X65Y109_SLICE_X98Y109_BQ;
  assign CLBLM_L_X74Y135_SLICE_X112Y135_D4 = 1'b1;
  assign CLBLM_L_X76Y122_SLICE_X117Y122_D1 = 1'b1;
  assign CLBLM_L_X76Y122_SLICE_X117Y122_D2 = 1'b1;
  assign CLBLM_L_X76Y122_SLICE_X117Y122_D3 = 1'b1;
  assign CLBLM_L_X76Y122_SLICE_X117Y122_D4 = 1'b1;
  assign CLBLM_L_X70Y102_SLICE_X105Y102_A1 = CLBLM_L_X70Y103_SLICE_X104Y103_DO6;
  assign CLBLM_L_X70Y102_SLICE_X105Y102_A2 = CLBLM_L_X70Y102_SLICE_X105Y102_BQ;
  assign CLBLM_L_X70Y102_SLICE_X105Y102_A3 = CLBLM_L_X70Y102_SLICE_X105Y102_AQ;
  assign CLBLM_L_X70Y102_SLICE_X105Y102_A4 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X70Y102_SLICE_X105Y102_A5 = CLBLL_R_X71Y103_SLICE_X106Y103_BO6;
  assign CLBLM_L_X70Y102_SLICE_X105Y102_A6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y135_SLICE_X112Y135_D5 = 1'b1;
  assign CLBLM_L_X74Y135_SLICE_X112Y135_D6 = 1'b1;
  assign CLBLM_L_X76Y122_SLICE_X116Y122_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y102_SLICE_X105Y102_B1 = CLBLM_L_X70Y102_SLICE_X105Y102_CQ;
  assign CLBLM_L_X70Y102_SLICE_X105Y102_B2 = CLBLM_L_X70Y102_SLICE_X105Y102_BQ;
  assign CLBLM_L_X70Y102_SLICE_X105Y102_B3 = CLBLM_L_X70Y103_SLICE_X104Y103_C5Q;
  assign CLBLM_L_X70Y102_SLICE_X105Y102_B4 = CLBLL_R_X71Y103_SLICE_X106Y103_BO5;
  assign CLBLM_L_X70Y102_SLICE_X105Y102_B5 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X70Y102_SLICE_X105Y102_B6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X76Y122_SLICE_X116Y122_A2 = CLBLM_L_X76Y122_SLICE_X116Y122_BQ;
  assign CLBLM_L_X70Y125_SLICE_X104Y125_A3 = 1'b1;
  assign CLBLM_L_X76Y122_SLICE_X116Y122_A3 = CLBLM_L_X76Y122_SLICE_X116Y122_AQ;
  assign CLBLM_L_X70Y102_SLICE_X105Y102_C1 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X70Y102_SLICE_X105Y102_C2 = CLBLM_L_X70Y102_SLICE_X105Y102_CQ;
  assign CLBLM_L_X70Y102_SLICE_X105Y102_C3 = CLBLL_R_X71Y103_SLICE_X106Y103_BO5;
  assign CLBLM_L_X70Y102_SLICE_X105Y102_C4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y102_SLICE_X105Y102_C5 = CLBLM_L_X70Y103_SLICE_X105Y103_DO5;
  assign CLBLM_L_X70Y102_SLICE_X105Y102_C6 = CLBLL_R_X71Y102_SLICE_X106Y102_CQ;
  assign CLBLM_L_X76Y122_SLICE_X116Y122_B1 = CLBLL_R_X77Y127_SLICE_X118Y127_AQ;
  assign CLBLM_L_X70Y102_SLICE_X105Y102_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X76Y122_SLICE_X116Y122_B2 = CLBLM_L_X76Y122_SLICE_X116Y122_BQ;
  assign CLBLM_L_X74Y135_SLICE_X112Y135_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X76Y122_SLICE_X116Y122_B4 = CLBLM_L_X76Y124_SLICE_X116Y124_BQ;
  assign CLBLM_L_X76Y122_SLICE_X116Y122_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y102_SLICE_X105Y102_D1 = CLBLM_L_X70Y100_SLICE_X105Y100_AQ;
  assign CLBLM_L_X70Y102_SLICE_X105Y102_D2 = CLBLM_L_X70Y100_SLICE_X105Y100_A5Q;
  assign CLBLM_L_X70Y102_SLICE_X105Y102_D3 = CLBLM_R_X65Y103_SLICE_X99Y103_DO6;
  assign CLBLM_L_X70Y102_SLICE_X105Y102_D4 = CLBLL_R_X71Y98_SLICE_X106Y98_A5Q;
  assign CLBLM_L_X70Y102_SLICE_X105Y102_D5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y102_SLICE_X105Y102_D6 = CLBLM_L_X60Y97_SLICE_X90Y97_BQ;
  assign CLBLM_L_X76Y122_SLICE_X116Y122_C3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X76Y122_SLICE_X116Y122_C4 = CLBLM_L_X76Y125_SLICE_X116Y125_C5Q;
  assign CLBLM_L_X70Y102_SLICE_X105Y102_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X76Y122_SLICE_X116Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X76Y122_SLICE_X116Y122_D1 = 1'b1;
  assign CLBLM_L_X70Y102_SLICE_X104Y102_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y102_SLICE_X104Y102_A2 = CLBLM_L_X70Y104_SLICE_X104Y104_CO5;
  assign CLBLM_L_X70Y102_SLICE_X104Y102_A3 = CLBLM_L_X70Y102_SLICE_X104Y102_AQ;
  assign CLBLM_L_X70Y102_SLICE_X104Y102_A4 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X70Y102_SLICE_X104Y102_A5 = CLBLM_L_X70Y101_SLICE_X105Y101_BQ;
  assign CLBLM_L_X70Y102_SLICE_X104Y102_A6 = 1'b1;
  assign CLBLM_L_X76Y122_SLICE_X116Y122_D2 = 1'b1;
  assign CLBLM_L_X76Y122_SLICE_X116Y122_D3 = 1'b1;
  assign CLBLM_L_X76Y122_SLICE_X116Y122_D4 = 1'b1;
  assign CLBLM_L_X76Y122_SLICE_X116Y122_D5 = 1'b1;
  assign CLBLM_L_X70Y102_SLICE_X104Y102_B1 = 1'b1;
  assign CLBLM_L_X70Y102_SLICE_X104Y102_B2 = CLBLL_R_X71Y98_SLICE_X106Y98_A5Q;
  assign CLBLM_L_X70Y102_SLICE_X104Y102_B3 = CLBLM_L_X70Y102_SLICE_X104Y102_AQ;
  assign CLBLM_L_X70Y102_SLICE_X104Y102_B4 = CLBLM_L_X60Y97_SLICE_X90Y97_BQ;
  assign CLBLM_L_X70Y102_SLICE_X104Y102_B5 = CLBLM_L_X70Y100_SLICE_X105Y100_AQ;
  assign CLBLM_L_X70Y102_SLICE_X104Y102_B6 = CLBLM_L_X70Y100_SLICE_X105Y100_A5Q;
  assign CLBLM_L_X76Y119_SLICE_X116Y119_A5 = CLBLM_L_X76Y119_SLICE_X116Y119_A5Q;
  assign LIOI3_X0Y95_OLOGIC_X0Y96_T1 = 1'b1;
  assign CLBLM_L_X70Y125_SLICE_X104Y125_B2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_D1 = CLBLM_L_X72Y107_SLICE_X109Y107_A5Q;
  assign CLBLM_L_X70Y102_SLICE_X104Y102_C1 = 1'b1;
  assign CLBLM_L_X70Y102_SLICE_X104Y102_C2 = 1'b1;
  assign CLBLM_L_X70Y102_SLICE_X104Y102_C3 = 1'b1;
  assign CLBLM_L_X70Y102_SLICE_X104Y102_C4 = 1'b1;
  assign CLBLM_L_X70Y102_SLICE_X104Y102_C5 = 1'b1;
  assign CLBLM_L_X70Y102_SLICE_X104Y102_C6 = 1'b1;
  assign LIOI3_X0Y95_OLOGIC_X0Y95_D1 = CLBLM_L_X70Y101_SLICE_X104Y101_AQ;
  assign CLBLM_L_X70Y102_SLICE_X104Y102_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_T1 = 1'b1;
  assign CLBLM_L_X70Y102_SLICE_X104Y102_D1 = 1'b1;
  assign CLBLM_L_X70Y102_SLICE_X104Y102_D2 = 1'b1;
  assign CLBLM_L_X70Y102_SLICE_X104Y102_D3 = 1'b1;
  assign CLBLM_L_X70Y102_SLICE_X104Y102_D4 = 1'b1;
  assign CLBLM_L_X70Y102_SLICE_X104Y102_D5 = 1'b1;
  assign CLBLM_L_X70Y102_SLICE_X104Y102_D6 = 1'b1;
  assign LIOI3_X0Y95_OLOGIC_X0Y95_T1 = 1'b1;
  assign RIOB33_X105Y109_IOB_X1Y110_O = CLBLM_L_X72Y111_SLICE_X108Y111_C5Q;
  assign CLBLM_L_X70Y102_SLICE_X104Y102_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign RIOB33_X105Y109_IOB_X1Y109_O = CLBLL_R_X79Y104_SLICE_X122Y104_AQ;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_D1 = CLBLL_R_X83Y132_SLICE_X130Y132_AQ;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_T1 = 1'b1;
  assign RIOB33_SING_X105Y150_IOB_X1Y150_O = 1'b1;
  assign CLBLM_R_X67Y105_SLICE_X101Y105_C1 = CLBLM_L_X68Y103_SLICE_X102Y103_B5Q;
  assign CLBLM_R_X67Y105_SLICE_X101Y105_C2 = CLBLM_L_X72Y104_SLICE_X108Y104_CQ;
  assign CLBLM_R_X67Y105_SLICE_X101Y105_C5 = CLBLM_R_X67Y108_SLICE_X100Y108_BO5;
  assign CLBLM_R_X67Y105_SLICE_X101Y105_C6 = CLBLM_L_X72Y105_SLICE_X109Y105_B5Q;
  assign LIOB33_X0Y151_IOB_X0Y152_O = CLBLM_L_X64Y105_SLICE_X97Y105_DO6;
  assign LIOB33_X0Y151_IOB_X0Y151_O = CLBLM_L_X72Y128_SLICE_X109Y128_AO6;
  assign RIOB33_SING_X105Y199_IOB_X1Y199_O = CLBLM_L_X74Y109_SLICE_X113Y109_AQ;
  assign LIOB33_X0Y187_IOB_X0Y188_O = CLBLL_R_X77Y124_SLICE_X118Y124_AO6;
  assign CLBLM_R_X67Y105_SLICE_X101Y105_D1 = CLBLM_R_X65Y105_SLICE_X99Y105_BO6;
  assign CLBLM_L_X76Y123_SLICE_X117Y123_A1 = CLBLL_R_X75Y113_SLICE_X114Y113_AQ;
  assign CLBLM_L_X76Y123_SLICE_X117Y123_A2 = 1'b1;
  assign CLBLM_L_X76Y123_SLICE_X117Y123_A3 = CLBLM_L_X76Y123_SLICE_X117Y123_AQ;
  assign CLBLM_L_X76Y123_SLICE_X117Y123_A4 = CLBLM_L_X74Y123_SLICE_X113Y123_A5Q;
  assign CLBLM_L_X76Y123_SLICE_X117Y123_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X76Y123_SLICE_X117Y123_A6 = 1'b1;
  assign CLBLM_L_X76Y123_SLICE_X117Y123_B1 = CLBLM_L_X76Y123_SLICE_X117Y123_B5Q;
  assign CLBLM_L_X76Y123_SLICE_X117Y123_B2 = CLBLM_L_X76Y123_SLICE_X117Y123_BQ;
  assign CLBLM_L_X76Y123_SLICE_X117Y123_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X76Y123_SLICE_X117Y123_B4 = CLBLM_L_X76Y125_SLICE_X117Y125_BQ;
  assign CLBLM_L_X76Y123_SLICE_X117Y123_B5 = CLBLM_L_X76Y130_SLICE_X116Y130_DQ;
  assign CLBLM_L_X76Y123_SLICE_X117Y123_B6 = 1'b1;
  assign CLBLM_R_X67Y105_SLICE_X101Y105_D5 = CLBLM_R_X67Y103_SLICE_X100Y103_AO6;
  assign CLBLM_L_X76Y123_SLICE_X117Y123_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X76Y123_SLICE_X117Y123_C2 = CLBLM_L_X76Y123_SLICE_X117Y123_CQ;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_C2 = 1'b1;
  assign CLBLM_L_X76Y123_SLICE_X117Y123_C3 = CLBLM_L_X76Y125_SLICE_X117Y125_BQ;
  assign CLBLM_L_X76Y123_SLICE_X117Y123_C4 = CLBLM_L_X76Y122_SLICE_X117Y122_AQ;
  assign CLBLM_L_X76Y123_SLICE_X117Y123_C5 = CLBLM_L_X76Y123_SLICE_X117Y123_B5Q;
  assign CLBLM_L_X76Y123_SLICE_X117Y123_C6 = CLBLL_R_X77Y113_SLICE_X118Y113_AQ;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_C3 = 1'b1;
  assign CLBLM_L_X76Y123_SLICE_X117Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X67Y105_SLICE_X101Y105_D6 = CLBLM_R_X67Y105_SLICE_X101Y105_BO6;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_C4 = 1'b1;
  assign CLBLM_L_X76Y123_SLICE_X117Y123_D1 = CLBLM_L_X76Y122_SLICE_X116Y122_C5Q;
  assign CLBLM_L_X76Y123_SLICE_X117Y123_D2 = CLBLL_R_X77Y123_SLICE_X119Y123_BO6;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_C5 = 1'b1;
  assign CLBLM_L_X76Y123_SLICE_X117Y123_D3 = CLBLM_L_X76Y125_SLICE_X117Y125_BQ;
  assign CLBLM_L_X76Y123_SLICE_X117Y123_D4 = CLBLM_L_X76Y124_SLICE_X116Y124_CQ;
  assign CLBLM_L_X70Y103_SLICE_X105Y103_A1 = CLBLM_L_X70Y103_SLICE_X104Y103_C5Q;
  assign CLBLM_L_X70Y103_SLICE_X105Y103_A2 = CLBLM_L_X70Y103_SLICE_X105Y103_BQ;
  assign CLBLM_L_X70Y103_SLICE_X105Y103_A3 = CLBLM_L_X70Y103_SLICE_X104Y103_B5Q;
  assign CLBLM_L_X70Y103_SLICE_X105Y103_A4 = CLBLM_L_X70Y103_SLICE_X105Y103_AQ;
  assign CLBLM_L_X70Y103_SLICE_X105Y103_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y103_SLICE_X105Y103_A6 = CLBLM_L_X70Y104_SLICE_X104Y104_A5Q;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_C6 = 1'b1;
  assign CLBLM_L_X76Y123_SLICE_X117Y123_D5 = CLBLM_L_X76Y124_SLICE_X117Y124_AQ;
  assign CLBLM_L_X76Y123_SLICE_X116Y123_A1 = 1'b1;
  assign CLBLM_L_X70Y103_SLICE_X105Y103_B1 = CLBLM_L_X70Y103_SLICE_X104Y103_C5Q;
  assign CLBLM_L_X70Y103_SLICE_X105Y103_B2 = CLBLM_L_X70Y103_SLICE_X105Y103_BQ;
  assign CLBLM_L_X70Y103_SLICE_X105Y103_B3 = CLBLM_L_X70Y103_SLICE_X104Y103_B5Q;
  assign CLBLM_L_X70Y103_SLICE_X105Y103_B4 = CLBLL_R_X79Y99_SLICE_X122Y99_AO6;
  assign CLBLM_L_X70Y103_SLICE_X105Y103_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y103_SLICE_X105Y103_B6 = CLBLM_L_X70Y104_SLICE_X104Y104_A5Q;
  assign CLBLM_L_X76Y123_SLICE_X116Y123_A2 = CLBLM_L_X76Y122_SLICE_X116Y122_A5Q;
  assign CLBLM_L_X76Y123_SLICE_X116Y123_A3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X76Y123_SLICE_X116Y123_A4 = CLBLM_L_X76Y122_SLICE_X116Y122_AQ;
  assign CLBLM_L_X70Y103_SLICE_X105Y103_C1 = 1'b1;
  assign CLBLM_L_X70Y103_SLICE_X105Y103_C2 = CLBLM_L_X70Y104_SLICE_X104Y104_A5Q;
  assign CLBLM_L_X70Y103_SLICE_X105Y103_C3 = CLBLM_L_X70Y103_SLICE_X104Y103_B5Q;
  assign CLBLM_L_X70Y103_SLICE_X105Y103_C4 = 1'b1;
  assign CLBLM_L_X70Y103_SLICE_X105Y103_C5 = 1'b1;
  assign CLBLM_L_X70Y103_SLICE_X105Y103_C6 = 1'b1;
  assign CLBLM_L_X76Y123_SLICE_X116Y123_AX = CLBLL_R_X75Y123_SLICE_X115Y123_AO6;
  assign CLBLM_L_X76Y123_SLICE_X116Y123_B1 = CLBLM_L_X76Y123_SLICE_X116Y123_CQ;
  assign CLBLM_L_X70Y103_SLICE_X105Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X76Y123_SLICE_X116Y123_C1 = CLBLM_L_X74Y123_SLICE_X113Y123_CO5;
  assign CLBLM_L_X76Y123_SLICE_X116Y123_C2 = CLBLM_L_X76Y123_SLICE_X116Y123_CQ;
  assign CLBLM_L_X76Y123_SLICE_X116Y123_C3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X76Y123_SLICE_X116Y123_C4 = CLBLL_R_X75Y121_SLICE_X114Y121_BQ;
  assign CLBLM_L_X70Y103_SLICE_X105Y103_D1 = 1'b1;
  assign CLBLM_L_X70Y103_SLICE_X105Y103_D2 = CLBLM_L_X70Y103_SLICE_X104Y103_BQ;
  assign CLBLM_L_X70Y103_SLICE_X105Y103_D3 = 1'b1;
  assign CLBLM_L_X70Y103_SLICE_X105Y103_D4 = CLBLM_L_X70Y103_SLICE_X104Y103_CQ;
  assign CLBLM_L_X70Y103_SLICE_X105Y103_D5 = 1'b1;
  assign CLBLM_L_X70Y103_SLICE_X105Y103_D6 = 1'b1;
  assign CLBLM_L_X76Y123_SLICE_X116Y123_C5 = 1'b1;
  assign CLBLM_L_X76Y123_SLICE_X116Y123_C6 = CLBLL_R_X75Y123_SLICE_X115Y123_AQ;
  assign CLBLM_L_X70Y103_SLICE_X105Y103_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X76Y123_SLICE_X116Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X70Y103_SLICE_X104Y103_A1 = CLBLM_L_X70Y103_SLICE_X104Y103_AQ;
  assign CLBLM_L_X70Y103_SLICE_X104Y103_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y103_SLICE_X104Y103_A3 = CLBLM_R_X65Y103_SLICE_X99Y103_DO6;
  assign CLBLM_L_X70Y103_SLICE_X104Y103_A4 = 1'b1;
  assign CLBLM_L_X70Y103_SLICE_X104Y103_A5 = CLBLM_L_X70Y102_SLICE_X104Y102_AQ;
  assign CLBLM_L_X70Y103_SLICE_X104Y103_A6 = CLBLM_L_X70Y101_SLICE_X105Y101_CO6;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_D1 = 1'b1;
  assign CLBLM_L_X76Y123_SLICE_X116Y123_D1 = CLBLM_L_X76Y123_SLICE_X117Y123_AQ;
  assign CLBLM_L_X76Y123_SLICE_X116Y123_D2 = CLBLM_L_X74Y123_SLICE_X113Y123_A5Q;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_D2 = 1'b1;
  assign CLBLM_L_X70Y103_SLICE_X104Y103_B1 = CLBLM_L_X70Y103_SLICE_X104Y103_B5Q;
  assign CLBLM_L_X70Y103_SLICE_X104Y103_B2 = CLBLM_L_X70Y103_SLICE_X104Y103_BQ;
  assign CLBLM_L_X70Y103_SLICE_X104Y103_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y103_SLICE_X104Y103_B4 = 1'b1;
  assign CLBLM_L_X70Y103_SLICE_X104Y103_B5 = CLBLM_L_X70Y103_SLICE_X104Y103_C5Q;
  assign CLBLM_L_X70Y103_SLICE_X104Y103_B6 = 1'b1;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_D3 = 1'b1;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_D4 = 1'b1;
  assign CLBLM_L_X70Y103_SLICE_X104Y103_C1 = CLBLM_L_X70Y103_SLICE_X104Y103_C5Q;
  assign CLBLM_L_X70Y103_SLICE_X104Y103_C2 = CLBLM_L_X70Y103_SLICE_X104Y103_CQ;
  assign CLBLM_L_X70Y103_SLICE_X104Y103_C3 = 1'b1;
  assign CLBLM_L_X70Y103_SLICE_X104Y103_C4 = CLBLM_L_X70Y103_SLICE_X104Y103_BQ;
  assign CLBLM_L_X70Y103_SLICE_X104Y103_C5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y103_SLICE_X104Y103_C6 = 1'b1;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_D5 = 1'b1;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_D6 = 1'b1;
  assign CLBLM_L_X70Y103_SLICE_X104Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X70Y103_SLICE_X104Y103_D1 = CLBLM_L_X70Y103_SLICE_X104Y103_C5Q;
  assign CLBLM_L_X70Y103_SLICE_X104Y103_D2 = CLBLM_L_X70Y103_SLICE_X104Y103_CQ;
  assign CLBLM_L_X70Y103_SLICE_X104Y103_D3 = CLBLM_L_X70Y103_SLICE_X104Y103_BQ;
  assign CLBLM_L_X70Y103_SLICE_X104Y103_D4 = 1'b1;
  assign CLBLM_L_X70Y103_SLICE_X104Y103_D5 = 1'b1;
  assign CLBLM_L_X70Y103_SLICE_X104Y103_D6 = 1'b1;
  assign CLBLM_L_X70Y103_SLICE_X104Y103_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_A1 = CLBLM_L_X72Y120_SLICE_X108Y120_A5Q;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_A2 = CLBLM_L_X72Y120_SLICE_X108Y120_BQ;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_A3 = CLBLM_L_X72Y120_SLICE_X108Y120_AQ;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_A5 = CLBLM_L_X72Y118_SLICE_X109Y118_AQ;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_A6 = 1'b1;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_B1 = 1'b1;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_B2 = CLBLM_L_X72Y120_SLICE_X108Y120_BQ;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_B3 = 1'b1;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_B5 = 1'b1;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_B6 = 1'b1;
  assign LIOB33_X0Y153_IOB_X0Y154_O = CLBLM_R_X67Y118_SLICE_X100Y118_A5Q;
  assign LIOB33_X0Y153_IOB_X0Y153_O = CLBLM_R_X65Y106_SLICE_X99Y106_DQ;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_C5 = 1'b1;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_C6 = 1'b1;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_A1 = CLBLM_L_X76Y122_SLICE_X116Y122_C5Q;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_A2 = CLBLM_L_X76Y124_SLICE_X116Y124_BO6;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_A3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_A4 = CLBLM_L_X76Y124_SLICE_X117Y124_AQ;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_A5 = CLBLM_L_X74Y123_SLICE_X113Y123_CO5;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_A6 = 1'b1;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_B1 = CLBLL_R_X77Y123_SLICE_X119Y123_CQ;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_B2 = CLBLM_L_X76Y124_SLICE_X117Y124_BQ;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_B3 = CLBLL_R_X75Y113_SLICE_X114Y113_AQ;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_B5 = CLBLM_L_X76Y123_SLICE_X117Y123_AQ;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_B6 = CLBLM_L_X74Y123_SLICE_X113Y123_A5Q;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_C2 = CLBLM_L_X76Y119_SLICE_X116Y119_BO6;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_C3 = CLBLL_R_X75Y122_SLICE_X114Y122_AQ;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_C4 = CLBLM_L_X76Y123_SLICE_X117Y123_AO5;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_C5 = CLBLM_L_X76Y125_SLICE_X117Y125_BQ;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_C6 = 1'b1;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_D1 = 1'b1;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_D1 = 1'b1;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_D2 = CLBLM_L_X76Y124_SLICE_X117Y124_AQ;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_D3 = CLBLM_L_X76Y124_SLICE_X116Y124_B5Q;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_D4 = CLBLM_L_X76Y125_SLICE_X117Y125_BQ;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_D2 = 1'b1;
  assign CLBLM_L_X70Y104_SLICE_X105Y104_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y104_SLICE_X105Y104_A2 = 1'b1;
  assign CLBLM_L_X70Y104_SLICE_X105Y104_A3 = CLBLM_L_X70Y104_SLICE_X105Y104_AQ;
  assign CLBLM_L_X70Y104_SLICE_X105Y104_A4 = CLBLM_L_X70Y101_SLICE_X105Y101_CO6;
  assign CLBLM_L_X70Y104_SLICE_X105Y104_A5 = CLBLM_L_X70Y103_SLICE_X105Y103_AQ;
  assign CLBLM_L_X70Y104_SLICE_X105Y104_A6 = CLBLM_L_X70Y101_SLICE_X104Y101_AO5;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_D3 = 1'b1;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_D5 = CLBLM_L_X76Y122_SLICE_X116Y122_C5Q;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_D4 = 1'b1;
  assign CLBLM_L_X70Y104_SLICE_X105Y104_B1 = CLBLM_L_X70Y102_SLICE_X105Y102_DO6;
  assign CLBLM_L_X70Y104_SLICE_X105Y104_B2 = CLBLM_L_X70Y104_SLICE_X105Y104_BQ;
  assign CLBLM_L_X70Y104_SLICE_X105Y104_B3 = CLBLM_L_X70Y104_SLICE_X105Y104_AQ;
  assign CLBLM_L_X70Y104_SLICE_X105Y104_B4 = 1'b1;
  assign CLBLM_L_X70Y104_SLICE_X105Y104_B5 = CLBLM_L_X70Y103_SLICE_X105Y103_AQ;
  assign CLBLM_L_X70Y104_SLICE_X105Y104_B6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_D5 = 1'b1;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_A1 = 1'b1;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_D6 = 1'b1;
  assign CLBLM_L_X70Y104_SLICE_X105Y104_C1 = CLBLM_L_X70Y104_SLICE_X105Y104_BQ;
  assign CLBLM_L_X70Y104_SLICE_X105Y104_C2 = CLBLM_L_X70Y104_SLICE_X105Y104_CQ;
  assign CLBLM_L_X70Y104_SLICE_X105Y104_C3 = CLBLM_L_X70Y103_SLICE_X104Y103_B5Q;
  assign CLBLM_L_X70Y104_SLICE_X105Y104_C4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y104_SLICE_X105Y104_C5 = CLBLM_L_X70Y104_SLICE_X104Y104_A5Q;
  assign CLBLM_L_X70Y104_SLICE_X105Y104_C6 = CLBLM_L_X70Y103_SLICE_X104Y103_C5Q;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_AX = CLBLM_L_X76Y124_SLICE_X116Y124_B5Q;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_B1 = CLBLM_L_X76Y124_SLICE_X116Y124_A5Q;
  assign CLBLM_L_X70Y104_SLICE_X105Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_B2 = CLBLM_L_X76Y124_SLICE_X116Y124_BQ;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_B3 = CLBLM_L_X76Y124_SLICE_X116Y124_AQ;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_B4 = CLBLL_R_X75Y124_SLICE_X115Y124_AQ;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_B5 = CLBLM_L_X76Y124_SLICE_X116Y124_CQ;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_BX = CLBLL_R_X75Y124_SLICE_X115Y124_DQ;
  assign CLBLM_L_X70Y104_SLICE_X105Y104_D1 = CLBLM_L_X70Y104_SLICE_X105Y104_DQ;
  assign CLBLM_L_X70Y104_SLICE_X105Y104_D2 = CLBLM_L_X70Y104_SLICE_X105Y104_CQ;
  assign CLBLM_L_X70Y104_SLICE_X105Y104_D3 = CLBLM_L_X70Y104_SLICE_X105Y104_D5Q;
  assign CLBLM_L_X70Y104_SLICE_X105Y104_D4 = CLBLM_L_X70Y102_SLICE_X105Y102_DO6;
  assign CLBLM_L_X70Y104_SLICE_X105Y104_D5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y104_SLICE_X105Y104_D6 = 1'b1;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_C4 = CLBLL_R_X75Y123_SLICE_X115Y123_AO5;
  assign CLBLM_L_X70Y104_SLICE_X105Y104_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_CX = CLBLM_L_X76Y124_SLICE_X117Y124_AQ;
  assign CLBLM_L_X70Y104_SLICE_X104Y104_A1 = CLBLM_L_X70Y105_SLICE_X105Y105_A5Q;
  assign CLBLM_L_X70Y104_SLICE_X104Y104_A2 = CLBLM_L_X70Y103_SLICE_X104Y103_C5Q;
  assign CLBLM_L_X70Y104_SLICE_X104Y104_A3 = CLBLM_L_X70Y104_SLICE_X104Y104_AQ;
  assign CLBLM_L_X70Y104_SLICE_X104Y104_A4 = CLBLM_L_X70Y103_SLICE_X104Y103_B5Q;
  assign CLBLM_L_X70Y104_SLICE_X104Y104_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y104_SLICE_X104Y104_A6 = CLBLM_L_X70Y104_SLICE_X104Y104_A5Q;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_D1 = 1'b1;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_D2 = 1'b1;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_D3 = 1'b1;
  assign CLBLM_L_X70Y104_SLICE_X104Y104_AX = CLBLM_L_X70Y104_SLICE_X104Y104_CO6;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_D4 = 1'b1;
  assign CLBLM_L_X70Y104_SLICE_X104Y104_B1 = CLBLM_L_X70Y105_SLICE_X105Y105_A5Q;
  assign CLBLM_L_X70Y104_SLICE_X104Y104_B2 = CLBLM_L_X70Y104_SLICE_X104Y104_BQ;
  assign CLBLM_L_X70Y104_SLICE_X104Y104_B3 = CLBLM_L_X70Y104_SLICE_X104Y104_AQ;
  assign CLBLM_L_X70Y104_SLICE_X104Y104_B4 = 1'b1;
  assign CLBLM_L_X70Y104_SLICE_X104Y104_B5 = CLBLM_L_X70Y104_SLICE_X104Y104_CO5;
  assign CLBLM_L_X70Y104_SLICE_X104Y104_B6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_B5 = 1'b1;
  assign CLBLM_L_X70Y104_SLICE_X104Y104_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y104_SLICE_X104Y104_C2 = 1'b1;
  assign CLBLM_L_X70Y104_SLICE_X104Y104_C3 = CLBLM_L_X70Y104_SLICE_X104Y104_A5Q;
  assign CLBLM_L_X70Y104_SLICE_X104Y104_C4 = CLBLM_L_X70Y103_SLICE_X104Y103_B5Q;
  assign CLBLM_L_X70Y104_SLICE_X104Y104_C5 = CLBLM_L_X70Y103_SLICE_X104Y103_C5Q;
  assign CLBLM_L_X70Y104_SLICE_X104Y104_C6 = 1'b1;
  assign CLBLM_L_X70Y104_SLICE_X104Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X70Y104_SLICE_X104Y104_D1 = 1'b1;
  assign CLBLM_L_X70Y104_SLICE_X104Y104_D2 = 1'b1;
  assign CLBLM_L_X70Y104_SLICE_X104Y104_D3 = 1'b1;
  assign CLBLM_L_X70Y104_SLICE_X104Y104_D4 = 1'b1;
  assign CLBLM_L_X70Y104_SLICE_X104Y104_D5 = 1'b1;
  assign CLBLM_L_X70Y104_SLICE_X104Y104_D6 = 1'b1;
  assign CLBLM_L_X70Y104_SLICE_X104Y104_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X67Y109_SLICE_X101Y109_D2 = CLBLM_L_X68Y108_SLICE_X102Y108_A5Q;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_D5 = 1'b1;
  assign LIOI3_X0Y97_OLOGIC_X0Y98_D1 = CLBLM_L_X68Y97_SLICE_X103Y97_AQ;
  assign LIOI3_X0Y97_OLOGIC_X0Y98_T1 = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_D1 = CLBLL_R_X73Y103_SLICE_X110Y103_A5Q;
  assign LIOB33_X0Y155_IOB_X0Y156_O = CLBLM_L_X64Y99_SLICE_X97Y99_B5Q;
  assign LIOB33_X0Y155_IOB_X0Y155_O = CLBLM_L_X76Y118_SLICE_X117Y118_CQ;
  assign LIOI3_X0Y97_OLOGIC_X0Y97_D1 = CLBLM_L_X62Y103_SLICE_X92Y103_A5Q;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_T1 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_A1 = 1'b1;
  assign LIOI3_X0Y97_OLOGIC_X0Y97_T1 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_A3 = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_D1 = CLBLM_R_X65Y110_SLICE_X99Y110_AQ;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_A5 = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_T1 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_A6 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_B1 = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_D1 = CLBLM_L_X64Y99_SLICE_X97Y99_B5Q;
  assign CLBLM_R_X67Y109_SLICE_X101Y109_D3 = CLBLM_R_X67Y109_SLICE_X100Y109_DO6;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_B3 = 1'b1;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_A1 = CLBLL_R_X77Y123_SLICE_X119Y123_DO6;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_A2 = CLBLM_L_X76Y126_SLICE_X117Y126_AQ;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_A3 = CLBLM_L_X76Y125_SLICE_X117Y125_AQ;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_A4 = CLBLL_R_X75Y123_SLICE_X115Y123_DO6;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_A6 = CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  assign CLBLM_L_X82Y130_SLICE_X129Y130_B3 = 1'b1;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_B1 = CLBLM_L_X76Y125_SLICE_X117Y125_DO6;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_B2 = CLBLM_L_X76Y125_SLICE_X117Y125_BQ;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_B3 = CLBLM_L_X76Y123_SLICE_X117Y123_AQ;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_B4 = CLBLL_R_X75Y113_SLICE_X114Y113_AQ;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_B5 = CLBLM_L_X76Y124_SLICE_X117Y124_CO6;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_B6 = CLBLM_L_X74Y123_SLICE_X113Y123_A5Q;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_A1 = 1'b1;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_A2 = 1'b1;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_A3 = 1'b1;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_A4 = 1'b1;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_A5 = 1'b1;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_A6 = 1'b1;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_C1 = CLBLL_R_X77Y125_SLICE_X118Y125_BQ;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_C2 = CLBLM_L_X76Y124_SLICE_X116Y124_CO6;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_B1 = 1'b1;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_B2 = 1'b1;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_B3 = 1'b1;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_B4 = 1'b1;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_B5 = 1'b1;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_B6 = 1'b1;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_C4 = CLBLM_L_X74Y123_SLICE_X113Y123_A5Q;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_C5 = CLBLM_L_X76Y123_SLICE_X117Y123_AQ;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_C1 = 1'b1;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_C2 = 1'b1;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_C3 = 1'b1;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_C4 = 1'b1;
  assign CLBLM_L_X70Y105_SLICE_X105Y105_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y105_SLICE_X105Y105_A2 = CLBLM_L_X70Y104_SLICE_X105Y104_D5Q;
  assign CLBLM_L_X70Y105_SLICE_X105Y105_A3 = CLBLM_L_X70Y105_SLICE_X105Y105_A5Q;
  assign CLBLM_L_X70Y105_SLICE_X105Y105_A4 = CLBLM_L_X70Y101_SLICE_X104Y101_AO5;
  assign CLBLM_L_X70Y105_SLICE_X105Y105_A5 = CLBLL_R_X75Y122_SLICE_X115Y122_AQ;
  assign CLBLM_L_X70Y105_SLICE_X105Y105_A6 = 1'b1;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_C5 = 1'b1;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_C6 = 1'b1;
  assign CLBLM_L_X70Y105_SLICE_X105Y105_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y105_SLICE_X105Y105_B2 = CLBLM_L_X70Y105_SLICE_X104Y105_BO6;
  assign CLBLM_L_X70Y105_SLICE_X105Y105_B3 = CLBLM_L_X72Y104_SLICE_X109Y104_DO6;
  assign CLBLM_L_X70Y105_SLICE_X105Y105_B4 = CLBLM_L_X68Y108_SLICE_X103Y108_CO6;
  assign CLBLM_L_X70Y105_SLICE_X105Y105_B5 = CLBLM_L_X68Y109_SLICE_X103Y109_B5Q;
  assign CLBLM_L_X70Y105_SLICE_X105Y105_B6 = CLBLM_L_X68Y109_SLICE_X103Y109_BQ;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_D1 = 1'b1;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_D2 = 1'b1;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_D3 = 1'b1;
  assign CLBLM_L_X70Y105_SLICE_X105Y105_C1 = 1'b1;
  assign CLBLM_L_X70Y105_SLICE_X105Y105_C2 = 1'b1;
  assign CLBLM_L_X70Y105_SLICE_X105Y105_C3 = 1'b1;
  assign CLBLM_L_X70Y105_SLICE_X105Y105_C4 = 1'b1;
  assign CLBLM_L_X70Y105_SLICE_X105Y105_C5 = 1'b1;
  assign CLBLM_L_X70Y105_SLICE_X105Y105_C6 = 1'b1;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_A1 = 1'b1;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_A2 = 1'b1;
  assign CLBLM_L_X70Y105_SLICE_X105Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_A3 = 1'b1;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_A4 = 1'b1;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_A5 = 1'b1;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_A6 = 1'b1;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_AX = CLBLM_L_X72Y116_SLICE_X108Y116_AQ;
  assign CLBLM_L_X70Y105_SLICE_X105Y105_D1 = 1'b1;
  assign CLBLM_L_X70Y105_SLICE_X105Y105_D2 = 1'b1;
  assign CLBLM_L_X70Y105_SLICE_X105Y105_D3 = 1'b1;
  assign CLBLM_L_X70Y105_SLICE_X105Y105_D4 = 1'b1;
  assign CLBLM_L_X70Y105_SLICE_X105Y105_D5 = 1'b1;
  assign CLBLM_L_X70Y105_SLICE_X105Y105_D6 = 1'b1;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_B1 = 1'b1;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_B2 = 1'b1;
  assign CLBLM_L_X70Y105_SLICE_X105Y105_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_B3 = 1'b1;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_B4 = 1'b1;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_B5 = 1'b1;
  assign CLBLM_L_X70Y105_SLICE_X104Y105_A1 = CLBLM_L_X68Y109_SLICE_X103Y109_B5Q;
  assign CLBLM_L_X70Y105_SLICE_X104Y105_A2 = CLBLM_L_X68Y109_SLICE_X103Y109_BQ;
  assign CLBLM_L_X70Y105_SLICE_X104Y105_A3 = CLBLM_L_X70Y105_SLICE_X104Y105_AQ;
  assign CLBLM_L_X70Y105_SLICE_X104Y105_A4 = CLBLM_L_X70Y105_SLICE_X105Y105_BQ;
  assign CLBLM_L_X70Y105_SLICE_X104Y105_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y105_SLICE_X104Y105_A6 = CLBLM_L_X68Y108_SLICE_X103Y108_CO6;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_C1 = 1'b1;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_C2 = 1'b1;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_C3 = 1'b1;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_C4 = 1'b1;
  assign CLBLM_L_X70Y105_SLICE_X104Y105_B1 = CLBLM_L_X68Y106_SLICE_X103Y106_DO6;
  assign CLBLM_L_X70Y105_SLICE_X104Y105_B2 = CLBLM_L_X68Y109_SLICE_X103Y109_B5Q;
  assign CLBLM_L_X70Y105_SLICE_X104Y105_B3 = CLBLM_L_X70Y105_SLICE_X104Y105_AQ;
  assign CLBLM_L_X70Y105_SLICE_X104Y105_B4 = CLBLM_L_X70Y106_SLICE_X104Y106_BQ;
  assign CLBLM_L_X70Y105_SLICE_X104Y105_B5 = 1'b1;
  assign CLBLM_L_X70Y105_SLICE_X104Y105_B6 = CLBLM_L_X68Y109_SLICE_X103Y109_BQ;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_D1 = 1'b1;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_D2 = 1'b1;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_D3 = 1'b1;
  assign CLBLM_L_X70Y105_SLICE_X104Y105_C1 = CLBLM_L_X68Y103_SLICE_X102Y103_AQ;
  assign CLBLM_L_X70Y105_SLICE_X104Y105_C2 = 1'b1;
  assign CLBLM_L_X70Y105_SLICE_X104Y105_C3 = CLBLM_L_X72Y104_SLICE_X108Y104_DQ;
  assign CLBLM_L_X70Y105_SLICE_X104Y105_C4 = CLBLM_L_X70Y106_SLICE_X104Y106_AQ;
  assign CLBLM_L_X70Y105_SLICE_X104Y105_C5 = 1'b1;
  assign CLBLM_L_X70Y105_SLICE_X104Y105_C6 = CLBLM_L_X70Y106_SLICE_X104Y106_BQ;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_D6 = 1'b1;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X70Y105_SLICE_X104Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X70Y105_SLICE_X104Y105_D1 = 1'b1;
  assign CLBLM_L_X70Y105_SLICE_X104Y105_D2 = 1'b1;
  assign CLBLM_L_X70Y105_SLICE_X104Y105_D3 = 1'b1;
  assign CLBLM_L_X70Y105_SLICE_X104Y105_D4 = 1'b1;
  assign CLBLM_L_X70Y105_SLICE_X104Y105_D5 = 1'b1;
  assign CLBLM_L_X70Y105_SLICE_X104Y105_D6 = 1'b1;
  assign CLBLM_L_X70Y105_SLICE_X104Y105_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X76Y129_SLICE_X116Y129_C3 = CLBLM_L_X76Y129_SLICE_X116Y129_AQ;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_T1 = 1'b1;
  assign RIOB33_X105Y167_IOB_X1Y167_O = 1'b1;
  assign LIOB33_X0Y157_IOB_X0Y158_O = CLBLM_L_X76Y125_SLICE_X116Y125_AQ;
  assign LIOB33_X0Y157_IOB_X0Y157_O = CLBLM_R_X63Y122_SLICE_X95Y122_CQ;
  assign CLBLM_L_X76Y129_SLICE_X116Y129_C5 = CLBLM_L_X76Y129_SLICE_X116Y129_B5Q;
  assign CLBLM_R_X67Y109_SLICE_X101Y109_D5 = CLBLM_L_X76Y111_SLICE_X116Y111_AQ;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_D1 = 1'b1;
  assign CLBLM_L_X76Y122_SLICE_X117Y122_D5 = 1'b1;
  assign CLBLM_L_X76Y122_SLICE_X117Y122_D6 = 1'b1;
  assign CLBLM_L_X76Y126_SLICE_X117Y126_A1 = CLBLM_L_X76Y126_SLICE_X116Y126_DQ;
  assign CLBLM_L_X76Y126_SLICE_X117Y126_A2 = CLBLL_R_X77Y127_SLICE_X119Y127_AO5;
  assign CLBLM_L_X76Y122_SLICE_X117Y122_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X76Y126_SLICE_X117Y126_A3 = CLBLM_L_X76Y126_SLICE_X117Y126_AQ;
  assign CLBLM_L_X76Y126_SLICE_X117Y126_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X76Y126_SLICE_X117Y126_A5 = 1'b1;
  assign CLBLM_L_X76Y126_SLICE_X117Y126_A6 = CLBLM_L_X76Y126_SLICE_X116Y126_AO6;
  assign CLBLM_L_X76Y126_SLICE_X117Y126_B1 = 1'b1;
  assign CLBLM_L_X76Y126_SLICE_X117Y126_B2 = 1'b1;
  assign CLBLM_L_X76Y126_SLICE_X117Y126_B3 = 1'b1;
  assign CLBLM_L_X76Y126_SLICE_X117Y126_B4 = 1'b1;
  assign CLBLM_L_X76Y126_SLICE_X117Y126_B5 = 1'b1;
  assign CLBLM_L_X76Y126_SLICE_X117Y126_B6 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_A1 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_A2 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_A3 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_A4 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_A5 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_A6 = 1'b1;
  assign CLBLM_L_X76Y126_SLICE_X117Y126_C1 = 1'b1;
  assign CLBLM_L_X76Y126_SLICE_X117Y126_C2 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_B1 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_B2 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_B3 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_B4 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_B5 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_B6 = 1'b1;
  assign CLBLM_L_X76Y126_SLICE_X117Y126_C4 = 1'b1;
  assign CLBLM_L_X76Y126_SLICE_X117Y126_C5 = 1'b1;
  assign CLBLM_L_X76Y126_SLICE_X117Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_C1 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_C2 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_C3 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_C4 = 1'b1;
  assign CLBLM_L_X70Y106_SLICE_X105Y106_A1 = CLBLM_L_X70Y106_SLICE_X105Y106_AQ;
  assign CLBLM_L_X70Y106_SLICE_X105Y106_A2 = CLBLM_L_X68Y108_SLICE_X103Y108_CO6;
  assign CLBLM_L_X70Y106_SLICE_X105Y106_A3 = CLBLM_L_X68Y109_SLICE_X103Y109_B5Q;
  assign CLBLM_L_X70Y106_SLICE_X105Y106_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y106_SLICE_X105Y106_A5 = CLBLM_L_X68Y109_SLICE_X103Y109_BQ;
  assign CLBLM_L_X70Y106_SLICE_X105Y106_A6 = CLBLM_L_X70Y107_SLICE_X105Y107_BQ;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_C5 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_C6 = 1'b1;
  assign CLBLM_L_X70Y106_SLICE_X105Y106_AX = CLBLM_L_X70Y106_SLICE_X104Y106_A5Q;
  assign CLBLM_L_X70Y106_SLICE_X105Y106_B1 = CLBLM_L_X68Y108_SLICE_X103Y108_CO6;
  assign CLBLM_L_X70Y106_SLICE_X105Y106_B2 = CLBLM_L_X70Y106_SLICE_X105Y106_BQ;
  assign CLBLM_L_X70Y106_SLICE_X105Y106_B3 = CLBLM_L_X68Y109_SLICE_X103Y109_B5Q;
  assign CLBLM_L_X70Y106_SLICE_X105Y106_B4 = CLBLM_L_X68Y108_SLICE_X103Y108_BQ;
  assign CLBLM_L_X70Y106_SLICE_X105Y106_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y106_SLICE_X105Y106_B6 = CLBLM_L_X68Y109_SLICE_X103Y109_BQ;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_D1 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_D2 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_D3 = 1'b1;
  assign CLBLM_L_X70Y106_SLICE_X105Y106_C1 = CLBLM_L_X70Y106_SLICE_X104Y106_A5Q;
  assign CLBLM_L_X70Y106_SLICE_X105Y106_C2 = CLBLM_L_X68Y109_SLICE_X103Y109_B5Q;
  assign CLBLM_L_X70Y106_SLICE_X105Y106_C3 = CLBLM_L_X68Y106_SLICE_X103Y106_DO6;
  assign CLBLM_L_X70Y106_SLICE_X105Y106_C4 = CLBLM_L_X68Y109_SLICE_X103Y109_BQ;
  assign CLBLM_L_X70Y106_SLICE_X105Y106_C5 = CLBLM_L_X70Y106_SLICE_X105Y106_AQ;
  assign CLBLM_L_X70Y106_SLICE_X105Y106_C6 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_A1 = CLBLM_L_X74Y119_SLICE_X112Y119_DQ;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_A2 = CLBLL_R_X75Y124_SLICE_X115Y124_BQ;
  assign CLBLM_L_X70Y106_SLICE_X105Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_A3 = CLBLM_L_X74Y118_SLICE_X112Y118_AQ;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_A4 = CLBLM_L_X74Y118_SLICE_X112Y118_BO6;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_A6 = CLBLM_L_X74Y119_SLICE_X113Y119_AO6;
  assign CLBLM_L_X70Y106_SLICE_X105Y106_D1 = 1'b1;
  assign CLBLM_L_X70Y106_SLICE_X105Y106_D2 = CLBLM_L_X68Y109_SLICE_X103Y109_BQ;
  assign CLBLM_L_X70Y106_SLICE_X105Y106_D3 = CLBLM_L_X70Y106_SLICE_X105Y106_BQ;
  assign CLBLM_L_X70Y106_SLICE_X105Y106_D4 = CLBLM_L_X68Y109_SLICE_X103Y109_B5Q;
  assign CLBLM_L_X70Y106_SLICE_X105Y106_D5 = CLBLM_L_X68Y106_SLICE_X103Y106_DO6;
  assign CLBLM_L_X70Y106_SLICE_X105Y106_D6 = CLBLM_L_X70Y106_SLICE_X105Y106_A5Q;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_B1 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_B2 = 1'b1;
  assign CLBLM_L_X70Y106_SLICE_X105Y106_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_B3 = CLBLM_L_X72Y118_SLICE_X108Y118_CQ;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_B4 = CLBLM_R_X65Y105_SLICE_X99Y105_CQ;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_B5 = 1'b1;
  assign CLBLM_L_X70Y106_SLICE_X104Y106_A1 = CLBLM_L_X70Y106_SLICE_X105Y106_A5Q;
  assign CLBLM_L_X70Y106_SLICE_X104Y106_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y106_SLICE_X104Y106_A3 = CLBLM_L_X70Y106_SLICE_X104Y106_AQ;
  assign CLBLM_L_X70Y106_SLICE_X104Y106_A4 = CLBLM_L_X68Y105_SLICE_X102Y105_CQ;
  assign CLBLM_L_X70Y106_SLICE_X104Y106_A5 = CLBLM_L_X68Y106_SLICE_X103Y106_AO6;
  assign CLBLM_L_X70Y106_SLICE_X104Y106_A6 = CLBLM_L_X70Y106_SLICE_X104Y106_A5Q;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_C2 = CLBLM_L_X74Y118_SLICE_X112Y118_CQ;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_C3 = CLBLM_L_X74Y118_SLICE_X112Y118_AQ;
  assign CLBLM_L_X70Y106_SLICE_X104Y106_AX = CLBLM_L_X70Y106_SLICE_X104Y106_AQ;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_C4 = CLBLM_L_X74Y119_SLICE_X113Y119_AO6;
  assign CLBLM_L_X70Y106_SLICE_X104Y106_B1 = CLBLM_L_X70Y106_SLICE_X105Y106_AQ;
  assign CLBLM_L_X70Y106_SLICE_X104Y106_B2 = CLBLM_L_X68Y105_SLICE_X103Y105_AQ;
  assign CLBLM_L_X70Y106_SLICE_X104Y106_B3 = CLBLM_L_X70Y105_SLICE_X104Y105_AQ;
  assign CLBLM_L_X70Y106_SLICE_X104Y106_B4 = CLBLM_L_X70Y106_SLICE_X105Y106_BQ;
  assign CLBLM_L_X70Y106_SLICE_X104Y106_B5 = CLBLM_L_X68Y109_SLICE_X103Y109_B5Q;
  assign CLBLM_L_X70Y106_SLICE_X104Y106_B6 = CLBLM_L_X68Y109_SLICE_X103Y109_BQ;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_D1 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_D2 = 1'b1;
  assign CLBLM_L_X70Y106_SLICE_X104Y106_BX = CLBLM_L_X70Y106_SLICE_X105Y106_A5Q;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_D3 = 1'b1;
  assign CLBLM_L_X70Y106_SLICE_X104Y106_C1 = CLBLM_L_X68Y105_SLICE_X103Y105_AQ;
  assign CLBLM_L_X70Y106_SLICE_X104Y106_C2 = CLBLM_L_X68Y109_SLICE_X103Y109_B5Q;
  assign CLBLM_L_X70Y106_SLICE_X104Y106_C3 = CLBLM_L_X68Y106_SLICE_X103Y106_DO6;
  assign CLBLM_L_X70Y106_SLICE_X104Y106_C4 = CLBLM_L_X68Y109_SLICE_X103Y109_BQ;
  assign CLBLM_L_X70Y106_SLICE_X104Y106_C5 = 1'b1;
  assign CLBLM_L_X70Y106_SLICE_X104Y106_C6 = CLBLM_L_X70Y106_SLICE_X104Y106_AQ;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_D6 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X70Y106_SLICE_X104Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X70Y106_SLICE_X104Y106_D1 = 1'b1;
  assign CLBLM_L_X70Y106_SLICE_X104Y106_D2 = 1'b1;
  assign CLBLM_L_X70Y106_SLICE_X104Y106_D3 = 1'b1;
  assign CLBLM_L_X70Y106_SLICE_X104Y106_D4 = CLBLM_L_X70Y106_SLICE_X104Y106_A5Q;
  assign CLBLM_L_X70Y106_SLICE_X104Y106_D5 = CLBLM_L_X70Y106_SLICE_X105Y106_A5Q;
  assign CLBLM_L_X70Y106_SLICE_X104Y106_D6 = CLBLM_L_X70Y106_SLICE_X104Y106_AQ;
  assign CLBLM_L_X76Y122_SLICE_X116Y122_C1 = CLBLM_L_X76Y122_SLICE_X116Y122_C5Q;
  assign CLBLM_L_X70Y106_SLICE_X104Y106_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X76Y122_SLICE_X116Y122_C2 = CLBLM_L_X74Y123_SLICE_X113Y123_CO5;
  assign CLBLM_L_X76Y122_SLICE_X116Y122_C5 = CLBLL_R_X77Y127_SLICE_X118Y127_AQ;
  assign CLBLM_L_X76Y122_SLICE_X116Y122_C6 = 1'b1;
  assign LIOB33_X0Y159_IOB_X0Y160_O = CLBLL_R_X71Y119_SLICE_X106Y119_AQ;
  assign LIOB33_X0Y159_IOB_X0Y159_O = CLBLM_R_X67Y116_SLICE_X100Y116_AQ;
  assign LIOB33_X0Y81_IOB_X0Y82_O = CLBLM_L_X62Y107_SLICE_X93Y107_A5Q;
  assign LIOB33_X0Y81_IOB_X0Y81_O = CLBLM_L_X60Y99_SLICE_X90Y99_BQ;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign RIOB33_X105Y63_IOB_X1Y64_O = CLBLM_R_X103Y67_SLICE_X163Y67_AQ;
  assign CLBLM_L_X82Y130_SLICE_X129Y130_B4 = 1'b1;
  assign CLBLM_L_X76Y129_SLICE_X116Y129_D3 = CLBLL_R_X77Y129_SLICE_X118Y129_CQ;
  assign CLBLM_L_X76Y122_SLICE_X116Y122_D6 = 1'b1;
  assign CLBLM_L_X76Y122_SLICE_X116Y122_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X65Y111_SLICE_X98Y111_A1 = CLBLM_L_X60Y97_SLICE_X91Y97_AQ;
  assign CLBLM_R_X65Y111_SLICE_X98Y111_A2 = CLBLM_L_X76Y111_SLICE_X116Y111_AQ;
  assign CLBLM_R_X65Y111_SLICE_X98Y111_A3 = CLBLM_R_X65Y111_SLICE_X98Y111_AQ;
  assign CLBLM_R_X65Y111_SLICE_X98Y111_A4 = CLBLM_R_X65Y111_SLICE_X98Y111_BO6;
  assign CLBLM_R_X65Y111_SLICE_X98Y111_A5 = CLBLM_L_X62Y92_SLICE_X92Y92_BQ;
  assign RIOB33_X105Y111_IOB_X1Y112_O = CLBLL_R_X71Y100_SLICE_X106Y100_BQ;
  assign RIOB33_X105Y111_IOB_X1Y111_O = CLBLM_L_X62Y107_SLICE_X93Y107_BQ;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_A1 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_A2 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_A3 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_A4 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_A5 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_A6 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_D1 = RIOB33_X105Y59_IOB_X1Y59_I;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_B1 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_B2 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_B3 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_B4 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_B5 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_B6 = 1'b1;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_A1 = CLBLM_L_X70Y105_SLICE_X105Y105_AQ;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_A2 = CLBLM_L_X76Y122_SLICE_X116Y122_CQ;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_A3 = CLBLL_R_X75Y121_SLICE_X114Y121_AQ;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_A4 = CLBLM_L_X74Y121_SLICE_X113Y121_AQ;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_A5 = CLBLL_R_X75Y122_SLICE_X115Y122_AQ;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_A6 = CLBLM_L_X76Y125_SLICE_X116Y125_C5Q;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_C1 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_C2 = 1'b1;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_B1 = 1'b1;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_B2 = 1'b1;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_B3 = 1'b1;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_B4 = 1'b1;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_B5 = 1'b1;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_B6 = 1'b1;
  assign CLBLM_L_X76Y119_SLICE_X116Y119_B6 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_C5 = 1'b1;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_C1 = 1'b1;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_C2 = 1'b1;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_C3 = 1'b1;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_C4 = 1'b1;
  assign CLBLM_L_X70Y107_SLICE_X105Y107_A1 = CLBLM_L_X72Y106_SLICE_X108Y106_CO6;
  assign CLBLM_L_X70Y107_SLICE_X105Y107_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y107_SLICE_X105Y107_A3 = CLBLM_L_X70Y107_SLICE_X105Y107_AQ;
  assign CLBLM_L_X70Y107_SLICE_X105Y107_A4 = CLBLM_L_X70Y106_SLICE_X105Y106_CO6;
  assign CLBLM_L_X70Y107_SLICE_X105Y107_A5 = 1'b1;
  assign CLBLM_L_X70Y107_SLICE_X105Y107_A6 = CLBLM_L_X72Y108_SLICE_X108Y108_DQ;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_C5 = 1'b1;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_C6 = 1'b1;
  assign CLBLM_L_X70Y107_SLICE_X105Y107_B1 = CLBLL_R_X71Y107_SLICE_X106Y107_DO6;
  assign CLBLM_L_X70Y107_SLICE_X105Y107_B2 = CLBLM_L_X68Y109_SLICE_X103Y109_BQ;
  assign CLBLM_L_X70Y107_SLICE_X105Y107_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y107_SLICE_X105Y107_B4 = CLBLM_L_X68Y108_SLICE_X103Y108_CO6;
  assign CLBLM_L_X70Y107_SLICE_X105Y107_B5 = CLBLM_L_X70Y106_SLICE_X105Y106_CO6;
  assign CLBLM_L_X70Y107_SLICE_X105Y107_B6 = CLBLM_L_X68Y109_SLICE_X103Y109_B5Q;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_D1 = 1'b1;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_D2 = 1'b1;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_D3 = 1'b1;
  assign CLBLM_L_X70Y107_SLICE_X105Y107_C1 = 1'b1;
  assign CLBLM_L_X70Y107_SLICE_X105Y107_C2 = 1'b1;
  assign CLBLM_L_X70Y107_SLICE_X105Y107_C3 = 1'b1;
  assign CLBLM_L_X70Y108_SLICE_X104Y108_D5 = 1'b1;
  assign CLBLM_L_X70Y107_SLICE_X105Y107_C4 = 1'b1;
  assign CLBLM_L_X70Y107_SLICE_X105Y107_C5 = 1'b1;
  assign CLBLM_L_X70Y107_SLICE_X105Y107_C6 = 1'b1;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_A1 = CLBLM_L_X70Y105_SLICE_X105Y105_AQ;
  assign CLBLM_L_X70Y107_SLICE_X105Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_A2 = CLBLL_R_X75Y122_SLICE_X115Y122_AQ;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_A3 = CLBLM_L_X74Y121_SLICE_X113Y121_AQ;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_A4 = CLBLM_L_X74Y119_SLICE_X112Y119_BO6;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_A5 = CLBLL_R_X75Y121_SLICE_X114Y121_AQ;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_A6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y107_SLICE_X105Y107_D1 = 1'b1;
  assign CLBLM_L_X70Y107_SLICE_X105Y107_D2 = 1'b1;
  assign CLBLM_L_X70Y107_SLICE_X105Y107_D3 = 1'b1;
  assign CLBLM_L_X70Y107_SLICE_X105Y107_D4 = 1'b1;
  assign CLBLM_L_X70Y107_SLICE_X105Y107_D5 = 1'b1;
  assign CLBLM_L_X70Y107_SLICE_X105Y107_D6 = 1'b1;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_B1 = 1'b1;
  assign CLBLM_L_X70Y107_SLICE_X105Y107_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_B2 = CLBLM_R_X65Y105_SLICE_X99Y105_CQ;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_C1 = CLBLM_L_X74Y119_SLICE_X113Y119_AO6;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_C2 = CLBLM_L_X74Y119_SLICE_X112Y119_CQ;
  assign CLBLM_L_X70Y107_SLICE_X104Y107_A1 = CLBLM_L_X68Y107_SLICE_X103Y107_DO6;
  assign CLBLM_L_X70Y107_SLICE_X104Y107_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y107_SLICE_X104Y107_A3 = 1'b1;
  assign CLBLM_L_X70Y107_SLICE_X104Y107_A4 = CLBLM_L_X70Y106_SLICE_X104Y106_DO6;
  assign CLBLM_L_X70Y107_SLICE_X104Y107_A5 = CLBLM_L_X70Y106_SLICE_X104Y106_BQ;
  assign CLBLM_L_X70Y107_SLICE_X104Y107_A6 = CLBLM_L_X70Y107_SLICE_X104Y107_CO6;
  assign CLBLM_L_X70Y108_SLICE_X104Y108_D6 = 1'b1;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_C3 = CLBLM_L_X72Y118_SLICE_X108Y118_CQ;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_C4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_C5 = CLBLM_R_X65Y105_SLICE_X99Y105_CQ;
  assign CLBLM_L_X70Y107_SLICE_X104Y107_B1 = CLBLM_L_X68Y107_SLICE_X103Y107_DO6;
  assign CLBLM_L_X70Y107_SLICE_X104Y107_B2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y107_SLICE_X104Y107_B3 = CLBLM_L_X70Y107_SLICE_X104Y107_AQ;
  assign CLBLM_L_X70Y107_SLICE_X104Y107_B4 = CLBLM_L_X70Y106_SLICE_X104Y106_DO6;
  assign CLBLM_L_X70Y107_SLICE_X104Y107_B5 = CLBLM_L_X70Y106_SLICE_X104Y106_BQ;
  assign CLBLM_L_X70Y107_SLICE_X104Y107_B6 = CLBLM_L_X70Y107_SLICE_X104Y107_CO6;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_D1 = CLBLM_L_X74Y119_SLICE_X113Y119_AO6;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_D2 = CLBLM_L_X74Y119_SLICE_X112Y119_CQ;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_D3 = CLBLM_L_X74Y119_SLICE_X112Y119_DQ;
  assign CLBLM_L_X70Y107_SLICE_X104Y107_C1 = 1'b1;
  assign CLBLM_L_X70Y107_SLICE_X104Y107_C2 = CLBLM_L_X70Y107_SLICE_X105Y107_AQ;
  assign CLBLM_L_X70Y107_SLICE_X104Y107_C3 = CLBLM_L_X70Y106_SLICE_X105Y106_A5Q;
  assign CLBLM_L_X70Y107_SLICE_X104Y107_C4 = CLBLM_L_X70Y106_SLICE_X104Y106_A5Q;
  assign CLBLM_L_X70Y107_SLICE_X104Y107_C5 = CLBLM_L_X68Y109_SLICE_X103Y109_AQ;
  assign CLBLM_L_X70Y107_SLICE_X104Y107_C6 = CLBLM_L_X70Y105_SLICE_X104Y105_CO6;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_D6 = CLBLL_R_X75Y124_SLICE_X115Y124_BQ;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X70Y107_SLICE_X104Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_A6 = 1'b1;
  assign CLBLM_R_X65Y111_SLICE_X98Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X70Y107_SLICE_X104Y107_D1 = 1'b1;
  assign CLBLM_L_X70Y107_SLICE_X104Y107_D2 = 1'b1;
  assign CLBLM_L_X70Y107_SLICE_X104Y107_D3 = 1'b1;
  assign CLBLM_L_X70Y107_SLICE_X104Y107_D4 = 1'b1;
  assign CLBLM_L_X70Y107_SLICE_X104Y107_D5 = 1'b1;
  assign CLBLM_L_X70Y107_SLICE_X104Y107_D6 = 1'b1;
  assign CLBLM_L_X70Y107_SLICE_X104Y107_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign LIOB33_X0Y161_IOB_X0Y162_O = CLBLL_R_X71Y124_SLICE_X106Y124_AQ;
  assign LIOB33_X0Y161_IOB_X0Y161_O = CLBLM_L_X70Y110_SLICE_X104Y110_CQ;
  assign CLBLM_L_X82Y130_SLICE_X129Y130_B6 = 1'b1;
  assign CLBLM_R_X65Y111_SLICE_X98Y111_D4 = 1'b1;
  assign CLBLM_R_X65Y111_SLICE_X98Y111_D5 = 1'b1;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_B1 = CLBLM_L_X76Y126_SLICE_X116Y126_AO6;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_D1 = 1'b1;
  assign CLBLM_L_X82Y130_SLICE_X129Y130_A3 = 1'b1;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_B2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y121_SLICE_X118Y121_A1 = CLBLL_R_X77Y121_SLICE_X119Y121_DQ;
  assign CLBLL_R_X77Y121_SLICE_X118Y121_A2 = CLBLM_L_X76Y118_SLICE_X116Y118_DQ;
  assign CLBLL_R_X77Y121_SLICE_X118Y121_A3 = 1'b1;
  assign CLBLL_R_X77Y121_SLICE_X118Y121_A4 = CLBLM_L_X78Y123_SLICE_X121Y123_A5Q;
  assign CLBLL_R_X77Y121_SLICE_X118Y121_A5 = CLBLL_R_X77Y121_SLICE_X119Y121_AQ;
  assign CLBLL_R_X77Y121_SLICE_X118Y121_A6 = CLBLM_L_X76Y118_SLICE_X116Y118_AQ;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_B3 = CLBLM_L_X74Y123_SLICE_X112Y123_BQ;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_A1 = CLBLM_L_X76Y128_SLICE_X117Y128_B5Q;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_A2 = CLBLM_L_X76Y128_SLICE_X117Y128_BQ;
  assign CLBLL_R_X77Y121_SLICE_X118Y121_B1 = 1'b1;
  assign CLBLL_R_X77Y121_SLICE_X118Y121_B2 = 1'b1;
  assign CLBLL_R_X77Y121_SLICE_X118Y121_B3 = 1'b1;
  assign CLBLL_R_X77Y121_SLICE_X118Y121_B4 = 1'b1;
  assign CLBLL_R_X77Y121_SLICE_X118Y121_B5 = 1'b1;
  assign CLBLL_R_X77Y121_SLICE_X118Y121_B6 = 1'b1;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_A3 = 1'b1;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_A4 = CLBLL_R_X77Y129_SLICE_X118Y129_AQ;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_A5 = CLBLM_L_X76Y128_SLICE_X116Y128_CQ;
  assign CLBLL_R_X77Y121_SLICE_X118Y121_C1 = 1'b1;
  assign CLBLL_R_X77Y121_SLICE_X118Y121_C2 = 1'b1;
  assign CLBLL_R_X77Y121_SLICE_X118Y121_C3 = 1'b1;
  assign CLBLL_R_X77Y121_SLICE_X118Y121_C4 = 1'b1;
  assign CLBLL_R_X77Y121_SLICE_X118Y121_C5 = 1'b1;
  assign CLBLL_R_X77Y121_SLICE_X118Y121_C6 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_A1 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_A2 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_A3 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_A4 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_A5 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_A6 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_B1 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_B2 = 1'b1;
  assign CLBLL_R_X77Y121_SLICE_X118Y121_D1 = 1'b1;
  assign CLBLL_R_X77Y121_SLICE_X118Y121_D2 = 1'b1;
  assign CLBLL_R_X77Y121_SLICE_X118Y121_D3 = 1'b1;
  assign CLBLL_R_X77Y121_SLICE_X118Y121_D4 = 1'b1;
  assign CLBLL_R_X77Y121_SLICE_X118Y121_D5 = 1'b1;
  assign CLBLL_R_X77Y121_SLICE_X118Y121_D6 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_B3 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_B4 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_B5 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_B6 = 1'b1;
  assign CLBLM_L_X70Y108_SLICE_X105Y108_A1 = CLBLL_R_X71Y108_SLICE_X107Y108_A5Q;
  assign CLBLM_L_X70Y108_SLICE_X105Y108_A2 = CLBLM_L_X72Y118_SLICE_X109Y118_BQ;
  assign CLBLM_L_X70Y108_SLICE_X105Y108_A3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y108_SLICE_X105Y108_A4 = CLBLM_R_X65Y106_SLICE_X98Y106_CQ;
  assign CLBLM_L_X70Y108_SLICE_X105Y108_A5 = CLBLM_L_X74Y109_SLICE_X113Y109_A5Q;
  assign CLBLM_L_X70Y108_SLICE_X105Y108_A6 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_C2 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_C3 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_C5 = 1'b1;
  assign CLBLM_L_X70Y108_SLICE_X105Y108_B1 = 1'b1;
  assign CLBLM_L_X70Y108_SLICE_X105Y108_B2 = 1'b1;
  assign CLBLM_L_X70Y108_SLICE_X105Y108_B3 = 1'b1;
  assign CLBLM_L_X70Y108_SLICE_X105Y108_B4 = 1'b1;
  assign CLBLM_L_X70Y108_SLICE_X105Y108_B5 = 1'b1;
  assign CLBLM_L_X70Y108_SLICE_X105Y108_B6 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_D1 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_D2 = 1'b1;
  assign CLBLM_L_X70Y108_SLICE_X105Y108_C1 = 1'b1;
  assign CLBLM_L_X70Y108_SLICE_X105Y108_C2 = 1'b1;
  assign CLBLM_L_X70Y108_SLICE_X105Y108_C3 = 1'b1;
  assign CLBLM_L_X70Y108_SLICE_X105Y108_C4 = 1'b1;
  assign CLBLL_R_X77Y121_SLICE_X119Y121_A1 = CLBLL_R_X77Y121_SLICE_X119Y121_BO5;
  assign CLBLL_R_X77Y121_SLICE_X119Y121_A2 = CLBLL_R_X77Y122_SLICE_X119Y122_AO6;
  assign CLBLL_R_X77Y121_SLICE_X119Y121_A3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y121_SLICE_X119Y121_A4 = CLBLL_R_X77Y121_SLICE_X119Y121_BO6;
  assign CLBLL_R_X77Y121_SLICE_X119Y121_A5 = CLBLL_R_X77Y121_SLICE_X119Y121_DQ;
  assign CLBLL_R_X77Y121_SLICE_X119Y121_A6 = CLBLM_L_X78Y122_SLICE_X120Y122_DO6;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_A2 = CLBLM_L_X64Y97_SLICE_X97Y97_AQ;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_A3 = CLBLM_L_X64Y96_SLICE_X97Y96_AQ;
  assign CLBLM_L_X70Y108_SLICE_X105Y108_D1 = 1'b1;
  assign CLBLM_L_X70Y108_SLICE_X105Y108_D2 = 1'b1;
  assign CLBLM_L_X70Y108_SLICE_X105Y108_D3 = 1'b1;
  assign CLBLM_L_X70Y108_SLICE_X105Y108_D4 = 1'b1;
  assign CLBLM_L_X70Y108_SLICE_X105Y108_D5 = 1'b1;
  assign CLBLM_L_X70Y108_SLICE_X105Y108_D6 = 1'b1;
  assign CLBLL_R_X77Y121_SLICE_X119Y121_B1 = CLBLL_R_X77Y122_SLICE_X119Y122_DQ;
  assign CLBLL_R_X77Y121_SLICE_X119Y121_B2 = CLBLL_R_X77Y113_SLICE_X118Y113_AQ;
  assign CLBLL_R_X77Y121_SLICE_X119Y121_C2 = CLBLL_R_X77Y121_SLICE_X119Y121_CQ;
  assign CLBLL_R_X77Y121_SLICE_X119Y121_C3 = CLBLL_R_X77Y122_SLICE_X119Y122_DQ;
  assign CLBLL_R_X77Y121_SLICE_X119Y121_C4 = CLBLL_R_X77Y122_SLICE_X119Y122_CQ;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_B6 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_C1 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_C2 = 1'b1;
  assign CLBLL_R_X77Y121_SLICE_X119Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_C3 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_C4 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_C5 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_C6 = 1'b1;
  assign CLBLL_R_X77Y121_SLICE_X119Y121_D1 = CLBLM_L_X78Y123_SLICE_X121Y123_CO6;
  assign CLBLL_R_X77Y121_SLICE_X119Y121_D2 = CLBLL_R_X77Y121_SLICE_X119Y121_CQ;
  assign CLBLL_R_X77Y121_SLICE_X119Y121_D3 = CLBLL_R_X77Y121_SLICE_X119Y121_DQ;
  assign CLBLL_R_X77Y121_SLICE_X119Y121_D4 = CLBLM_L_X78Y122_SLICE_X120Y122_DO6;
  assign CLBLL_R_X77Y121_SLICE_X119Y121_D5 = CLBLL_R_X77Y121_SLICE_X119Y121_BO5;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_D1 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_D2 = 1'b1;
  assign CLBLL_R_X77Y121_SLICE_X119Y121_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_D3 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_D4 = 1'b1;
  assign CLBLM_L_X70Y108_SLICE_X104Y108_C2 = 1'b1;
  assign CLBLM_L_X70Y108_SLICE_X104Y108_C3 = 1'b1;
  assign CLBLM_L_X70Y108_SLICE_X104Y108_C4 = 1'b1;
  assign CLBLM_L_X70Y108_SLICE_X104Y108_C5 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_A1 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_A2 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_A3 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_A4 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_A5 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_B1 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_B2 = 1'b1;
  assign CLBLM_L_X70Y108_SLICE_X104Y108_D1 = 1'b1;
  assign CLBLM_L_X70Y108_SLICE_X104Y108_D2 = 1'b1;
  assign CLBLM_L_X70Y108_SLICE_X104Y108_D3 = 1'b1;
  assign CLBLM_L_X70Y108_SLICE_X104Y108_D4 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_B3 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_B4 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_B5 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_C1 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_C2 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_B6 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_C3 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_C4 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_C5 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_C6 = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_T1 = 1'b1;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_D1 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_D2 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_D3 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_D4 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_D5 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_D6 = 1'b1;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_A1 = CLBLM_L_X72Y121_SLICE_X108Y121_CQ;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_A2 = CLBLM_L_X72Y121_SLICE_X108Y121_DQ;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_A3 = CLBLM_L_X76Y119_SLICE_X116Y119_AQ;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_A4 = CLBLM_L_X72Y121_SLICE_X109Y121_A5Q;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_A5 = CLBLM_L_X72Y121_SLICE_X109Y121_AQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1 = 1'b1;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_A6 = 1'b1;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_AX = CLBLM_L_X72Y121_SLICE_X108Y121_DQ;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_B1 = CLBLM_L_X72Y122_SLICE_X108Y122_CQ;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_B2 = CLBLM_L_X72Y121_SLICE_X108Y121_BQ;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_B3 = CLBLM_L_X74Y122_SLICE_X112Y122_BQ;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_B4 = CLBLM_L_X72Y118_SLICE_X108Y118_AQ;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_B5 = CLBLM_L_X72Y128_SLICE_X109Y128_AQ;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_B6 = CLBLM_L_X72Y121_SLICE_X108Y121_A5Q;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1 = 1'b1;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_BX = CLBLM_L_X72Y120_SLICE_X108Y120_A5Q;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_C1 = 1'b1;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_C2 = 1'b1;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_C3 = 1'b1;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_C4 = 1'b1;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_C5 = 1'b1;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_A1 = CLBLM_L_X76Y122_SLICE_X117Y122_AQ;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_A2 = CLBLM_L_X78Y122_SLICE_X120Y122_BO6;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_A3 = CLBLL_R_X77Y122_SLICE_X118Y122_AQ;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_A4 = CLBLL_R_X77Y113_SLICE_X118Y113_AQ;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_A6 = CLBLM_L_X78Y122_SLICE_X121Y122_BQ;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_C6 = 1'b1;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_CE = CLBLM_L_X76Y109_SLICE_X116Y109_AO6;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_B1 = CLBLM_L_X76Y122_SLICE_X117Y122_AQ;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_B2 = CLBLL_R_X77Y122_SLICE_X118Y122_BQ;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_B3 = CLBLL_R_X77Y122_SLICE_X118Y122_AQ;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_B4 = CLBLL_R_X77Y113_SLICE_X118Y113_AQ;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_B5 = CLBLM_L_X78Y122_SLICE_X120Y122_BO6;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_B6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X76Y129_SLICE_X117Y129_A1 = 1'b1;
  assign CLBLM_L_X76Y129_SLICE_X117Y129_A2 = 1'b1;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_C5 = CLBLL_R_X77Y127_SLICE_X119Y127_AQ;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_C1 = CLBLL_R_X77Y121_SLICE_X118Y121_AO6;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_C2 = CLBLL_R_X75Y123_SLICE_X114Y123_AO6;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_C3 = 1'b1;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_C4 = CLBLM_L_X76Y125_SLICE_X117Y125_BQ;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_C5 = CLBLM_L_X78Y123_SLICE_X120Y123_DO6;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_C6 = CLBLL_R_X75Y123_SLICE_X115Y123_CO6;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_A2 = CLBLM_L_X76Y122_SLICE_X116Y122_CQ;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_A3 = 1'b1;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_A4 = CLBLM_L_X74Y123_SLICE_X112Y123_B5Q;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_A5 = CLBLM_L_X74Y121_SLICE_X113Y121_A5Q;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_A6 = 1'b1;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_D1 = 1'b1;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_D2 = 1'b1;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_D3 = 1'b1;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_D4 = 1'b1;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_D5 = 1'b1;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_D6 = 1'b1;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_B1 = CLBLM_L_X74Y121_SLICE_X113Y121_B5Q;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_CX = CLBLM_L_X72Y121_SLICE_X108Y121_BQ;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_B2 = CLBLM_L_X74Y121_SLICE_X113Y121_BQ;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_B4 = CLBLM_L_X74Y123_SLICE_X112Y123_B5Q;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_B5 = CLBLM_L_X74Y121_SLICE_X113Y121_A5Q;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_B6 = 1'b1;
  assign CLBLM_L_X70Y109_SLICE_X105Y109_A1 = 1'b1;
  assign CLBLM_L_X70Y109_SLICE_X105Y109_A2 = 1'b1;
  assign CLBLM_L_X70Y109_SLICE_X105Y109_A3 = 1'b1;
  assign CLBLM_L_X70Y109_SLICE_X105Y109_A4 = 1'b1;
  assign CLBLM_L_X70Y109_SLICE_X105Y109_A5 = 1'b1;
  assign CLBLM_L_X70Y109_SLICE_X105Y109_A6 = 1'b1;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_D1 = 1'b1;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_C3 = 1'b1;
  assign CLBLM_L_X70Y109_SLICE_X105Y109_AX = CLBLM_L_X70Y109_SLICE_X104Y109_B5Q;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_D2 = 1'b1;
  assign CLBLM_L_X70Y109_SLICE_X105Y109_B1 = 1'b1;
  assign CLBLM_L_X70Y109_SLICE_X105Y109_B2 = 1'b1;
  assign CLBLM_L_X70Y109_SLICE_X105Y109_B3 = 1'b1;
  assign CLBLM_L_X70Y109_SLICE_X105Y109_B4 = 1'b1;
  assign CLBLM_L_X70Y109_SLICE_X105Y109_B5 = 1'b1;
  assign CLBLM_L_X70Y109_SLICE_X105Y109_B6 = 1'b1;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_D3 = 1'b1;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_A1 = CLBLL_R_X77Y122_SLICE_X118Y122_AQ;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_A2 = CLBLL_R_X77Y113_SLICE_X118Y113_AQ;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_A3 = CLBLM_L_X76Y122_SLICE_X117Y122_AQ;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_A4 = CLBLL_R_X77Y122_SLICE_X118Y122_BQ;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_A5 = CLBLL_R_X77Y121_SLICE_X119Y121_CQ;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_A6 = 1'b1;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_A1 = CLBLM_R_X63Y98_SLICE_X94Y98_AO5;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_A3 = CLBLM_L_X64Y96_SLICE_X97Y96_AQ;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_B1 = CLBLL_R_X77Y122_SLICE_X118Y122_AQ;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_B2 = CLBLL_R_X77Y122_SLICE_X119Y122_BQ;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_B4 = CLBLL_R_X77Y122_SLICE_X118Y122_BQ;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_B5 = CLBLM_L_X78Y122_SLICE_X120Y122_BO6;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_B6 = CLBLM_L_X78Y123_SLICE_X121Y123_CO6;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_A6 = 1'b1;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_B3 = 1'b1;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_B4 = 1'b1;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_C1 = CLBLL_R_X77Y113_SLICE_X118Y113_AQ;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_C2 = CLBLL_R_X77Y122_SLICE_X119Y122_CQ;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_C3 = CLBLM_L_X76Y122_SLICE_X117Y122_AQ;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_C4 = CLBLL_R_X77Y122_SLICE_X119Y122_BQ;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_C5 = CLBLM_L_X78Y122_SLICE_X120Y122_CO6;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_C6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_B6 = 1'b1;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_C1 = CLBLM_L_X64Y98_SLICE_X96Y98_AO6;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_C2 = CLBLM_L_X64Y97_SLICE_X97Y97_CQ;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_C5 = CLBLM_R_X63Y99_SLICE_X94Y99_A5Q;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_C6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_D1 = CLBLL_R_X77Y122_SLICE_X119Y122_DQ;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_D2 = CLBLL_R_X77Y122_SLICE_X119Y122_CQ;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_D3 = CLBLL_R_X77Y122_SLICE_X119Y122_BQ;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_D4 = CLBLM_L_X78Y123_SLICE_X121Y123_CO6;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_D5 = CLBLM_L_X78Y122_SLICE_X120Y122_CO6;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_D6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_D1 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_D2 = CLBLM_L_X64Y98_SLICE_X96Y98_AO6;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_D3 = CLBLM_L_X64Y97_SLICE_X97Y97_DQ;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_D4 = CLBLM_R_X63Y96_SLICE_X95Y96_DQ;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_D5 = CLBLM_R_X63Y99_SLICE_X94Y99_CO5;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_D6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X70Y109_SLICE_X104Y109_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_A1 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_A2 = CLBLM_R_X63Y99_SLICE_X94Y99_BO6;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_A3 = CLBLM_L_X64Y97_SLICE_X96Y97_AQ;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_A4 = CLBLM_L_X64Y99_SLICE_X96Y99_BQ;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_A5 = CLBLM_L_X64Y99_SLICE_X96Y99_A5Q;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_A6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y109_SLICE_X104Y109_C1 = 1'b1;
  assign CLBLM_L_X70Y109_SLICE_X104Y109_C2 = 1'b1;
  assign CLBLM_L_X70Y109_SLICE_X104Y109_C3 = 1'b1;
  assign CLBLM_L_X70Y109_SLICE_X104Y109_C4 = 1'b1;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_B1 = CLBLM_R_X63Y99_SLICE_X94Y99_A5Q;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_B2 = CLBLM_L_X64Y97_SLICE_X96Y97_BQ;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_B3 = CLBLM_L_X64Y97_SLICE_X97Y97_BO5;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_B4 = CLBLM_L_X64Y97_SLICE_X96Y97_DQ;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_B5 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_B6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y109_SLICE_X104Y109_D1 = 1'b1;
  assign CLBLM_L_X70Y109_SLICE_X104Y109_D2 = 1'b1;
  assign CLBLM_L_X70Y109_SLICE_X104Y109_D3 = 1'b1;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_C1 = CLBLM_R_X63Y99_SLICE_X94Y99_BO6;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_C2 = CLBLM_L_X64Y97_SLICE_X96Y97_CQ;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_C3 = CLBLM_R_X63Y97_SLICE_X94Y97_BQ;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_C4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_C5 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_C6 = CLBLM_L_X64Y98_SLICE_X96Y98_AO6;
  assign CLBLM_L_X70Y109_SLICE_X104Y109_D6 = 1'b1;
  assign CLBLM_L_X70Y109_SLICE_X104Y109_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign RIOI3_X105Y147_OLOGIC_X1Y148_D1 = CLBLM_L_X62Y103_SLICE_X92Y103_B5Q;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_D1 = RIOB33_X105Y55_IOB_X1Y56_I;
  assign RIOI3_X105Y147_OLOGIC_X1Y148_T1 = 1'b1;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_D1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_D2 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_D3 = CLBLM_L_X64Y97_SLICE_X97Y97_BO5;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_D4 = CLBLM_L_X64Y97_SLICE_X96Y97_DQ;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_D5 = CLBLM_R_X63Y99_SLICE_X94Y99_CO5;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_D6 = CLBLM_R_X63Y96_SLICE_X95Y96_CQ;
  assign LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y88_D1 = CLBLM_L_X60Y94_SLICE_X90Y94_CQ;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_T1 = 1'b1;
  assign CLBLL_R_X79Y127_SLICE_X122Y127_C4 = CLBLL_R_X83Y130_SLICE_X130Y130_CQ;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign RIOI3_X105Y147_OLOGIC_X1Y147_D1 = CLBLL_R_X77Y108_SLICE_X118Y108_AQ;
  assign LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y88_T1 = 1'b1;
  assign RIOI3_X105Y147_OLOGIC_X1Y147_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y87_D1 = CLBLM_R_X63Y97_SLICE_X94Y97_B5Q;
  assign LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y87_T1 = 1'b1;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_A5 = CLBLM_L_X64Y102_SLICE_X96Y102_AQ;
  assign CLBLM_L_X76Y134_SLICE_X117Y134_D1 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X118Y104_B3 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X118Y104_B4 = 1'b1;
  assign CLBLL_R_X77Y123_SLICE_X118Y123_A1 = CLBLL_R_X77Y124_SLICE_X118Y124_DO6;
  assign CLBLL_R_X77Y123_SLICE_X118Y123_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y123_SLICE_X118Y123_A3 = CLBLL_R_X77Y123_SLICE_X118Y123_AQ;
  assign CLBLL_R_X77Y123_SLICE_X118Y123_A4 = CLBLL_R_X77Y123_SLICE_X118Y123_BO6;
  assign CLBLL_R_X77Y123_SLICE_X118Y123_A5 = CLBLL_R_X77Y123_SLICE_X119Y123_AQ;
  assign CLBLL_R_X77Y123_SLICE_X118Y123_A6 = CLBLM_L_X78Y124_SLICE_X120Y124_CQ;
  assign CLBLL_R_X77Y123_SLICE_X118Y123_B1 = CLBLM_L_X76Y123_SLICE_X117Y123_AQ;
  assign CLBLL_R_X77Y123_SLICE_X118Y123_B2 = CLBLM_L_X74Y123_SLICE_X113Y123_A5Q;
  assign CLBLL_R_X77Y123_SLICE_X118Y123_B3 = CLBLL_R_X75Y113_SLICE_X114Y113_AQ;
  assign CLBLL_R_X77Y123_SLICE_X118Y123_B4 = CLBLM_L_X78Y124_SLICE_X120Y124_CQ;
  assign CLBLL_R_X77Y123_SLICE_X118Y123_B5 = CLBLL_R_X77Y123_SLICE_X119Y123_AQ;
  assign CLBLL_R_X77Y123_SLICE_X118Y123_B6 = 1'b1;
  assign CLBLM_L_X76Y130_SLICE_X117Y130_A1 = 1'b1;
  assign CLBLM_L_X76Y130_SLICE_X117Y130_A2 = 1'b1;
  assign CLBLM_L_X76Y130_SLICE_X117Y130_A3 = 1'b1;
  assign CLBLL_R_X77Y123_SLICE_X118Y123_C1 = CLBLM_L_X76Y123_SLICE_X117Y123_AO5;
  assign CLBLL_R_X77Y123_SLICE_X118Y123_C2 = CLBLL_R_X77Y123_SLICE_X118Y123_CQ;
  assign CLBLL_R_X77Y123_SLICE_X118Y123_C3 = CLBLL_R_X77Y123_SLICE_X118Y123_AQ;
  assign CLBLL_R_X77Y123_SLICE_X118Y123_C4 = CLBLL_R_X77Y123_SLICE_X119Y123_CQ;
  assign CLBLL_R_X77Y123_SLICE_X118Y123_C5 = CLBLM_L_X76Y124_SLICE_X117Y124_BQ;
  assign CLBLL_R_X77Y123_SLICE_X118Y123_C6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X76Y130_SLICE_X117Y130_A4 = 1'b1;
  assign CLBLM_L_X76Y130_SLICE_X117Y130_A5 = 1'b1;
  assign CLBLL_R_X77Y123_SLICE_X118Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X76Y130_SLICE_X117Y130_A6 = 1'b1;
  assign CLBLM_L_X76Y130_SLICE_X117Y130_B1 = 1'b1;
  assign CLBLM_L_X74Y122_SLICE_X113Y122_A1 = CLBLL_R_X75Y123_SLICE_X114Y123_BQ;
  assign CLBLM_L_X74Y122_SLICE_X113Y122_A2 = CLBLM_L_X74Y123_SLICE_X113Y123_CO5;
  assign CLBLL_R_X77Y123_SLICE_X118Y123_D1 = CLBLM_L_X78Y124_SLICE_X120Y124_BQ;
  assign CLBLL_R_X77Y123_SLICE_X118Y123_D2 = CLBLL_R_X77Y123_SLICE_X118Y123_CQ;
  assign CLBLL_R_X77Y123_SLICE_X118Y123_D3 = CLBLL_R_X77Y124_SLICE_X118Y124_BQ;
  assign CLBLL_R_X77Y123_SLICE_X118Y123_D4 = CLBLM_L_X78Y124_SLICE_X120Y124_AQ;
  assign CLBLL_R_X77Y123_SLICE_X118Y123_D5 = CLBLM_L_X74Y123_SLICE_X113Y123_CO5;
  assign CLBLL_R_X77Y123_SLICE_X118Y123_D6 = CLBLL_R_X77Y123_SLICE_X118Y123_AQ;
  assign CLBLM_L_X74Y122_SLICE_X113Y122_A3 = CLBLM_L_X74Y122_SLICE_X113Y122_AQ;
  assign CLBLM_L_X74Y122_SLICE_X113Y122_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y123_SLICE_X118Y123_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y122_SLICE_X113Y122_A5 = CLBLM_L_X74Y123_SLICE_X113Y123_DQ;
  assign CLBLM_L_X74Y122_SLICE_X113Y122_A6 = CLBLL_R_X75Y121_SLICE_X114Y121_AO5;
  assign CLBLM_L_X74Y122_SLICE_X113Y122_B1 = 1'b1;
  assign CLBLM_L_X74Y122_SLICE_X113Y122_B2 = 1'b1;
  assign CLBLM_L_X74Y122_SLICE_X113Y122_B3 = 1'b1;
  assign CLBLM_L_X74Y122_SLICE_X113Y122_B4 = 1'b1;
  assign CLBLM_L_X74Y122_SLICE_X113Y122_C1 = 1'b1;
  assign CLBLM_L_X74Y122_SLICE_X113Y122_C2 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X118Y104_C5 = 1'b1;
  assign CLBLM_L_X74Y122_SLICE_X113Y122_C3 = 1'b1;
  assign CLBLM_L_X70Y110_SLICE_X105Y110_A1 = 1'b1;
  assign CLBLM_L_X70Y110_SLICE_X105Y110_A2 = 1'b1;
  assign CLBLM_L_X70Y110_SLICE_X105Y110_A3 = 1'b1;
  assign CLBLM_L_X70Y110_SLICE_X105Y110_A4 = 1'b1;
  assign CLBLM_L_X70Y110_SLICE_X105Y110_A5 = 1'b1;
  assign CLBLM_L_X70Y110_SLICE_X105Y110_A6 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X118Y104_C6 = 1'b1;
  assign CLBLM_L_X74Y122_SLICE_X113Y122_C4 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X118Y104_CE = CLBLM_L_X76Y109_SLICE_X116Y109_AO6;
  assign CLBLM_L_X70Y110_SLICE_X105Y110_B1 = 1'b1;
  assign CLBLM_L_X70Y110_SLICE_X105Y110_B2 = 1'b1;
  assign CLBLM_L_X70Y110_SLICE_X105Y110_B3 = 1'b1;
  assign CLBLM_L_X70Y110_SLICE_X105Y110_B4 = 1'b1;
  assign CLBLL_R_X77Y123_SLICE_X119Y123_A1 = CLBLL_R_X77Y123_SLICE_X119Y123_CQ;
  assign CLBLL_R_X77Y123_SLICE_X119Y123_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y123_SLICE_X119Y123_A3 = CLBLL_R_X77Y123_SLICE_X119Y123_AQ;
  assign CLBLL_R_X77Y123_SLICE_X119Y123_A4 = CLBLM_L_X76Y123_SLICE_X117Y123_AO5;
  assign CLBLL_R_X77Y123_SLICE_X119Y123_A5 = CLBLM_L_X76Y124_SLICE_X117Y124_BQ;
  assign CLBLL_R_X77Y123_SLICE_X119Y123_A6 = CLBLL_R_X77Y123_SLICE_X118Y123_CQ;
  assign CLBLM_L_X70Y110_SLICE_X105Y110_C1 = 1'b1;
  assign CLBLM_L_X70Y110_SLICE_X105Y110_C2 = 1'b1;
  assign CLBLL_R_X77Y123_SLICE_X119Y123_B1 = CLBLM_L_X78Y124_SLICE_X120Y124_CQ;
  assign CLBLL_R_X77Y123_SLICE_X119Y123_B2 = CLBLL_R_X77Y124_SLICE_X118Y124_AO5;
  assign CLBLL_R_X77Y123_SLICE_X119Y123_B3 = CLBLL_R_X75Y123_SLICE_X114Y123_AO6;
  assign CLBLL_R_X77Y123_SLICE_X119Y123_B4 = CLBLL_R_X77Y121_SLICE_X118Y121_AO6;
  assign CLBLL_R_X77Y123_SLICE_X119Y123_B5 = CLBLL_R_X77Y123_SLICE_X118Y123_AQ;
  assign CLBLL_R_X77Y123_SLICE_X119Y123_B6 = 1'b1;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_A1 = 1'b1;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_A2 = 1'b1;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_A3 = 1'b1;
  assign CLBLL_R_X77Y123_SLICE_X119Y123_C1 = CLBLM_L_X76Y123_SLICE_X117Y123_AO5;
  assign CLBLL_R_X77Y123_SLICE_X119Y123_C2 = CLBLM_L_X76Y125_SLICE_X117Y125_BQ;
  assign CLBLL_R_X77Y123_SLICE_X119Y123_C3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y123_SLICE_X119Y123_C4 = CLBLL_R_X75Y122_SLICE_X114Y122_AQ;
  assign CLBLL_R_X77Y123_SLICE_X119Y123_C5 = CLBLL_R_X77Y123_SLICE_X119Y123_CQ;
  assign CLBLL_R_X77Y123_SLICE_X119Y123_C6 = CLBLM_L_X76Y119_SLICE_X116Y119_BO6;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_B1 = 1'b1;
  assign CLBLL_R_X77Y123_SLICE_X119Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_B2 = 1'b1;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_B3 = 1'b1;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_B4 = 1'b1;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_B5 = 1'b1;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_B6 = 1'b1;
  assign CLBLL_R_X77Y123_SLICE_X119Y123_D1 = CLBLL_R_X75Y123_SLICE_X114Y123_AO6;
  assign CLBLL_R_X77Y123_SLICE_X119Y123_D2 = CLBLL_R_X77Y121_SLICE_X118Y121_AO6;
  assign CLBLL_R_X77Y123_SLICE_X119Y123_D3 = CLBLL_R_X77Y124_SLICE_X118Y124_AO5;
  assign CLBLL_R_X77Y123_SLICE_X119Y123_D4 = CLBLM_L_X76Y125_SLICE_X117Y125_BQ;
  assign CLBLL_R_X77Y123_SLICE_X119Y123_D5 = CLBLL_R_X77Y123_SLICE_X118Y123_AQ;
  assign CLBLL_R_X77Y123_SLICE_X119Y123_D6 = CLBLM_L_X78Y124_SLICE_X120Y124_CQ;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_C3 = 1'b1;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_C4 = 1'b1;
  assign CLBLL_R_X77Y123_SLICE_X119Y123_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X70Y110_SLICE_X104Y110_B1 = CLBLM_L_X70Y110_SLICE_X104Y110_B5Q;
  assign CLBLM_L_X70Y110_SLICE_X104Y110_B2 = CLBLM_L_X70Y110_SLICE_X104Y110_BQ;
  assign CLBLM_L_X70Y110_SLICE_X104Y110_B4 = CLBLM_L_X70Y111_SLICE_X104Y111_CO6;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_D1 = 1'b1;
  assign CLBLM_L_X70Y110_SLICE_X104Y110_B6 = 1'b1;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_D2 = 1'b1;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_D3 = 1'b1;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_D4 = 1'b1;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_D5 = 1'b1;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_D6 = 1'b1;
  assign CLBLM_L_X70Y110_SLICE_X104Y110_C2 = CLBLM_L_X70Y110_SLICE_X104Y110_AQ;
  assign CLBLM_L_X70Y110_SLICE_X104Y110_C3 = CLBLM_L_X70Y112_SLICE_X104Y112_A5Q;
  assign CLBLM_L_X70Y110_SLICE_X104Y110_C4 = CLBLM_L_X70Y110_SLICE_X104Y110_BQ;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_A1 = CLBLM_L_X64Y99_SLICE_X96Y99_A5Q;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_A4 = 1'b1;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_A5 = 1'b1;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_A6 = 1'b1;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_A2 = CLBLM_L_X64Y99_SLICE_X96Y99_BQ;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_A3 = 1'b1;
  assign CLBLM_L_X70Y110_SLICE_X104Y110_C5 = CLBLM_L_X70Y110_SLICE_X104Y110_B5Q;
  assign CLBLM_L_X70Y110_SLICE_X104Y110_C6 = CLBLL_R_X71Y111_SLICE_X107Y111_BO6;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_B2 = CLBLM_L_X64Y98_SLICE_X96Y98_BQ;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_B3 = CLBLM_L_X64Y97_SLICE_X97Y97_CQ;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_B4 = CLBLM_R_X63Y99_SLICE_X94Y99_BO6;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_B5 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_B6 = CLBLM_L_X64Y98_SLICE_X96Y98_AO5;
  assign CLBLM_L_X70Y110_SLICE_X104Y110_D1 = 1'b1;
  assign CLBLM_L_X70Y110_SLICE_X104Y110_D2 = 1'b1;
  assign CLBLM_L_X70Y110_SLICE_X104Y110_D3 = 1'b1;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_C1 = CLBLM_L_X62Y99_SLICE_X93Y99_AQ;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_C2 = CLBLM_R_X63Y97_SLICE_X94Y97_AQ;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_C3 = CLBLM_R_X63Y96_SLICE_X95Y96_CQ;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_C4 = CLBLM_L_X76Y111_SLICE_X116Y111_BQ;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_C5 = CLBLM_L_X64Y97_SLICE_X97Y97_A5Q;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_C6 = CLBLM_R_X63Y96_SLICE_X94Y96_BQ;
  assign CLBLM_L_X70Y110_SLICE_X104Y110_D6 = 1'b1;
  assign CLBLM_L_X70Y110_SLICE_X104Y110_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_D1 = 1'b1;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_D2 = 1'b1;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_D3 = 1'b1;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_D4 = 1'b1;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_D5 = 1'b1;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_D6 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X95Y122_A1 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X95Y122_A2 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X95Y122_A3 = 1'b1;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X63Y122_SLICE_X95Y122_A4 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X95Y122_A5 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X95Y122_A6 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X95Y122_B5 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X95Y122_B6 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X95Y122_AX = CLBLM_L_X64Y122_SLICE_X96Y122_AQ;
  assign CLBLM_R_X63Y122_SLICE_X95Y122_B1 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X95Y122_B2 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X95Y122_C1 = 1'b1;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_D2 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X95Y122_C2 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X95Y122_C3 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X95Y122_C4 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_A4 = CLBLM_L_X64Y99_SLICE_X97Y99_A5Q;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_D3 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X95Y122_C5 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X95Y122_C6 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X95Y122_CE = CLBLM_L_X76Y109_SLICE_X116Y109_AO6;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_A5 = 1'b1;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_D4 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X95Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X63Y122_SLICE_X95Y122_CX = CLBLM_R_X53Y122_SLICE_X80Y122_AQ;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_A6 = CLBLM_L_X64Y96_SLICE_X97Y96_A5Q;
  assign CLBLM_R_X63Y122_SLICE_X95Y122_D1 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X95Y122_D2 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X95Y122_D3 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X95Y122_D4 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X95Y122_D5 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X95Y122_D6 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X95Y122_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X63Y122_SLICE_X94Y122_A1 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X94Y122_A2 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_AX = CLBLM_L_X64Y99_SLICE_X97Y99_A5Q;
  assign CLBLM_R_X63Y122_SLICE_X94Y122_A3 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X94Y122_A4 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X94Y122_A5 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X94Y122_A6 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X94Y122_B1 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_B1 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X94Y122_B2 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X94Y122_B3 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X94Y122_B4 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X94Y122_B5 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_B2 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X94Y122_B6 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_B3 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X94Y122_C1 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X94Y122_C2 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X94Y122_C3 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X94Y122_C4 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_B4 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X94Y122_C5 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X94Y122_C6 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_B5 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X94Y122_D1 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X94Y122_D2 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X94Y122_D3 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X94Y122_D4 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X94Y122_D5 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X94Y122_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1 = 1'b1;
  assign CLBLL_R_X77Y124_SLICE_X118Y124_A1 = CLBLL_R_X77Y125_SLICE_X118Y125_CQ;
  assign CLBLL_R_X77Y124_SLICE_X118Y124_A2 = CLBLL_R_X77Y124_SLICE_X118Y124_BQ;
  assign CLBLL_R_X77Y124_SLICE_X118Y124_A3 = CLBLM_L_X76Y123_SLICE_X116Y123_AQ;
  assign CLBLL_R_X77Y124_SLICE_X118Y124_A4 = CLBLM_L_X78Y124_SLICE_X120Y124_AQ;
  assign CLBLL_R_X77Y124_SLICE_X118Y124_A5 = CLBLM_L_X78Y124_SLICE_X120Y124_BQ;
  assign CLBLL_R_X77Y124_SLICE_X118Y124_A6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_D1 = CLBLL_R_X77Y129_SLICE_X118Y129_AQ;
  assign CLBLL_R_X77Y124_SLICE_X118Y124_B1 = CLBLL_R_X77Y123_SLICE_X118Y123_BO5;
  assign CLBLL_R_X77Y124_SLICE_X118Y124_B2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y124_SLICE_X118Y124_B3 = CLBLL_R_X77Y126_SLICE_X118Y126_AO5;
  assign CLBLL_R_X77Y124_SLICE_X118Y124_B4 = CLBLM_L_X78Y124_SLICE_X120Y124_CQ;
  assign CLBLL_R_X77Y124_SLICE_X118Y124_B5 = CLBLL_R_X77Y124_SLICE_X118Y124_BQ;
  assign CLBLL_R_X77Y124_SLICE_X118Y124_B6 = CLBLL_R_X77Y124_SLICE_X118Y124_CO6;
  assign CLBLM_L_X76Y123_SLICE_X117Y123_D6 = CLBLL_R_X75Y123_SLICE_X114Y123_AO6;
  assign CLBLL_R_X77Y124_SLICE_X118Y124_C1 = CLBLM_L_X78Y124_SLICE_X120Y124_BQ;
  assign CLBLL_R_X77Y124_SLICE_X118Y124_C2 = CLBLM_L_X78Y124_SLICE_X120Y124_CQ;
  assign CLBLL_R_X77Y124_SLICE_X118Y124_C3 = CLBLM_L_X78Y124_SLICE_X120Y124_AQ;
  assign CLBLL_R_X77Y124_SLICE_X118Y124_C4 = CLBLL_R_X77Y124_SLICE_X118Y124_BQ;
  assign CLBLL_R_X77Y124_SLICE_X118Y124_C5 = CLBLL_R_X77Y123_SLICE_X119Y123_AQ;
  assign CLBLL_R_X77Y124_SLICE_X118Y124_C6 = CLBLL_R_X77Y123_SLICE_X118Y123_BO6;
  assign CLBLL_R_X77Y124_SLICE_X118Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X76Y123_SLICE_X117Y123_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X77Y124_SLICE_X118Y124_D1 = CLBLM_L_X76Y124_SLICE_X117Y124_BQ;
  assign CLBLL_R_X77Y124_SLICE_X118Y124_D2 = 1'b1;
  assign CLBLL_R_X77Y124_SLICE_X118Y124_D3 = 1'b1;
  assign CLBLL_R_X77Y124_SLICE_X118Y124_D4 = CLBLL_R_X77Y123_SLICE_X119Y123_CQ;
  assign CLBLL_R_X77Y124_SLICE_X118Y124_D5 = 1'b1;
  assign CLBLL_R_X77Y124_SLICE_X118Y124_D6 = 1'b1;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_A1 = CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_A2 = CLBLL_R_X73Y125_SLICE_X111Y125_AQ;
  assign CLBLL_R_X77Y124_SLICE_X118Y124_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_A3 = CLBLM_L_X74Y123_SLICE_X113Y123_AQ;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_A5 = CLBLL_R_X75Y123_SLICE_X115Y123_BO6;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_A6 = 1'b1;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_AX = CLBLM_L_X74Y123_SLICE_X113Y123_CO6;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_B2 = CLBLM_L_X74Y123_SLICE_X113Y123_BQ;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_B3 = CLBLM_L_X74Y109_SLICE_X113Y109_AQ;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_B4 = CLBLM_L_X76Y123_SLICE_X117Y123_AQ;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_B5 = CLBLL_R_X75Y113_SLICE_X114Y113_AQ;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_B6 = CLBLM_L_X74Y123_SLICE_X113Y123_A5Q;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_C1 = CLBLM_L_X76Y123_SLICE_X117Y123_AQ;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_C2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_C3 = CLBLM_L_X74Y123_SLICE_X113Y123_BQ;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_C4 = CLBLM_L_X74Y123_SLICE_X113Y123_A5Q;
  assign CLBLM_L_X70Y111_SLICE_X105Y111_A1 = CLBLL_R_X71Y111_SLICE_X106Y111_CQ;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_D5 = 1'b1;
  assign CLBLM_L_X70Y111_SLICE_X105Y111_A2 = CLBLM_L_X70Y111_SLICE_X105Y111_BQ;
  assign CLBLM_L_X70Y111_SLICE_X105Y111_A3 = CLBLM_L_X70Y111_SLICE_X105Y111_AQ;
  assign CLBLM_L_X70Y111_SLICE_X105Y111_A4 = CLBLM_L_X70Y111_SLICE_X104Y111_BO5;
  assign CLBLM_L_X70Y111_SLICE_X105Y111_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_D6 = 1'b1;
  assign CLBLM_L_X70Y111_SLICE_X105Y111_A6 = CLBLL_R_X71Y111_SLICE_X106Y111_BQ;
  assign CLBLL_R_X77Y124_SLICE_X119Y124_A1 = CLBLL_R_X77Y124_SLICE_X119Y124_AQ;
  assign CLBLM_L_X70Y111_SLICE_X105Y111_B1 = 1'b1;
  assign CLBLL_R_X77Y124_SLICE_X119Y124_A2 = CLBLL_R_X77Y123_SLICE_X118Y123_DO6;
  assign CLBLL_R_X77Y124_SLICE_X119Y124_A3 = CLBLM_L_X76Y124_SLICE_X117Y124_BQ;
  assign CLBLL_R_X77Y124_SLICE_X119Y124_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y124_SLICE_X119Y124_A5 = CLBLM_L_X76Y119_SLICE_X116Y119_BO6;
  assign CLBLL_R_X77Y124_SLICE_X119Y124_A6 = CLBLL_R_X75Y122_SLICE_X114Y122_AQ;
  assign CLBLM_L_X70Y111_SLICE_X105Y111_B2 = CLBLM_L_X70Y111_SLICE_X105Y111_BQ;
  assign CLBLL_R_X77Y124_SLICE_X119Y124_B1 = CLBLL_R_X77Y124_SLICE_X119Y124_AQ;
  assign CLBLL_R_X77Y124_SLICE_X119Y124_B2 = CLBLL_R_X77Y123_SLICE_X118Y123_DO6;
  assign CLBLL_R_X77Y124_SLICE_X119Y124_B3 = CLBLM_L_X76Y119_SLICE_X116Y119_BO6;
  assign CLBLL_R_X77Y124_SLICE_X119Y124_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y124_SLICE_X119Y124_B5 = CLBLL_R_X75Y122_SLICE_X114Y122_AQ;
  assign CLBLL_R_X77Y124_SLICE_X119Y124_B6 = CLBLL_R_X77Y124_SLICE_X119Y124_BQ;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_A1 = CLBLM_R_X65Y99_SLICE_X99Y99_DQ;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_A3 = CLBLM_L_X64Y99_SLICE_X97Y99_AQ;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_A4 = CLBLM_L_X64Y99_SLICE_X96Y99_BQ;
  assign CLBLL_R_X77Y124_SLICE_X119Y124_C1 = CLBLL_R_X77Y123_SLICE_X118Y123_DO6;
  assign CLBLL_R_X77Y124_SLICE_X119Y124_C2 = CLBLL_R_X77Y124_SLICE_X119Y124_CQ;
  assign CLBLL_R_X77Y124_SLICE_X119Y124_C3 = CLBLL_R_X77Y124_SLICE_X119Y124_BQ;
  assign CLBLL_R_X77Y124_SLICE_X119Y124_C4 = CLBLL_R_X77Y124_SLICE_X119Y124_AQ;
  assign CLBLL_R_X77Y124_SLICE_X119Y124_C5 = CLBLL_R_X77Y124_SLICE_X119Y124_DO6;
  assign CLBLL_R_X77Y124_SLICE_X119Y124_C6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_A6 = 1'b1;
  assign CLBLL_R_X77Y124_SLICE_X119Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_B1 = CLBLM_L_X64Y99_SLICE_X97Y99_B5Q;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_B2 = CLBLM_L_X64Y99_SLICE_X97Y99_BQ;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_B3 = CLBLM_L_X64Y99_SLICE_X97Y99_AQ;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_B5 = CLBLM_R_X65Y99_SLICE_X99Y99_DQ;
  assign CLBLL_R_X77Y124_SLICE_X119Y124_D1 = CLBLL_R_X75Y122_SLICE_X114Y122_AQ;
  assign CLBLL_R_X77Y124_SLICE_X119Y124_D2 = CLBLL_R_X77Y123_SLICE_X118Y123_DO6;
  assign CLBLL_R_X77Y124_SLICE_X119Y124_D3 = CLBLM_L_X76Y119_SLICE_X116Y119_BO6;
  assign CLBLL_R_X77Y124_SLICE_X119Y124_D4 = 1'b1;
  assign CLBLL_R_X77Y124_SLICE_X119Y124_D5 = 1'b1;
  assign CLBLL_R_X77Y124_SLICE_X119Y124_D6 = 1'b1;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_C2 = 1'b1;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_C3 = 1'b1;
  assign CLBLL_R_X77Y124_SLICE_X119Y124_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_C5 = 1'b1;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_C6 = 1'b1;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X70Y111_SLICE_X104Y111_A2 = CLBLM_L_X72Y111_SLICE_X109Y111_AQ;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_D1 = 1'b1;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_D2 = 1'b1;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_D3 = 1'b1;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_D4 = 1'b1;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_D5 = 1'b1;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_D6 = 1'b1;
  assign CLBLM_L_X70Y111_SLICE_X104Y111_AX = CLBLM_L_X70Y111_SLICE_X104Y111_BO6;
  assign CLBLM_L_X70Y111_SLICE_X104Y111_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X70Y111_SLICE_X104Y111_B2 = CLBLM_L_X70Y110_SLICE_X104Y110_BQ;
  assign CLBLM_L_X70Y111_SLICE_X104Y111_B3 = CLBLM_L_X70Y111_SLICE_X104Y111_AQ;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_A6 = 1'b1;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_A1 = CLBLM_R_X63Y99_SLICE_X94Y99_A5Q;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_A2 = CLBLM_L_X64Y99_SLICE_X96Y99_A5Q;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_A3 = CLBLM_L_X64Y99_SLICE_X96Y99_AQ;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_A5 = 1'b1;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_A6 = 1'b1;
  assign CLBLM_L_X70Y111_SLICE_X104Y111_C1 = CLBLM_L_X70Y111_SLICE_X104Y111_BQ;
  assign CLBLM_L_X70Y111_SLICE_X104Y111_C2 = CLBLL_R_X71Y111_SLICE_X107Y111_AQ;
  assign CLBLM_L_X70Y111_SLICE_X104Y111_C3 = CLBLM_L_X72Y111_SLICE_X109Y111_A5Q;
  assign CLBLM_L_X70Y111_SLICE_X104Y111_C4 = CLBLM_L_X70Y112_SLICE_X104Y112_A5Q;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_B1 = CLBLM_R_X63Y99_SLICE_X94Y99_A5Q;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_B2 = CLBLM_L_X64Y99_SLICE_X96Y99_BQ;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_B3 = 1'b1;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_B5 = CLBLM_L_X64Y99_SLICE_X96Y99_A5Q;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_B6 = 1'b1;
  assign CLBLM_L_X70Y111_SLICE_X104Y111_D1 = CLBLM_L_X70Y110_SLICE_X104Y110_BQ;
  assign CLBLM_L_X70Y111_SLICE_X104Y111_D2 = CLBLL_R_X71Y111_SLICE_X107Y111_AQ;
  assign CLBLM_L_X70Y111_SLICE_X104Y111_D3 = CLBLM_L_X70Y110_SLICE_X104Y110_B5Q;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_C1 = CLBLM_L_X62Y98_SLICE_X93Y98_CQ;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_C2 = CLBLM_L_X64Y99_SLICE_X96Y99_CQ;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_C3 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_C4 = 1'b1;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_C5 = CLBLM_L_X64Y99_SLICE_X96Y99_BO5;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_C6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y111_SLICE_X104Y111_D6 = CLBLM_L_X70Y112_SLICE_X104Y112_AQ;
  assign CLBLM_L_X70Y111_SLICE_X104Y111_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X76Y119_SLICE_X116Y119_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_D1 = CLBLL_R_X77Y104_SLICE_X119Y104_A5Q;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_D1 = 1'b1;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_D2 = 1'b1;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_D3 = 1'b1;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_D4 = 1'b1;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_D5 = 1'b1;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_D6 = 1'b1;
  assign RIOB33_X105Y113_IOB_X1Y114_O = 1'b0;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign RIOB33_X105Y113_IOB_X1Y113_O = CLBLM_L_X62Y99_SLICE_X93Y99_AQ;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_T1 = 1'b1;
  assign CLBLM_L_X76Y123_SLICE_X116Y123_D3 = CLBLL_R_X75Y113_SLICE_X114Y113_AQ;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_D1 = RIOB33_X105Y59_IOB_X1Y60_I;
  assign CLBLM_L_X76Y123_SLICE_X116Y123_D4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X76Y123_SLICE_X116Y123_D5 = 1'b1;
  assign RIOI3_SING_X105Y50_ILOGIC_X1Y50_D = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_T1 = 1'b1;
  assign CLBLM_L_X76Y123_SLICE_X116Y123_D6 = CLBLM_L_X74Y123_SLICE_X113Y123_BQ;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_D1 = 1'b1;
  assign RIOB33_X105Y161_IOB_X1Y162_O = 1'b1;
  assign RIOB33_X105Y161_IOB_X1Y161_O = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_D1 = RIOB33_X105Y53_IOB_X1Y54_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1 = CLBLL_R_X71Y124_SLICE_X106Y124_AQ;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_T1 = 1'b1;
  assign CLBLM_L_X76Y123_SLICE_X116Y123_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_D1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_T1 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_A1 = CLBLL_R_X77Y125_SLICE_X118Y125_CQ;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_A2 = CLBLL_R_X77Y125_SLICE_X118Y125_BQ;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_A3 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_A5 = CLBLM_R_X67Y116_SLICE_X100Y116_AQ;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_A6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1 = CLBLM_R_X63Y122_SLICE_X95Y122_CQ;
  assign LIOB33_X0Y171_IOB_X0Y171_O = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_B1 = CLBLL_R_X77Y125_SLICE_X118Y125_CQ;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_B2 = CLBLL_R_X77Y125_SLICE_X118Y125_BQ;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_B3 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_B5 = CLBLL_R_X77Y125_SLICE_X118Y125_A5Q;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_B6 = 1'b1;
  assign LIOB33_X0Y171_IOB_X0Y172_O = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_C1 = CLBLL_R_X77Y127_SLICE_X118Y127_AQ;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_C2 = CLBLL_R_X77Y125_SLICE_X118Y125_CQ;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_C3 = CLBLL_R_X77Y125_SLICE_X118Y125_BQ;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_C4 = CLBLL_R_X77Y125_SLICE_X118Y125_A5Q;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_C5 = CLBLM_L_X76Y125_SLICE_X117Y125_CO6;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_C6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_D1 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_D2 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_D3 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_D4 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_D5 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_D6 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X70Y112_SLICE_X105Y112_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y112_SLICE_X105Y112_A2 = CLBLM_L_X70Y112_SLICE_X105Y112_BQ;
  assign CLBLM_L_X70Y112_SLICE_X105Y112_A3 = CLBLM_L_X70Y112_SLICE_X105Y112_AQ;
  assign CLBLM_L_X70Y112_SLICE_X105Y112_A4 = CLBLL_R_X71Y112_SLICE_X106Y112_BQ;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_A1 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_A2 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_A3 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_A4 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_A5 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_A6 = 1'b1;
  assign CLBLM_L_X70Y112_SLICE_X105Y112_B1 = CLBLL_R_X71Y112_SLICE_X106Y112_B5Q;
  assign CLBLM_L_X70Y112_SLICE_X105Y112_A5 = CLBLM_L_X70Y112_SLICE_X105Y112_A5Q;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_B1 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_B2 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_B3 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_B4 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_B5 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_B6 = 1'b1;
  assign CLBLM_L_X70Y112_SLICE_X105Y112_B2 = CLBLM_L_X70Y112_SLICE_X105Y112_A5Q;
  assign CLBLM_L_X70Y112_SLICE_X105Y112_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y112_SLICE_X105Y112_B5 = CLBLL_R_X71Y112_SLICE_X106Y112_BQ;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_C1 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_C2 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_C3 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_C4 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_C5 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_C6 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_A2 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_A3 = CLBLM_L_X64Y100_SLICE_X97Y100_AQ;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_A4 = CLBLM_L_X64Y99_SLICE_X96Y99_CQ;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_A5 = CLBLM_R_X63Y98_SLICE_X95Y98_AO6;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_A6 = CLBLM_L_X64Y103_SLICE_X97Y103_CO6;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_B1 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_D1 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_D2 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_D3 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_D4 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_D5 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_D6 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_B3 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_B4 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_B6 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_C1 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_C2 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_C3 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_C4 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_C5 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_C6 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X70Y112_SLICE_X104Y112_A2 = CLBLM_L_X70Y111_SLICE_X104Y111_BQ;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_D1 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_D2 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_D3 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_D4 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_D5 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_D6 = 1'b1;
  assign CLBLM_L_X70Y112_SLICE_X104Y112_AX = CLBLM_L_X70Y112_SLICE_X104Y112_BO6;
  assign CLBLM_L_X70Y112_SLICE_X104Y112_B1 = CLBLL_R_X71Y111_SLICE_X107Y111_AQ;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X70Y112_SLICE_X104Y112_B2 = CLBLM_L_X70Y111_SLICE_X104Y111_AO6;
  assign CLBLM_L_X70Y112_SLICE_X104Y112_B3 = CLBLM_L_X70Y112_SLICE_X104Y112_AQ;
  assign CLBLM_L_X70Y112_SLICE_X104Y112_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_A1 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_A2 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_A3 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_A4 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_A5 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_A6 = 1'b1;
  assign CLBLM_L_X70Y112_SLICE_X104Y112_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y112_SLICE_X104Y112_C2 = CLBLM_L_X70Y112_SLICE_X105Y112_C5Q;
  assign CLBLM_L_X70Y112_SLICE_X104Y112_C3 = CLBLM_L_X70Y112_SLICE_X104Y112_DQ;
  assign CLBLM_L_X70Y112_SLICE_X104Y112_C4 = CLBLM_L_X70Y112_SLICE_X105Y112_B5Q;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_B1 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_B2 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_B3 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_B4 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_B5 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_B6 = 1'b1;
  assign CLBLM_L_X70Y112_SLICE_X104Y112_D1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y112_SLICE_X104Y112_D2 = CLBLL_R_X71Y111_SLICE_X107Y111_AQ;
  assign CLBLM_L_X70Y112_SLICE_X104Y112_D3 = CLBLM_L_X72Y111_SLICE_X109Y111_CQ;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_C1 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_C2 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_C3 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_C4 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_C5 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_C6 = 1'b1;
  assign CLBLM_L_X70Y112_SLICE_X104Y112_D6 = CLBLM_L_X70Y110_SLICE_X104Y110_AO5;
  assign CLBLM_L_X70Y112_SLICE_X104Y112_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_D1 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_D2 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_D3 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_D4 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_D5 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_D6 = 1'b1;
  assign CLBLM_R_X67Y109_SLICE_X101Y109_D1 = CLBLM_L_X68Y108_SLICE_X102Y108_AQ;
  assign LIOB33_X0Y173_IOB_X0Y174_O = CLBLM_L_X62Y107_SLICE_X92Y107_AO5;
  assign LIOB33_X0Y173_IOB_X0Y173_O = CLBLM_L_X68Y107_SLICE_X102Y107_BO6;
  assign CLBLL_R_X77Y126_SLICE_X118Y126_A1 = CLBLL_R_X77Y123_SLICE_X119Y123_CQ;
  assign CLBLL_R_X77Y126_SLICE_X118Y126_A2 = CLBLL_R_X77Y126_SLICE_X118Y126_BQ;
  assign CLBLL_R_X77Y126_SLICE_X118Y126_A3 = CLBLL_R_X77Y126_SLICE_X118Y126_AQ;
  assign CLBLL_R_X77Y126_SLICE_X118Y126_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y126_SLICE_X118Y126_A5 = CLBLM_L_X76Y124_SLICE_X117Y124_BQ;
  assign CLBLL_R_X77Y126_SLICE_X118Y126_A6 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X118Y126_AX = CLBLM_L_X62Y105_SLICE_X93Y105_A5Q;
  assign CLBLL_R_X77Y126_SLICE_X118Y126_B1 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X118Y126_B2 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X118Y126_B3 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X118Y126_B4 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X118Y126_B5 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X118Y126_B6 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X118Y126_BX = CLBLL_R_X77Y126_SLICE_X118Y126_AO6;
  assign CLBLL_R_X77Y126_SLICE_X118Y126_C1 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X118Y126_C2 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X118Y126_C3 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X118Y126_C4 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X118Y126_C5 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X118Y126_C6 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X118Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_A1 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_A2 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_A3 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X118Y126_D1 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X118Y126_D2 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X118Y126_D3 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X118Y126_D4 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X118Y126_D5 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X118Y126_D6 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_A4 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_A5 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X118Y126_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_A6 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_A1 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_A2 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_A3 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_A4 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_A5 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_A6 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_B4 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_B5 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_B1 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_B2 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_B3 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_B4 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_B5 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_B6 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_C4 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_C5 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_C1 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_C2 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_C3 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X119Y126_A1 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X119Y126_A2 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X119Y126_A3 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X119Y126_A4 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X119Y126_A5 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X119Y126_A6 = 1'b1;
  assign CLBLM_L_X70Y113_SLICE_X105Y113_A1 = 1'b1;
  assign CLBLM_L_X70Y113_SLICE_X105Y113_A2 = 1'b1;
  assign CLBLM_L_X70Y113_SLICE_X105Y113_A3 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X119Y126_B1 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X119Y126_B2 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X119Y126_B3 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X119Y126_B4 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X119Y126_B5 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X119Y126_B6 = 1'b1;
  assign CLBLM_L_X70Y113_SLICE_X105Y113_B1 = 1'b1;
  assign CLBLM_L_X70Y113_SLICE_X105Y113_B2 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X119Y126_C1 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X119Y126_C2 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X119Y126_C3 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X119Y126_C4 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X119Y126_C5 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X119Y126_C6 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_A1 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_A2 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_A3 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_A4 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_A5 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_A6 = 1'b1;
  assign CLBLM_L_X70Y113_SLICE_X105Y113_C3 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X119Y126_D1 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X119Y126_D2 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X119Y126_D3 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X119Y126_D4 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X119Y126_D5 = 1'b1;
  assign CLBLL_R_X77Y126_SLICE_X119Y126_D6 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_B1 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_B2 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_B3 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_B4 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_B5 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_C3 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_B6 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_C1 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_C2 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_C4 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_C5 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_C6 = 1'b1;
  assign CLBLM_L_X70Y113_SLICE_X104Y113_A1 = 1'b1;
  assign CLBLM_L_X70Y113_SLICE_X104Y113_A2 = CLBLM_L_X70Y112_SLICE_X105Y112_D5Q;
  assign CLBLM_L_X70Y113_SLICE_X104Y113_A3 = CLBLM_L_X70Y113_SLICE_X104Y113_AQ;
  assign CLBLM_L_X70Y113_SLICE_X104Y113_A4 = CLBLM_L_X70Y112_SLICE_X105Y112_B5Q;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_D1 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_D2 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_D3 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_D4 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_D5 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_D6 = 1'b1;
  assign CLBLM_L_X70Y113_SLICE_X104Y113_B1 = CLBLM_L_X70Y107_SLICE_X104Y107_AQ;
  assign CLBLM_L_X70Y113_SLICE_X104Y113_B2 = CLBLM_L_X70Y113_SLICE_X104Y113_A5Q;
  assign CLBLM_L_X70Y113_SLICE_X104Y113_B3 = CLBLM_L_X70Y112_SLICE_X104Y112_C5Q;
  assign CLBLM_L_X70Y113_SLICE_X104Y113_B4 = CLBLM_L_X70Y112_SLICE_X105Y112_B5Q;
  assign CLBLM_L_X70Y113_SLICE_X104Y113_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_A1 = CLBLM_R_X63Y101_SLICE_X94Y101_BQ;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_A2 = CLBLM_L_X68Y101_SLICE_X102Y101_AQ;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_A3 = CLBLM_L_X62Y100_SLICE_X93Y100_AO6;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_A5 = CLBLM_L_X64Y101_SLICE_X96Y101_A5Q;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_A6 = 1'b1;
  assign CLBLM_L_X70Y113_SLICE_X104Y113_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y113_SLICE_X104Y113_C2 = CLBLM_R_X65Y106_SLICE_X99Y106_DQ;
  assign CLBLM_L_X70Y113_SLICE_X104Y113_C3 = CLBLM_L_X70Y113_SLICE_X104Y113_BQ;
  assign CLBLM_L_X70Y113_SLICE_X104Y113_C4 = CLBLM_L_X70Y112_SLICE_X105Y112_B5Q;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_B1 = CLBLM_L_X64Y101_SLICE_X96Y101_B5Q;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_B2 = CLBLM_L_X64Y101_SLICE_X96Y101_BQ;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_B4 = CLBLM_L_X64Y103_SLICE_X97Y103_DO6;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_B5 = CLBLM_L_X64Y101_SLICE_X96Y101_C5Q;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_B6 = 1'b1;
  assign CLBLM_L_X70Y113_SLICE_X104Y113_D1 = 1'b1;
  assign CLBLM_L_X70Y113_SLICE_X104Y113_D2 = 1'b1;
  assign CLBLM_L_X70Y113_SLICE_X104Y113_D3 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_C1 = CLBLM_L_X62Y100_SLICE_X93Y100_AO6;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_C2 = CLBLM_L_X64Y101_SLICE_X96Y101_CQ;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_C3 = CLBLM_L_X64Y101_SLICE_X96Y101_C5Q;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_C4 = CLBLM_L_X64Y101_SLICE_X96Y101_A5Q;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_C5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_C6 = 1'b1;
  assign CLBLM_L_X70Y113_SLICE_X104Y113_D6 = 1'b1;
  assign CLBLM_L_X70Y113_SLICE_X104Y113_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_D1 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_D2 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_D3 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_D4 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_D5 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_D6 = 1'b1;
  assign RIOI3_X105Y75_OLOGIC_X1Y76_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_D1 = CLBLM_R_X103Y67_SLICE_X163Y67_AQ;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_A4 = CLBLM_L_X72Y121_SLICE_X108Y121_BO6;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_A5 = CLBLL_R_X71Y121_SLICE_X106Y121_AQ;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_A6 = CLBLM_L_X72Y122_SLICE_X108Y122_AQ;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_T1 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_T1 = 1'b1;
  assign RIOI3_X105Y75_OLOGIC_X1Y75_D1 = CLBLM_R_X103Y75_SLICE_X162Y75_CQ;
  assign RIOI3_SING_X105Y100_OLOGIC_X1Y100_D1 = CLBLM_L_X78Y104_SLICE_X120Y104_A5Q;
  assign LIOB33_X0Y175_IOB_X0Y176_O = CLBLM_L_X70Y135_SLICE_X104Y135_CO6;
  assign LIOB33_X0Y175_IOB_X0Y175_O = CLBLM_R_X63Y105_SLICE_X95Y105_A5Q;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_B2 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_B3 = 1'b1;
  assign RIOI3_SING_X105Y100_OLOGIC_X1Y100_T1 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_B4 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_B5 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_B6 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_D1 = CLBLM_R_X103Y67_SLICE_X162Y67_AQ;
  assign RIOI3_X105Y75_OLOGIC_X1Y75_T1 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X118Y127_A1 = CLBLL_R_X77Y125_SLICE_X118Y125_BO5;
  assign CLBLL_R_X77Y127_SLICE_X118Y127_A2 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X118Y127_A3 = CLBLL_R_X77Y127_SLICE_X118Y127_AQ;
  assign CLBLL_R_X77Y127_SLICE_X118Y127_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y127_SLICE_X118Y127_A5 = CLBLL_R_X79Y127_SLICE_X122Y127_BQ;
  assign CLBLL_R_X77Y127_SLICE_X118Y127_A6 = CLBLL_R_X79Y127_SLICE_X122Y127_A5Q;
  assign CLBLM_L_X68Y112_SLICE_X103Y112_C6 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X118Y127_B1 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X118Y127_B2 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X118Y127_B3 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X118Y127_B4 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X118Y127_B5 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X118Y127_B6 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X118Y127_C1 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X118Y127_C2 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X118Y127_C3 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X118Y127_C4 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X118Y127_C5 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X118Y127_C6 = 1'b1;
  assign CLBLM_R_X67Y118_SLICE_X100Y118_D5 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X118Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_C5 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X118Y127_D1 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X118Y127_D2 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X118Y127_D3 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X118Y127_D4 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X118Y127_D5 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X118Y127_D6 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_C6 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_CE = CLBLM_L_X76Y109_SLICE_X116Y109_AO6;
  assign CLBLL_R_X77Y127_SLICE_X118Y127_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X76Y134_SLICE_X117Y134_A1 = CLBLM_L_X76Y134_SLICE_X116Y134_CO6;
  assign CLBLM_L_X76Y134_SLICE_X117Y134_A2 = 1'b1;
  assign CLBLM_L_X76Y134_SLICE_X117Y134_A3 = CLBLM_L_X76Y134_SLICE_X117Y134_AQ;
  assign CLBLM_L_X76Y134_SLICE_X117Y134_A4 = CLBLM_L_X76Y134_SLICE_X116Y134_BQ;
  assign CLBLM_L_X76Y134_SLICE_X117Y134_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X76Y134_SLICE_X117Y134_A6 = CLBLM_L_X76Y134_SLICE_X117Y134_CO6;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_A2 = CLBLL_R_X75Y128_SLICE_X115Y128_AO6;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_A3 = CLBLM_L_X74Y126_SLICE_X113Y126_AQ;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_A4 = CLBLM_L_X74Y126_SLICE_X112Y126_A5Q;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_A5 = CLBLM_L_X74Y126_SLICE_X113Y126_A5Q;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_A6 = 1'b1;
  assign CLBLM_L_X76Y134_SLICE_X117Y134_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_B2 = CLBLM_L_X74Y126_SLICE_X113Y126_BQ;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_B3 = CLBLM_L_X74Y126_SLICE_X113Y126_AQ;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_B4 = CLBLL_R_X75Y128_SLICE_X115Y128_AO6;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_B5 = CLBLM_L_X74Y128_SLICE_X113Y128_AO6;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_B6 = CLBLM_L_X74Y126_SLICE_X113Y126_A5Q;
  assign CLBLM_L_X76Y134_SLICE_X117Y134_C4 = CLBLM_L_X76Y133_SLICE_X116Y133_BQ;
  assign CLBLM_L_X76Y134_SLICE_X117Y134_C5 = CLBLM_L_X76Y134_SLICE_X116Y134_AQ;
  assign CLBLL_R_X77Y127_SLICE_X119Y127_A1 = CLBLM_L_X78Y127_SLICE_X121Y127_CO6;
  assign CLBLL_R_X77Y127_SLICE_X119Y127_A2 = CLBLL_R_X77Y123_SLICE_X119Y123_DO6;
  assign CLBLL_R_X77Y127_SLICE_X119Y127_A3 = CLBLL_R_X77Y127_SLICE_X119Y127_AQ;
  assign CLBLL_R_X77Y127_SLICE_X119Y127_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y127_SLICE_X119Y127_A5 = CLBLM_L_X78Y127_SLICE_X121Y127_BO6;
  assign CLBLL_R_X77Y127_SLICE_X119Y127_A6 = 1'b1;
  assign CLBLM_L_X70Y114_SLICE_X105Y114_A1 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X103Y112_D6 = 1'b1;
  assign CLBLM_L_X70Y114_SLICE_X105Y114_A2 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X119Y127_B1 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X119Y127_B2 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X119Y127_B3 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X119Y127_B4 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X119Y127_B5 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X119Y127_B6 = 1'b1;
  assign CLBLM_L_X70Y114_SLICE_X105Y114_A3 = 1'b1;
  assign CLBLM_L_X70Y114_SLICE_X105Y114_A4 = 1'b1;
  assign CLBLM_L_X70Y114_SLICE_X105Y114_A5 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X119Y127_C1 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X119Y127_C2 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X119Y127_C3 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X119Y127_C4 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X119Y127_C5 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X119Y127_C6 = 1'b1;
  assign CLBLM_L_X70Y114_SLICE_X105Y114_B2 = 1'b1;
  assign CLBLM_L_X70Y114_SLICE_X105Y114_B3 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X119Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X70Y114_SLICE_X105Y114_B5 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_A1 = CLBLM_R_X65Y104_SLICE_X99Y104_DO6;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_A2 = CLBLM_R_X65Y104_SLICE_X98Y104_CQ;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_A3 = CLBLM_R_X63Y99_SLICE_X95Y99_CO6;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y127_SLICE_X119Y127_D1 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X119Y127_D2 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X119Y127_D3 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X119Y127_D4 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X119Y127_D5 = 1'b1;
  assign CLBLL_R_X77Y127_SLICE_X119Y127_D6 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_A5 = CLBLM_R_X65Y104_SLICE_X98Y104_C5Q;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_A6 = CLBLM_L_X64Y103_SLICE_X97Y103_CO6;
  assign CLBLL_R_X77Y127_SLICE_X119Y127_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_B2 = CLBLM_R_X65Y104_SLICE_X98Y104_CQ;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_B3 = CLBLM_R_X65Y104_SLICE_X98Y104_C5Q;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_B4 = CLBLM_L_X64Y103_SLICE_X97Y103_DO6;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_C1 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_C2 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_C3 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_C4 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_C5 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_C6 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X70Y114_SLICE_X104Y114_A1 = CLBLL_R_X71Y117_SLICE_X106Y117_B5Q;
  assign CLBLM_L_X70Y114_SLICE_X104Y114_A2 = 1'b1;
  assign CLBLM_L_X70Y114_SLICE_X104Y114_A3 = CLBLM_L_X70Y114_SLICE_X104Y114_AQ;
  assign CLBLM_L_X70Y114_SLICE_X104Y114_A4 = CLBLM_L_X68Y109_SLICE_X102Y109_AQ;
  assign CLBLM_L_X70Y114_SLICE_X104Y114_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_D1 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_D2 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_D3 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_D4 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_D5 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_D6 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X102Y112_A5 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X102Y112_A6 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X70Y114_SLICE_X104Y114_B3 = 1'b1;
  assign CLBLM_L_X70Y114_SLICE_X104Y114_C2 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_A1 = CLBLM_R_X63Y102_SLICE_X95Y102_AQ;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_A2 = CLBLM_L_X64Y102_SLICE_X96Y102_A5Q;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_A3 = CLBLM_L_X64Y102_SLICE_X96Y102_AQ;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_A5 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_A6 = 1'b1;
  assign CLBLM_L_X70Y114_SLICE_X104Y114_C1 = 1'b1;
  assign CLBLM_L_X70Y114_SLICE_X104Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X70Y114_SLICE_X104Y114_C3 = 1'b1;
  assign CLBLM_L_X70Y114_SLICE_X104Y114_C4 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_B1 = CLBLM_L_X64Y105_SLICE_X96Y105_CQ;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_B2 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_B3 = CLBLM_L_X64Y105_SLICE_X96Y105_C5Q;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_B4 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_B5 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_B6 = 1'b1;
  assign CLBLM_L_X70Y114_SLICE_X104Y114_D1 = 1'b1;
  assign CLBLM_L_X70Y114_SLICE_X104Y114_D6 = 1'b1;
  assign CLBLM_L_X70Y114_SLICE_X104Y114_D2 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_C1 = CLBLM_R_X63Y102_SLICE_X94Y102_DO5;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_C2 = CLBLM_L_X64Y102_SLICE_X96Y102_CQ;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_C3 = CLBLM_R_X63Y102_SLICE_X94Y102_BQ;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_C4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_C5 = CLBLM_L_X64Y102_SLICE_X96Y102_BO5;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_C6 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X68Y112_SLICE_X102Y112_B1 = 1'b1;
  assign CLBLM_L_X70Y114_SLICE_X104Y114_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X68Y112_SLICE_X102Y112_B3 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_D1 = CLBLM_L_X64Y101_SLICE_X96Y101_BQ;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_D2 = CLBLM_L_X64Y101_SLICE_X96Y101_CQ;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_D3 = CLBLM_L_X64Y101_SLICE_X96Y101_C5Q;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_D4 = CLBLM_L_X64Y101_SLICE_X96Y101_B5Q;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_D5 = CLBLM_L_X64Y102_SLICE_X97Y102_BQ;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_D6 = CLBLM_L_X64Y103_SLICE_X97Y103_DO6;
  assign CLBLM_L_X68Y112_SLICE_X102Y112_B4 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_D1 = CLBLL_R_X75Y133_SLICE_X114Y133_AQ;
  assign LIOB33_X0Y177_IOB_X0Y178_O = CLBLM_L_X72Y122_SLICE_X108Y122_AO6;
  assign LIOB33_X0Y177_IOB_X0Y177_O = CLBLM_L_X70Y134_SLICE_X104Y134_CO5;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_D4 = 1'b1;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_D5 = 1'b1;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_D6 = 1'b1;
  assign CLBLL_R_X77Y128_SLICE_X118Y128_A1 = CLBLL_R_X77Y128_SLICE_X119Y128_BQ;
  assign CLBLL_R_X77Y128_SLICE_X118Y128_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y128_SLICE_X118Y128_A3 = CLBLL_R_X77Y129_SLICE_X118Y129_CQ;
  assign CLBLL_R_X77Y128_SLICE_X118Y128_A4 = CLBLL_R_X77Y129_SLICE_X119Y129_AO6;
  assign CLBLL_R_X77Y128_SLICE_X118Y128_A5 = CLBLL_R_X77Y128_SLICE_X118Y128_CQ;
  assign CLBLL_R_X77Y128_SLICE_X118Y128_A6 = 1'b1;
  assign RIOI3_SING_X105Y149_OLOGIC_X1Y149_D1 = CLBLM_L_X76Y111_SLICE_X116Y111_BQ;
  assign CLBLL_R_X77Y128_SLICE_X118Y128_AX = CLBLM_L_X76Y127_SLICE_X116Y127_AQ;
  assign CLBLM_L_X68Y112_SLICE_X102Y112_D3 = 1'b1;
  assign CLBLL_R_X77Y128_SLICE_X118Y128_B1 = CLBLM_L_X76Y128_SLICE_X116Y128_A5Q;
  assign CLBLL_R_X77Y128_SLICE_X118Y128_B2 = CLBLM_L_X76Y128_SLICE_X116Y128_CQ;
  assign CLBLL_R_X77Y128_SLICE_X118Y128_B3 = CLBLL_R_X77Y128_SLICE_X119Y128_A5Q;
  assign CLBLL_R_X77Y128_SLICE_X118Y128_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y128_SLICE_X118Y128_B5 = 1'b1;
  assign CLBLL_R_X77Y128_SLICE_X118Y128_B6 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X102Y112_D4 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X102Y112_D5 = 1'b1;
  assign CLBLL_R_X77Y128_SLICE_X118Y128_C1 = CLBLL_R_X77Y129_SLICE_X118Y129_AQ;
  assign CLBLL_R_X77Y128_SLICE_X118Y128_C2 = CLBLL_R_X77Y128_SLICE_X119Y128_BQ;
  assign CLBLL_R_X77Y128_SLICE_X118Y128_C3 = CLBLM_L_X76Y128_SLICE_X116Y128_CQ;
  assign CLBLL_R_X77Y128_SLICE_X118Y128_C4 = CLBLL_R_X77Y130_SLICE_X119Y130_AQ;
  assign CLBLL_R_X77Y128_SLICE_X118Y128_C5 = 1'b1;
  assign CLBLL_R_X77Y128_SLICE_X118Y128_C6 = 1'b1;
  assign RIOI3_SING_X105Y149_OLOGIC_X1Y149_T1 = 1'b1;
  assign CLBLL_R_X77Y128_SLICE_X118Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X77Y128_SLICE_X118Y128_CX = CLBLL_R_X77Y128_SLICE_X118Y128_AO5;
  assign CLBLL_R_X77Y128_SLICE_X118Y128_D1 = 1'b1;
  assign CLBLL_R_X77Y128_SLICE_X118Y128_D2 = 1'b1;
  assign CLBLL_R_X77Y128_SLICE_X118Y128_D3 = 1'b1;
  assign CLBLL_R_X77Y128_SLICE_X118Y128_D4 = 1'b1;
  assign CLBLL_R_X77Y128_SLICE_X118Y128_D5 = 1'b1;
  assign CLBLL_R_X77Y128_SLICE_X118Y128_D6 = 1'b1;
  assign CLBLL_R_X77Y128_SLICE_X118Y128_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X76Y134_SLICE_X116Y134_A1 = CLBLM_L_X76Y134_SLICE_X116Y134_AQ;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_A1 = CLBLM_L_X74Y127_SLICE_X113Y127_AQ;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_A2 = CLBLM_L_X74Y128_SLICE_X112Y128_AQ;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_A3 = CLBLL_R_X75Y128_SLICE_X114Y128_DO6;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_A4 = CLBLM_L_X74Y127_SLICE_X113Y127_BO6;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_A6 = CLBLM_L_X74Y127_SLICE_X113Y127_A5Q;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_AX = CLBLM_L_X74Y127_SLICE_X112Y127_AO5;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_B1 = CLBLL_R_X75Y128_SLICE_X115Y128_DO6;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_B2 = CLBLM_L_X74Y127_SLICE_X113Y127_A5Q;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_B3 = 1'b1;
  assign CLBLL_R_X77Y128_SLICE_X119Y128_A1 = CLBLL_R_X77Y128_SLICE_X119Y128_AQ;
  assign CLBLL_R_X77Y128_SLICE_X119Y128_A2 = CLBLM_L_X78Y128_SLICE_X120Y128_AQ;
  assign CLBLL_R_X77Y128_SLICE_X119Y128_A3 = CLBLL_R_X77Y128_SLICE_X118Y128_AO6;
  assign CLBLL_R_X77Y128_SLICE_X119Y128_A4 = CLBLL_R_X77Y128_SLICE_X118Y128_BQ;
  assign CLBLL_R_X77Y128_SLICE_X119Y128_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y128_SLICE_X119Y128_A6 = CLBLL_R_X77Y128_SLICE_X118Y128_CQ;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_B4 = CLBLM_L_X74Y129_SLICE_X112Y129_A5Q;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_B5 = 1'b1;
  assign CLBLL_R_X77Y128_SLICE_X119Y128_AX = CLBLL_R_X77Y128_SLICE_X119Y128_DQ;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_B6 = 1'b1;
  assign CLBLL_R_X77Y128_SLICE_X119Y128_B1 = CLBLM_L_X76Y127_SLICE_X116Y127_AQ;
  assign CLBLL_R_X77Y128_SLICE_X119Y128_B2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y128_SLICE_X119Y128_B3 = CLBLL_R_X77Y128_SLICE_X118Y128_CO5;
  assign CLBLL_R_X77Y128_SLICE_X119Y128_B4 = CLBLL_R_X77Y128_SLICE_X118Y128_BQ;
  assign CLBLL_R_X77Y128_SLICE_X119Y128_B5 = CLBLM_L_X78Y129_SLICE_X120Y129_AO6;
  assign CLBLL_R_X77Y128_SLICE_X119Y128_B6 = CLBLM_L_X80Y132_SLICE_X124Y132_AQ;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_C2 = CLBLM_L_X74Y127_SLICE_X113Y127_CQ;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_C4 = CLBLM_L_X74Y127_SLICE_X113Y127_AQ;
  assign CLBLL_R_X77Y128_SLICE_X119Y128_C1 = CLBLM_L_X78Y128_SLICE_X120Y128_AQ;
  assign CLBLL_R_X77Y128_SLICE_X119Y128_C2 = CLBLL_R_X77Y128_SLICE_X119Y128_CQ;
  assign CLBLL_R_X77Y128_SLICE_X119Y128_C3 = CLBLL_R_X77Y128_SLICE_X119Y128_BQ;
  assign CLBLL_R_X77Y128_SLICE_X119Y128_C4 = 1'b1;
  assign CLBLL_R_X77Y128_SLICE_X119Y128_C5 = CLBLL_R_X77Y128_SLICE_X119Y128_AQ;
  assign CLBLL_R_X77Y128_SLICE_X119Y128_C6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_B6 = 1'b1;
  assign CLBLL_R_X77Y128_SLICE_X119Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_D1 = 1'b1;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_D2 = 1'b1;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_D3 = 1'b1;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_D4 = 1'b1;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_D5 = 1'b1;
  assign CLBLL_R_X77Y128_SLICE_X119Y128_D1 = CLBLL_R_X77Y128_SLICE_X119Y128_DQ;
  assign CLBLL_R_X77Y128_SLICE_X119Y128_D2 = CLBLM_L_X62Y105_SLICE_X93Y105_A5Q;
  assign CLBLL_R_X77Y128_SLICE_X119Y128_D3 = CLBLL_R_X77Y128_SLICE_X118Y128_B5Q;
  assign CLBLL_R_X77Y128_SLICE_X119Y128_D4 = CLBLM_L_X76Y128_SLICE_X116Y128_CQ;
  assign CLBLL_R_X77Y128_SLICE_X119Y128_D5 = 1'b1;
  assign CLBLL_R_X77Y128_SLICE_X119Y128_D6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_A1 = CLBLM_L_X64Y103_SLICE_X97Y103_AQ;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_A3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y128_SLICE_X119Y128_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_B1 = CLBLM_R_X65Y104_SLICE_X99Y104_DO6;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_B2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_B3 = CLBLM_L_X64Y102_SLICE_X97Y102_BQ;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_A5 = CLBLM_L_X64Y102_SLICE_X97Y102_AQ;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_A6 = CLBLM_R_X65Y104_SLICE_X98Y104_C5Q;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_B4 = CLBLM_R_X65Y104_SLICE_X98Y104_CQ;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_B5 = CLBLM_R_X65Y104_SLICE_X98Y104_C5Q;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_B6 = CLBLM_L_X64Y103_SLICE_X97Y103_BQ;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_C1 = CLBLM_R_X65Y104_SLICE_X98Y104_C5Q;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_C2 = CLBLM_R_X65Y103_SLICE_X99Y103_CO6;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_C3 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_C4 = CLBLM_L_X64Y103_SLICE_X97Y103_AQ;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_C5 = CLBLM_R_X65Y104_SLICE_X99Y104_B5Q;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_C6 = CLBLM_R_X65Y104_SLICE_X98Y104_CQ;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_BX = CLBLM_L_X74Y129_SLICE_X112Y129_AQ;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_C1 = CLBLM_L_X72Y127_SLICE_X108Y127_AQ;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_C2 = CLBLM_L_X74Y127_SLICE_X113Y127_AQ;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_C3 = CLBLM_L_X74Y128_SLICE_X112Y128_DQ;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_C4 = CLBLM_L_X72Y127_SLICE_X108Y127_A5Q;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_C5 = 1'b1;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_C6 = CLBLM_L_X72Y128_SLICE_X108Y128_A5Q;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_D1 = CLBLM_R_X65Y104_SLICE_X98Y104_CQ;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_D2 = CLBLM_R_X65Y104_SLICE_X98Y104_C5Q;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_D3 = CLBLM_L_X64Y103_SLICE_X97Y103_BQ;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_C2 = CLBLM_L_X62Y102_SLICE_X92Y102_CQ;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_D4 = CLBLM_R_X65Y103_SLICE_X98Y103_A5Q;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_D5 = 1'b1;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_C3 = CLBLM_R_X63Y103_SLICE_X94Y103_AO5;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_D6 = CLBLM_R_X65Y103_SLICE_X99Y103_CO6;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_C5 = 1'b1;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_C6 = 1'b1;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_D1 = CLBLM_L_X72Y127_SLICE_X108Y127_AQ;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_A1 = CLBLM_R_X63Y102_SLICE_X95Y102_DQ;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_A2 = CLBLM_L_X64Y103_SLICE_X97Y103_DO6;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_A3 = CLBLM_L_X64Y103_SLICE_X96Y103_AQ;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_C5 = CLBLM_R_X63Y102_SLICE_X94Y102_DO6;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_A5 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_A6 = CLBLM_R_X63Y101_SLICE_X94Y101_DO6;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_CE = CLBLM_L_X76Y109_SLICE_X116Y109_AO6;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_B1 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_B2 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_B3 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_B4 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_B5 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_B6 = 1'b1;
  assign CLBLM_L_X76Y134_SLICE_X116Y134_A2 = CLBLL_R_X75Y133_SLICE_X115Y133_BQ;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_C1 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_C2 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_C3 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_C4 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_C5 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_C6 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_D1 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_D2 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_D3 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_D4 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_D5 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_D6 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign LIOB33_X0Y179_IOB_X0Y180_O = 1'b1;
  assign LIOB33_X0Y179_IOB_X0Y179_O = 1'b1;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_D4 = 1'b1;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_A4 = CLBLM_R_X63Y97_SLICE_X94Y97_CQ;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_D5 = 1'b1;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_A5 = CLBLM_L_X64Y97_SLICE_X97Y97_A5Q;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_A4 = CLBLL_R_X77Y113_SLICE_X118Y113_AQ;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_A5 = CLBLM_L_X78Y122_SLICE_X121Y122_AQ;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_A6 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0 = RIOB33_X105Y77_IOB_X1Y78_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_B1 = CLBLM_L_X64Y99_SLICE_X96Y99_A5Q;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_B2 = CLBLM_L_X64Y99_SLICE_X96Y99_BQ;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign RIOB33_X105Y67_IOB_X1Y68_O = CLBLM_R_X103Y67_SLICE_X163Y67_CQ;
  assign RIOB33_X105Y67_IOB_X1Y67_O = CLBLM_R_X103Y67_SLICE_X163Y67_BQ;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_B5 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_B2 = CLBLM_L_X78Y121_SLICE_X120Y121_BQ;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_B3 = CLBLM_L_X78Y120_SLICE_X120Y120_AQ;
  assign CLBLM_L_X76Y134_SLICE_X116Y134_A3 = CLBLM_L_X76Y134_SLICE_X117Y134_CO6;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_B4 = CLBLM_L_X78Y122_SLICE_X121Y122_BQ;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_B5 = CLBLM_L_X78Y122_SLICE_X121Y122_AQ;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_B6 = CLBLM_L_X78Y123_SLICE_X120Y123_CO6;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_A1 = CLBLL_R_X77Y130_SLICE_X118Y130_AO5;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_A2 = CLBLL_R_X77Y128_SLICE_X119Y128_A5Q;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_A3 = CLBLL_R_X77Y128_SLICE_X118Y128_AQ;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_A4 = CLBLL_R_X77Y128_SLICE_X118Y128_BQ;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_A6 = CLBLL_R_X77Y130_SLICE_X119Y130_AQ;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_B1 = CLBLL_R_X77Y129_SLICE_X119Y129_AO6;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_B2 = CLBLL_R_X77Y129_SLICE_X118Y129_BQ;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_B3 = CLBLL_R_X77Y129_SLICE_X118Y129_DQ;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_B4 = 1'b1;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_B6 = CLBLL_R_X77Y129_SLICE_X119Y129_DO6;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_C3 = CLBLM_L_X64Y97_SLICE_X97Y97_DQ;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_C4 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_C1 = CLBLL_R_X77Y128_SLICE_X119Y128_BQ;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_C2 = CLBLL_R_X77Y129_SLICE_X118Y129_CQ;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_C3 = CLBLL_R_X77Y128_SLICE_X118Y128_CQ;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_C4 = CLBLL_R_X77Y130_SLICE_X119Y130_CO6;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_C5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_C6 = CLBLL_R_X77Y129_SLICE_X119Y129_BQ;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_D1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_D2 = CLBLL_R_X77Y129_SLICE_X119Y129_AO6;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_D3 = CLBLL_R_X77Y129_SLICE_X118Y129_DQ;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_D4 = CLBLL_R_X77Y129_SLICE_X119Y129_DO6;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_D5 = 1'b1;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_D6 = CLBLL_R_X77Y129_SLICE_X119Y129_BQ;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_D6 = CLBLL_R_X75Y124_SLICE_X115Y124_AQ;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_D1 = CLBLM_L_X80Y132_SLICE_X124Y132_AQ;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1 = 1'b1;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_A1 = CLBLL_R_X77Y128_SLICE_X118Y128_B5Q;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_A2 = CLBLM_L_X74Y129_SLICE_X113Y129_CO6;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_A3 = CLBLL_R_X75Y130_SLICE_X115Y130_AQ;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_A4 = 1'b1;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_A5 = CLBLL_R_X75Y129_SLICE_X114Y129_DQ;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_A6 = 1'b1;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_A1 = CLBLL_R_X77Y130_SLICE_X119Y130_CO6;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_A2 = CLBLL_R_X77Y129_SLICE_X119Y129_BQ;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_A3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_A4 = CLBLL_R_X77Y128_SLICE_X118Y128_CQ;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_A5 = CLBLL_R_X77Y129_SLICE_X118Y129_CQ;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_A6 = 1'b1;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_B1 = CLBLL_R_X75Y128_SLICE_X115Y128_DO6;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_B2 = 1'b1;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_B1 = CLBLL_R_X77Y130_SLICE_X119Y130_CO6;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_B2 = CLBLL_R_X77Y129_SLICE_X119Y129_BQ;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_B4 = CLBLL_R_X77Y129_SLICE_X118Y129_BQ;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_B5 = CLBLL_R_X77Y129_SLICE_X119Y129_CO6;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_B6 = CLBLL_R_X77Y128_SLICE_X119Y128_CQ;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_B6 = 1'b1;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_C1 = CLBLM_L_X74Y129_SLICE_X112Y129_AQ;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_C1 = CLBLM_L_X78Y128_SLICE_X120Y128_AQ;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_C2 = CLBLL_R_X77Y128_SLICE_X119Y128_CQ;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_C3 = CLBLL_R_X77Y128_SLICE_X119Y128_BQ;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_C4 = CLBLL_R_X77Y129_SLICE_X119Y129_AO5;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_C5 = CLBLL_R_X77Y129_SLICE_X118Y129_DQ;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_C6 = CLBLL_R_X77Y128_SLICE_X118Y128_BQ;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_C6 = CLBLM_L_X74Y129_SLICE_X112Y129_A5Q;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_D1 = 1'b1;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_D2 = 1'b1;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_D3 = 1'b1;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_D4 = 1'b1;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_D1 = CLBLL_R_X77Y128_SLICE_X119Y128_BQ;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_D2 = CLBLL_R_X77Y128_SLICE_X119Y128_CQ;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_D3 = CLBLL_R_X77Y128_SLICE_X118Y128_BQ;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_D4 = CLBLL_R_X77Y129_SLICE_X118Y129_CQ;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_D5 = CLBLL_R_X77Y128_SLICE_X118Y128_CQ;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_D6 = CLBLM_L_X78Y128_SLICE_X120Y128_AQ;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_A3 = CLBLM_L_X64Y104_SLICE_X97Y104_AQ;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_A4 = CLBLM_L_X64Y105_SLICE_X96Y105_CQ;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_A5 = CLBLM_L_X64Y105_SLICE_X96Y105_C5Q;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_A6 = CLBLM_L_X64Y102_SLICE_X96Y102_A5Q;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_A2 = CLBLM_R_X65Y105_SLICE_X99Y105_C5Q;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_B1 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_B2 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_B3 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_B4 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_B5 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_B6 = 1'b1;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_B1 = CLBLL_R_X75Y128_SLICE_X114Y128_DO6;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_B2 = CLBLM_L_X74Y128_SLICE_X112Y128_BQ;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_C1 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_C2 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_C3 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_C4 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X91Y92_A1 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X91Y92_A2 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X91Y92_A3 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X91Y92_A4 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X91Y92_A5 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X91Y92_A6 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_C5 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_C6 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X60Y92_SLICE_X91Y92_B1 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X91Y92_B2 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X91Y92_B3 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X91Y92_B4 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X91Y92_B5 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X91Y92_B6 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_D1 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_D2 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X91Y92_C1 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X91Y92_C2 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X91Y92_C3 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X91Y92_C4 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X91Y92_C5 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X91Y92_C6 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_A1 = CLBLM_R_X63Y101_SLICE_X94Y101_BO5;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_A2 = CLBLM_L_X64Y104_SLICE_X96Y104_BQ;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_A3 = CLBLM_L_X64Y104_SLICE_X96Y104_AQ;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_A4 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_A6 = CLBLM_R_X63Y101_SLICE_X94Y101_DO6;
  assign CLBLM_L_X60Y92_SLICE_X91Y92_D1 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X91Y92_D2 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X91Y92_D3 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X91Y92_D4 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X91Y92_D5 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X91Y92_D6 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_B1 = CLBLM_L_X64Y105_SLICE_X96Y105_CQ;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_B2 = CLBLM_L_X64Y104_SLICE_X96Y104_BQ;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_B3 = CLBLM_L_X64Y105_SLICE_X96Y105_C5Q;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_C2 = CLBLM_L_X64Y104_SLICE_X96Y104_CQ;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_C3 = CLBLM_R_X63Y101_SLICE_X94Y101_BO5;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_C4 = CLBLM_L_X64Y104_SLICE_X96Y104_BQ;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_C5 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_C6 = CLBLM_L_X64Y104_SLICE_X96Y104_AQ;
  assign CLBLM_L_X60Y92_SLICE_X90Y92_A1 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X90Y92_A2 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X90Y92_A3 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X90Y92_A4 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X90Y92_A5 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X90Y92_A6 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X90Y92_AX = CLBLL_R_X71Y134_SLICE_X106Y134_AQ;
  assign CLBLM_L_X60Y92_SLICE_X90Y92_B1 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X90Y92_B2 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_D1 = CLBLM_L_X64Y105_SLICE_X96Y105_C5Q;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_D2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_D3 = CLBLM_L_X64Y104_SLICE_X96Y104_DQ;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_D4 = CLBLL_R_X79Y99_SLICE_X122Y99_AO6;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_D5 = CLBLM_L_X64Y105_SLICE_X96Y105_CQ;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_D6 = CLBLM_L_X64Y102_SLICE_X96Y102_A5Q;
  assign CLBLM_L_X60Y92_SLICE_X90Y92_B3 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X90Y92_B4 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X90Y92_B5 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X90Y92_B6 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X90Y92_BX = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_L_X60Y92_SLICE_X90Y92_C1 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X90Y92_C2 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X90Y92_C3 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X90Y92_C4 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X90Y92_C5 = 1'b1;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_A3 = CLBLM_L_X70Y129_SLICE_X104Y129_AQ;
  assign CLBLM_L_X60Y92_SLICE_X90Y92_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X60Y92_SLICE_X90Y92_C6 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_A5 = CLBLM_L_X70Y129_SLICE_X105Y129_AQ;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_C3 = CLBLM_L_X76Y124_SLICE_X117Y124_DO6;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_C5 = CLBLM_L_X76Y122_SLICE_X116Y122_BQ;
  assign CLBLM_L_X60Y92_SLICE_X90Y92_D1 = 1'b1;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_A6 = CLBLM_L_X70Y128_SLICE_X105Y128_CO6;
  assign CLBLM_L_X60Y92_SLICE_X90Y92_D2 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X90Y92_D4 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X90Y92_D5 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X90Y92_D3 = 1'b1;
  assign CLBLM_L_X60Y92_SLICE_X90Y92_D6 = 1'b1;
  assign CLBLM_L_X74Y133_SLICE_X112Y133_B6 = CLBLM_L_X74Y133_SLICE_X113Y133_AO5;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_C6 = CLBLM_L_X76Y124_SLICE_X116Y124_BO6;
  assign CLBLM_L_X60Y92_SLICE_X90Y92_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_CE = CLBLM_L_X76Y123_SLICE_X116Y123_DO6;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_D1 = CLBLL_R_X73Y123_SLICE_X110Y123_AQ;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_D1 = 1'b1;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_AX = CLBLM_L_X70Y128_SLICE_X104Y128_AQ;
  assign RIOI3_X105Y101_OLOGIC_X1Y101_D1 = CLBLM_L_X72Y109_SLICE_X109Y109_DQ;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_T1 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_T1 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_D1 = CLBLM_R_X63Y106_SLICE_X95Y106_AQ;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_T1 = 1'b1;
  assign CLBLM_R_X103Y75_SLICE_X163Y75_B3 = 1'b1;
  assign RIOI3_X105Y101_OLOGIC_X1Y101_T1 = 1'b1;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_D5 = 1'b1;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_D6 = 1'b1;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_A1 = CLBLL_R_X77Y130_SLICE_X118Y130_DO6;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_A2 = CLBLM_L_X78Y131_SLICE_X120Y131_AQ;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_A3 = CLBLL_R_X77Y130_SLICE_X118Y130_AQ;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_A4 = CLBLL_R_X77Y131_SLICE_X118Y131_AO6;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_A6 = 1'b1;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_C4 = CLBLM_L_X70Y129_SLICE_X105Y129_BQ;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_C5 = CLBLM_L_X70Y128_SLICE_X104Y128_AQ;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_B1 = CLBLL_R_X77Y130_SLICE_X118Y130_DO6;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_B2 = CLBLL_R_X77Y130_SLICE_X118Y130_BQ;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_B3 = CLBLL_R_X77Y130_SLICE_X118Y130_AQ;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_B4 = CLBLL_R_X77Y130_SLICE_X118Y130_CQ;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_B6 = 1'b1;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_C6 = CLBLM_L_X70Y128_SLICE_X104Y128_BQ;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_CE = CLBLM_L_X76Y109_SLICE_X116Y109_AO6;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_DX = CLBLL_R_X75Y124_SLICE_X115Y124_CQ;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_C2 = CLBLL_R_X77Y130_SLICE_X118Y130_CQ;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_C3 = CLBLL_R_X77Y131_SLICE_X119Y131_BQ;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_C4 = 1'b1;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_C5 = CLBLL_R_X77Y130_SLICE_X118Y130_DO6;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_C6 = CLBLL_R_X77Y130_SLICE_X118Y130_AQ;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_D1 = CLBLL_R_X77Y128_SLICE_X118Y128_BQ;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_D2 = CLBLL_R_X77Y130_SLICE_X119Y130_AQ;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_D3 = CLBLM_L_X78Y131_SLICE_X120Y131_AQ;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_D4 = CLBLL_R_X77Y130_SLICE_X118Y130_AQ;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_D5 = CLBLL_R_X77Y128_SLICE_X118Y128_AQ;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_D6 = 1'b1;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_A2 = CLBLL_R_X75Y128_SLICE_X115Y128_DO6;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_A3 = CLBLM_L_X74Y129_SLICE_X112Y129_A5Q;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_A1 = CLBLL_R_X77Y131_SLICE_X119Y131_BQ;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_A2 = CLBLL_R_X77Y130_SLICE_X119Y130_BQ;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_A3 = CLBLL_R_X77Y128_SLICE_X118Y128_BQ;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_A4 = CLBLM_L_X78Y130_SLICE_X120Y130_AQ;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_A5 = CLBLL_R_X77Y128_SLICE_X118Y128_AQ;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_A6 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_A4 = CLBLL_R_X75Y128_SLICE_X114Y128_DO5;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_A5 = CLBLM_L_X74Y129_SLICE_X112Y129_AQ;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_AX = CLBLM_L_X80Y132_SLICE_X124Y132_AQ;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_A6 = CLBLM_L_X74Y129_SLICE_X113Y129_AQ;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_B1 = CLBLM_L_X78Y130_SLICE_X120Y130_DO6;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_B2 = CLBLL_R_X77Y130_SLICE_X119Y130_BQ;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_B4 = CLBLL_R_X77Y130_SLICE_X119Y130_DO6;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_B5 = CLBLM_L_X78Y130_SLICE_X120Y130_AQ;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_B6 = CLBLM_L_X78Y130_SLICE_X120Y130_BQ;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_B2 = CLBLM_L_X78Y131_SLICE_X120Y131_AQ;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_B4 = CLBLL_R_X77Y130_SLICE_X118Y130_AQ;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_C1 = CLBLL_R_X77Y128_SLICE_X119Y128_BQ;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_C2 = CLBLL_R_X77Y130_SLICE_X118Y130_AQ;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_C3 = CLBLM_L_X78Y131_SLICE_X120Y131_AQ;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_C4 = CLBLL_R_X77Y130_SLICE_X119Y130_AO5;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_C5 = CLBLL_R_X77Y130_SLICE_X119Y130_DO6;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_C6 = CLBLM_L_X78Y129_SLICE_X120Y129_BO6;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_C1 = CLBLL_R_X77Y129_SLICE_X119Y129_BQ;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_C2 = 1'b1;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_C4 = CLBLM_L_X78Y131_SLICE_X120Y131_AQ;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_C5 = CLBLM_L_X76Y130_SLICE_X116Y130_DQ;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_C6 = CLBLL_R_X77Y130_SLICE_X118Y130_AQ;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_D1 = CLBLL_R_X77Y128_SLICE_X118Y128_AQ;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_D2 = 1'b1;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_D3 = 1'b1;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_D4 = CLBLL_R_X77Y130_SLICE_X119Y130_AQ;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_D5 = 1'b1;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_D6 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_D1 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_D2 = 1'b1;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_A2 = CLBLM_L_X64Y105_SLICE_X97Y105_BQ;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_A3 = CLBLM_L_X64Y105_SLICE_X97Y105_AQ;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_A4 = CLBLM_R_X65Y104_SLICE_X98Y104_CQ;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_A5 = CLBLM_R_X65Y104_SLICE_X98Y104_C5Q;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_A6 = CLBLM_R_X65Y104_SLICE_X99Y104_DO6;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_A2 = CLBLM_L_X74Y127_SLICE_X113Y127_A5Q;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_A3 = CLBLM_L_X74Y129_SLICE_X112Y129_AQ;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_B1 = CLBLM_R_X65Y104_SLICE_X99Y104_DO6;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_B2 = CLBLM_R_X65Y104_SLICE_X98Y104_CQ;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_B3 = CLBLM_R_X65Y104_SLICE_X98Y104_C5Q;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_B4 = CLBLM_L_X64Y105_SLICE_X97Y105_DO6;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_B6 = CLBLM_R_X63Y105_SLICE_X95Y105_DO6;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_B1 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_B2 = 1'b1;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_C2 = CLBLM_L_X64Y105_SLICE_X97Y105_CQ;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_C3 = CLBLM_L_X64Y105_SLICE_X96Y105_C5Q;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_C4 = CLBLM_L_X64Y105_SLICE_X96Y105_CQ;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_C5 = CLBLM_L_X64Y102_SLICE_X96Y102_A5Q;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_C6 = CLBLM_L_X64Y104_SLICE_X96Y104_CQ;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_A3 = CLBLM_L_X70Y128_SLICE_X104Y128_AQ;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_A4 = CLBLM_L_X70Y126_SLICE_X105Y126_CO6;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_BX = CLBLL_R_X75Y133_SLICE_X114Y133_AQ;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_C1 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_C2 = 1'b1;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_A5 = CLBLM_L_X70Y128_SLICE_X105Y128_AQ;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_C4 = 1'b1;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_D1 = CLBLM_R_X65Y105_SLICE_X98Y105_AQ;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_D2 = CLBLM_R_X65Y103_SLICE_X99Y103_CO6;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_D3 = 1'b1;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_D4 = CLBLM_L_X64Y105_SLICE_X97Y105_AQ;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_D5 = CLBLM_R_X65Y104_SLICE_X98Y104_C5Q;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_D6 = CLBLM_R_X65Y104_SLICE_X98Y104_CQ;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_A6 = 1'b1;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_D1 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_D2 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_D3 = 1'b1;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_A1 = CLBLM_L_X64Y106_SLICE_X97Y106_B5Q;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_A2 = 1'b1;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_A3 = CLBLM_L_X64Y106_SLICE_X97Y106_AQ;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_A4 = 1'b1;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_A5 = 1'b1;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_A6 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign LIOB33_X0Y183_IOB_X0Y183_O = CLBLM_L_X70Y125_SLICE_X104Y125_DO6;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_B1 = CLBLM_L_X64Y106_SLICE_X97Y106_B5Q;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_B2 = 1'b1;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_B3 = CLBLM_L_X64Y106_SLICE_X97Y106_AQ;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_B4 = 1'b1;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_B5 = 1'b1;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_B6 = 1'b1;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_C1 = CLBLM_L_X64Y105_SLICE_X96Y105_C5Q;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_C2 = CLBLM_L_X64Y105_SLICE_X96Y105_CQ;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_C3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_C4 = CLBLM_L_X64Y102_SLICE_X96Y102_A5Q;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_C5 = 1'b1;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_C6 = 1'b1;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_B3 = CLBLM_L_X70Y128_SLICE_X104Y128_AQ;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_B4 = CLBLM_L_X70Y126_SLICE_X105Y126_CO6;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_D1 = 1'b1;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_D2 = 1'b1;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_D3 = 1'b1;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_D4 = 1'b1;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_D5 = 1'b1;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_D6 = 1'b1;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_B5 = CLBLM_L_X70Y129_SLICE_X104Y129_AQ;
  assign CLBLM_L_X76Y119_SLICE_X116Y119_D5 = 1'b1;
  assign CLBLM_R_X103Y75_SLICE_X163Y75_B5 = 1'b1;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X67Y108_SLICE_X101Y108_A4 = CLBLM_L_X70Y106_SLICE_X105Y106_DO6;
  assign CLBLM_R_X67Y108_SLICE_X101Y108_A5 = CLBLM_L_X62Y92_SLICE_X92Y92_BQ;
  assign CLBLM_R_X67Y108_SLICE_X101Y108_A6 = 1'b1;
  assign CLBLM_R_X67Y108_SLICE_X101Y108_B3 = CLBLM_R_X67Y111_SLICE_X101Y111_B5Q;
  assign CLBLM_R_X67Y108_SLICE_X101Y108_B4 = CLBLM_R_X67Y111_SLICE_X101Y111_A5Q;
  assign CLBLM_R_X67Y108_SLICE_X101Y108_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y108_SLICE_X101Y108_B6 = CLBLM_R_X67Y111_SLICE_X100Y111_A5Q;
  assign CLBLM_R_X103Y75_SLICE_X163Y75_B4 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_A1 = CLBLL_R_X77Y130_SLICE_X119Y130_AQ;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_A2 = CLBLL_R_X77Y128_SLICE_X118Y128_BQ;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_A3 = CLBLL_R_X77Y128_SLICE_X118Y128_AQ;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_A4 = CLBLM_L_X78Y131_SLICE_X120Y131_AQ;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_A5 = CLBLL_R_X77Y130_SLICE_X118Y130_BO6;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_A6 = CLBLL_R_X77Y131_SLICE_X119Y131_DO6;
  assign CLBLM_R_X67Y108_SLICE_X101Y108_C1 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_B1 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_B2 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_B3 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_B4 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_B5 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_B6 = 1'b1;
  assign CLBLM_R_X67Y108_SLICE_X101Y108_C2 = 1'b1;
  assign CLBLM_R_X67Y108_SLICE_X101Y108_C3 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_C1 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_C2 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_C3 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_C4 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_C5 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_C6 = 1'b1;
  assign CLBLM_R_X67Y108_SLICE_X101Y108_C4 = 1'b1;
  assign CLBLM_R_X103Y75_SLICE_X163Y75_B6 = 1'b1;
  assign CLBLM_R_X67Y108_SLICE_X101Y108_C5 = 1'b1;
  assign CLBLM_R_X67Y108_SLICE_X101Y108_C6 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_D1 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_D2 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_D3 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_D4 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_D5 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_D6 = 1'b1;
  assign CLBLM_R_X67Y108_SLICE_X101Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_A1 = CLBLM_L_X78Y130_SLICE_X120Y130_DO6;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_A3 = CLBLL_R_X77Y131_SLICE_X119Y131_AQ;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_A4 = CLBLL_R_X77Y130_SLICE_X119Y130_BQ;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_A5 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_A6 = CLBLL_R_X77Y131_SLICE_X119Y131_CO6;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_B1 = CLBLM_L_X78Y130_SLICE_X120Y130_DO6;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_B2 = CLBLL_R_X77Y131_SLICE_X119Y131_BQ;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_B3 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_B4 = CLBLL_R_X77Y131_SLICE_X119Y131_AQ;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_B6 = CLBLL_R_X77Y131_SLICE_X119Y131_CO6;
  assign CLBLM_R_X67Y108_SLICE_X101Y108_D1 = 1'b1;
  assign CLBLM_R_X67Y108_SLICE_X101Y108_D2 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_C1 = CLBLL_R_X77Y128_SLICE_X118Y128_AQ;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_C2 = CLBLL_R_X77Y130_SLICE_X119Y130_AQ;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_C3 = CLBLM_L_X78Y130_SLICE_X120Y130_AQ;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_C4 = CLBLM_L_X78Y130_SLICE_X120Y130_DO6;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_C5 = CLBLL_R_X77Y130_SLICE_X119Y130_BQ;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_C6 = CLBLM_L_X78Y130_SLICE_X120Y130_BQ;
  assign CLBLM_R_X67Y108_SLICE_X101Y108_D3 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X67Y108_SLICE_X101Y108_D4 = 1'b1;
  assign CLBLM_R_X67Y108_SLICE_X101Y108_D5 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_D1 = CLBLM_L_X78Y130_SLICE_X120Y130_BQ;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_D2 = CLBLL_R_X77Y131_SLICE_X119Y131_AQ;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_D3 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_D4 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_D5 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_D6 = 1'b1;
  assign CLBLM_R_X67Y108_SLICE_X101Y108_D6 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_A1 = CLBLM_L_X64Y106_SLICE_X97Y106_B5Q;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_A2 = 1'b1;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_A3 = CLBLM_L_X64Y106_SLICE_X97Y106_AQ;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_A5 = CLBLM_L_X64Y106_SLICE_X97Y106_C5Q;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_A6 = 1'b1;
  assign CLBLM_R_X67Y108_SLICE_X101Y108_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_B1 = CLBLM_L_X64Y106_SLICE_X97Y106_B5Q;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_B2 = CLBLM_L_X64Y106_SLICE_X97Y106_BQ;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_B4 = 1'b1;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_B5 = CLBLM_L_X64Y106_SLICE_X97Y106_C5Q;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_B6 = 1'b1;
  assign LIOB33_X0Y185_IOB_X0Y186_O = 1'b1;
  assign LIOB33_X0Y185_IOB_X0Y185_O = 1'b1;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_C1 = CLBLM_L_X64Y106_SLICE_X97Y106_C5Q;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_C2 = CLBLM_L_X64Y106_SLICE_X97Y106_CQ;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_C3 = CLBLM_L_X64Y106_SLICE_X97Y106_BQ;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_C4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X60Y94_SLICE_X91Y94_A1 = 1'b1;
  assign CLBLM_L_X60Y94_SLICE_X91Y94_A2 = 1'b1;
  assign CLBLM_L_X60Y94_SLICE_X91Y94_A3 = 1'b1;
  assign CLBLM_L_X60Y94_SLICE_X91Y94_A4 = 1'b1;
  assign CLBLM_L_X60Y94_SLICE_X91Y94_A5 = 1'b1;
  assign CLBLM_L_X60Y94_SLICE_X91Y94_A6 = 1'b1;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_C5 = 1'b1;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_C6 = 1'b1;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X60Y94_SLICE_X91Y94_B1 = 1'b1;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_D1 = 1'b1;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_D2 = 1'b1;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_D3 = 1'b1;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_D4 = 1'b1;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_D5 = 1'b1;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_D6 = 1'b1;
  assign CLBLM_L_X60Y94_SLICE_X91Y94_B2 = 1'b1;
  assign CLBLM_L_X60Y94_SLICE_X91Y94_B3 = 1'b1;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X60Y94_SLICE_X91Y94_B4 = 1'b1;
  assign CLBLM_L_X60Y94_SLICE_X91Y94_B5 = 1'b1;
  assign CLBLM_L_X60Y94_SLICE_X91Y94_B6 = 1'b1;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_A1 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_A2 = CLBLM_L_X64Y106_SLICE_X97Y106_B5Q;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_A3 = CLBLM_L_X64Y106_SLICE_X96Y106_AQ;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_A4 = CLBLM_L_X64Y106_SLICE_X96Y106_BO6;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_A5 = CLBLM_L_X64Y106_SLICE_X97Y106_AQ;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_A6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X60Y94_SLICE_X91Y94_C2 = 1'b1;
  assign CLBLM_L_X60Y94_SLICE_X91Y94_C3 = 1'b1;
  assign CLBLM_L_X60Y94_SLICE_X91Y94_C4 = 1'b1;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_AX = CLBLM_L_X62Y106_SLICE_X92Y106_BQ;
  assign CLBLM_L_X60Y94_SLICE_X91Y94_C6 = 1'b1;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_B1 = 1'b1;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_B2 = 1'b1;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_B3 = CLBLM_L_X64Y106_SLICE_X97Y106_C5Q;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_B4 = CLBLM_L_X64Y106_SLICE_X97Y106_BQ;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_B5 = CLBLM_L_X64Y106_SLICE_X97Y106_CQ;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_B6 = 1'b1;
  assign CLBLM_L_X60Y94_SLICE_X91Y94_D1 = 1'b1;
  assign CLBLM_L_X60Y94_SLICE_X91Y94_D2 = 1'b1;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_BX = CLBLM_L_X64Y106_SLICE_X96Y106_A5Q;
  assign CLBLM_L_X60Y94_SLICE_X91Y94_D3 = 1'b1;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_C1 = CLBLM_L_X64Y105_SLICE_X96Y105_BO6;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_C2 = CLBLM_L_X64Y106_SLICE_X96Y106_CQ;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_C3 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_C4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_C5 = CLBLM_R_X63Y106_SLICE_X95Y106_CQ;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_C6 = CLBLM_L_X64Y106_SLICE_X96Y106_BO6;
  assign CLBLM_L_X60Y94_SLICE_X90Y94_A1 = 1'b1;
  assign CLBLM_L_X60Y94_SLICE_X90Y94_A2 = 1'b1;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X60Y94_SLICE_X90Y94_A3 = 1'b1;
  assign CLBLM_L_X60Y94_SLICE_X90Y94_A4 = 1'b1;
  assign CLBLM_L_X60Y94_SLICE_X90Y94_A5 = 1'b1;
  assign CLBLM_L_X60Y94_SLICE_X90Y94_A6 = 1'b1;
  assign CLBLM_L_X60Y94_SLICE_X90Y94_AX = CLBLM_L_X60Y92_SLICE_X90Y92_AQ;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_D1 = 1'b1;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_D2 = CLBLM_L_X64Y106_SLICE_X97Y106_BQ;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_D3 = 1'b1;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_D4 = CLBLM_L_X64Y106_SLICE_X97Y106_CQ;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_D5 = 1'b1;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_D6 = 1'b1;
  assign CLBLM_L_X60Y94_SLICE_X90Y94_B1 = 1'b1;
  assign CLBLM_L_X60Y94_SLICE_X90Y94_B2 = 1'b1;
  assign CLBLM_L_X60Y94_SLICE_X90Y94_B3 = 1'b1;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X60Y94_SLICE_X90Y94_B6 = 1'b1;
  assign CLBLM_L_X60Y94_SLICE_X90Y94_C1 = 1'b1;
  assign CLBLM_L_X60Y94_SLICE_X90Y94_C2 = 1'b1;
  assign CLBLM_L_X60Y94_SLICE_X90Y94_C3 = 1'b1;
  assign CLBLM_L_X60Y94_SLICE_X90Y94_BX = CLBLM_L_X62Y95_SLICE_X92Y95_BQ;
  assign CLBLM_L_X60Y94_SLICE_X90Y94_C4 = 1'b1;
  assign CLBLM_L_X60Y94_SLICE_X90Y94_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X60Y94_SLICE_X90Y94_C5 = 1'b1;
  assign CLBLM_L_X60Y94_SLICE_X90Y94_C6 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X128Y98_D5 = 1'b1;
  assign CLBLM_R_X67Y108_SLICE_X100Y108_B5 = CLBLM_R_X67Y108_SLICE_X100Y108_C5Q;
  assign CLBLM_L_X60Y94_SLICE_X90Y94_CX = CLBLM_L_X60Y94_SLICE_X90Y94_BQ;
  assign CLBLM_R_X67Y108_SLICE_X100Y108_B6 = 1'b1;
  assign CLBLM_L_X60Y94_SLICE_X90Y94_D1 = 1'b1;
  assign CLBLM_L_X60Y94_SLICE_X90Y94_D2 = 1'b1;
  assign CLBLM_L_X60Y94_SLICE_X90Y94_D3 = 1'b1;
  assign CLBLM_L_X60Y94_SLICE_X90Y94_D4 = 1'b1;
  assign CLBLM_L_X60Y94_SLICE_X90Y94_D5 = 1'b1;
  assign CLBLM_L_X60Y94_SLICE_X90Y94_D6 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X128Y98_D6 = 1'b1;
  assign CLBLM_L_X60Y94_SLICE_X90Y94_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X82Y98_SLICE_X128Y98_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_A4 = 1'b1;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_A6 = CLBLL_R_X71Y124_SLICE_X106Y124_CO6;
  assign CLBLM_R_X67Y108_SLICE_X100Y108_C5 = CLBLM_R_X67Y108_SLICE_X101Y108_BQ;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X67Y108_SLICE_X100Y108_C6 = 1'b1;
  assign CLBLM_R_X67Y109_SLICE_X101Y109_D4 = CLBLM_R_X67Y109_SLICE_X101Y109_CO6;
  assign CLBLM_R_X67Y108_SLICE_X100Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_B4 = CLBLM_L_X72Y125_SLICE_X109Y125_CO6;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_D1 = CLBLM_L_X76Y118_SLICE_X117Y118_CQ;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_B5 = CLBLM_L_X72Y123_SLICE_X108Y123_A5Q;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_B6 = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_T1 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_D1 = CLBLM_L_X74Y120_SLICE_X112Y120_AO6;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_D1 = CLBLM_R_X67Y118_SLICE_X100Y118_A5Q;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1 = CLBLL_R_X77Y124_SLICE_X118Y124_AO6;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_T1 = 1'b1;
  assign CLBLM_R_X67Y108_SLICE_X100Y108_D4 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_D1 = 1'b1;
  assign CLBLM_R_X67Y108_SLICE_X100Y108_D5 = CLBLM_R_X67Y109_SLICE_X100Y109_CQ;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X106Y98_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y98_SLICE_X106Y98_A2 = CLBLM_L_X72Y98_SLICE_X108Y98_AQ;
  assign CLBLL_R_X71Y98_SLICE_X106Y98_A3 = CLBLL_R_X71Y100_SLICE_X106Y100_AO5;
  assign CLBLL_R_X71Y98_SLICE_X106Y98_A4 = CLBLM_L_X70Y98_SLICE_X104Y98_AQ;
  assign CLBLL_R_X71Y98_SLICE_X106Y98_A5 = CLBLL_R_X71Y98_SLICE_X106Y98_A5Q;
  assign CLBLL_R_X71Y98_SLICE_X106Y98_A6 = 1'b1;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_A1 = CLBLL_R_X75Y128_SLICE_X115Y128_DO6;
  assign CLBLL_R_X71Y98_SLICE_X106Y98_B1 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X106Y98_B2 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X106Y98_B3 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X106Y98_B4 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X106Y98_B5 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X106Y98_B6 = 1'b1;
  assign CLBLM_L_X74Y131_SLICE_X113Y131_A2 = 1'b1;
  assign CLBLM_L_X74Y131_SLICE_X113Y131_A3 = 1'b1;
  assign CLBLM_L_X74Y131_SLICE_X113Y131_A4 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X106Y98_C1 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X106Y98_C2 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X106Y98_C3 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X106Y98_C4 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X106Y98_C5 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X106Y98_C6 = 1'b1;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y131_SLICE_X113Y131_B1 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X106Y98_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X74Y131_SLICE_X113Y131_B2 = 1'b1;
  assign CLBLM_L_X74Y131_SLICE_X113Y131_B3 = 1'b1;
  assign CLBLM_L_X74Y131_SLICE_X113Y131_B4 = 1'b1;
  assign CLBLM_L_X74Y131_SLICE_X113Y131_B5 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_A1 = CLBLM_L_X70Y123_SLICE_X104Y123_A5Q;
  assign CLBLL_R_X71Y98_SLICE_X106Y98_D1 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X106Y98_D2 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X106Y98_D3 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X106Y98_D4 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X106Y98_D5 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X106Y98_D6 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_A2 = CLBLL_R_X71Y108_SLICE_X107Y108_A5Q;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_A3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y98_SLICE_X106Y98_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_A4 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_A5 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_A6 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_B1 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_B2 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_B3 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_B4 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_B5 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_B6 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_C1 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_C2 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_C3 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_C4 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_C5 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_C6 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_A3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y131_SLICE_X112Y131_A1 = 1'b1;
  assign CLBLM_L_X74Y131_SLICE_X112Y131_A2 = 1'b1;
  assign CLBLM_L_X74Y131_SLICE_X112Y131_A3 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_D1 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_D2 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X107Y98_A1 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X107Y98_A2 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X107Y98_A3 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X107Y98_A4 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X107Y98_A5 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X107Y98_A6 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_D3 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_D4 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_D5 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X107Y98_B1 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X107Y98_B2 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X107Y98_B3 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X107Y98_B4 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X107Y98_B5 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X107Y98_B6 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_A2 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_A4 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_A5 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X107Y98_C1 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X107Y98_C2 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X107Y98_C3 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X107Y98_C4 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X107Y98_C5 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X107Y98_C6 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_B4 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_B6 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_B1 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_B2 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_B3 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_B5 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_C2 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X107Y98_D1 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X107Y98_D2 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X107Y98_D3 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X107Y98_D4 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X107Y98_D5 = 1'b1;
  assign CLBLL_R_X71Y98_SLICE_X107Y98_D6 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_C3 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_C4 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_C5 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_C6 = 1'b1;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_A5 = CLBLM_L_X74Y129_SLICE_X112Y129_AQ;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_D1 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_D2 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_D3 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_D4 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_D5 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_D6 = 1'b1;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_A6 = 1'b1;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_AX = CLBLL_R_X71Y127_SLICE_X107Y127_AQ;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_D4 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_D5 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_D6 = 1'b1;
  assign LIOI3_X0Y85_OLOGIC_X0Y86_D1 = CLBLM_L_X70Y100_SLICE_X105Y100_CQ;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_B1 = CLBLM_L_X74Y127_SLICE_X112Y127_DO6;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_B2 = CLBLM_L_X74Y128_SLICE_X112Y128_CQ;
  assign CLBLM_L_X74Y132_SLICE_X113Y132_A1 = CLBLM_L_X74Y133_SLICE_X112Y133_CQ;
  assign CLBLM_L_X74Y132_SLICE_X113Y132_A2 = CLBLM_L_X74Y133_SLICE_X113Y133_AO6;
  assign CLBLM_L_X74Y132_SLICE_X113Y132_A3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y132_SLICE_X113Y132_A4 = CLBLM_L_X74Y133_SLICE_X112Y133_DO5;
  assign CLBLM_L_X74Y132_SLICE_X113Y132_A5 = CLBLM_L_X74Y132_SLICE_X113Y132_BQ;
  assign CLBLM_L_X74Y132_SLICE_X113Y132_A6 = CLBLM_L_X74Y132_SLICE_X113Y132_CO6;
  assign LIOB33_X0Y189_IOB_X0Y189_O = 1'b1;
  assign LIOB33_X0Y189_IOB_X0Y190_O = 1'b1;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_B3 = CLBLM_L_X72Y127_SLICE_X108Y127_AQ;
  assign CLBLM_L_X74Y132_SLICE_X113Y132_B1 = CLBLM_L_X74Y133_SLICE_X112Y133_DO5;
  assign CLBLM_L_X74Y132_SLICE_X113Y132_B2 = CLBLM_L_X74Y132_SLICE_X113Y132_BQ;
  assign CLBLM_L_X74Y132_SLICE_X113Y132_B3 = CLBLM_L_X74Y132_SLICE_X113Y132_AQ;
  assign CLBLM_L_X74Y132_SLICE_X113Y132_B4 = CLBLM_L_X74Y134_SLICE_X113Y134_BQ;
  assign CLBLM_L_X74Y132_SLICE_X113Y132_B5 = CLBLM_L_X74Y132_SLICE_X112Y132_AQ;
  assign CLBLM_L_X74Y132_SLICE_X113Y132_B6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y132_SLICE_X113Y132_C1 = CLBLM_L_X74Y132_SLICE_X112Y132_AQ;
  assign CLBLM_L_X74Y132_SLICE_X113Y132_C2 = CLBLM_L_X74Y132_SLICE_X112Y132_A5Q;
  assign CLBLM_L_X74Y132_SLICE_X113Y132_C3 = CLBLM_L_X74Y129_SLICE_X112Y129_BQ;
  assign CLBLM_L_X74Y132_SLICE_X113Y132_C4 = CLBLM_L_X74Y134_SLICE_X113Y134_A5Q;
  assign CLBLM_L_X74Y132_SLICE_X113Y132_C5 = CLBLM_L_X74Y134_SLICE_X113Y134_CQ;
  assign CLBLM_L_X74Y132_SLICE_X113Y132_C6 = CLBLM_L_X74Y132_SLICE_X113Y132_AQ;
  assign LIOI3_X0Y85_OLOGIC_X0Y86_T1 = 1'b1;
  assign CLBLM_L_X74Y132_SLICE_X113Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_B4 = CLBLM_L_X74Y128_SLICE_X112Y128_BQ;
  assign CLBLM_L_X74Y132_SLICE_X113Y132_D1 = 1'b1;
  assign CLBLM_L_X74Y132_SLICE_X113Y132_D2 = 1'b1;
  assign CLBLM_L_X74Y132_SLICE_X113Y132_D3 = 1'b1;
  assign CLBLM_L_X74Y132_SLICE_X113Y132_D4 = 1'b1;
  assign CLBLM_L_X74Y132_SLICE_X113Y132_D5 = 1'b1;
  assign CLBLM_L_X74Y132_SLICE_X113Y132_D6 = 1'b1;
  assign CLBLM_L_X74Y132_SLICE_X113Y132_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y132_SLICE_X112Y132_A1 = CLBLM_L_X74Y134_SLICE_X113Y134_BQ;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_B6 = 1'b1;
  assign CLBLM_L_X74Y132_SLICE_X112Y132_A2 = CLBLM_L_X74Y134_SLICE_X113Y134_CQ;
  assign CLBLM_L_X74Y132_SLICE_X112Y132_A3 = CLBLM_L_X74Y132_SLICE_X112Y132_AQ;
  assign CLBLM_L_X74Y132_SLICE_X112Y132_A4 = CLBLM_L_X74Y129_SLICE_X112Y129_BQ;
  assign CLBLM_L_X74Y132_SLICE_X112Y132_A5 = CLBLM_L_X74Y134_SLICE_X113Y134_A5Q;
  assign CLBLM_L_X74Y132_SLICE_X112Y132_A6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y132_SLICE_X112Y132_AX = CLBLM_L_X74Y132_SLICE_X112Y132_BO5;
  assign CLBLM_L_X74Y132_SLICE_X112Y132_B1 = CLBLM_L_X74Y134_SLICE_X113Y134_BQ;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_B5 = CLBLM_L_X74Y127_SLICE_X112Y127_CO6;
  assign CLBLM_L_X74Y132_SLICE_X112Y132_B2 = CLBLM_L_X74Y133_SLICE_X112Y133_DO5;
  assign CLBLM_L_X74Y132_SLICE_X112Y132_B3 = CLBLM_L_X74Y132_SLICE_X112Y132_AQ;
  assign CLBLM_L_X74Y132_SLICE_X112Y132_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y132_SLICE_X112Y132_B5 = CLBLM_L_X74Y132_SLICE_X112Y132_A5Q;
  assign CLBLM_L_X74Y132_SLICE_X112Y132_B6 = 1'b1;
  assign CLBLM_L_X70Y108_SLICE_X105Y108_C5 = 1'b1;
  assign CLBLM_L_X74Y132_SLICE_X112Y132_C1 = CLBLM_L_X74Y131_SLICE_X112Y131_AQ;
  assign CLBLM_L_X70Y108_SLICE_X105Y108_C6 = 1'b1;
  assign CLBLM_L_X74Y132_SLICE_X112Y132_C2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y132_SLICE_X112Y132_C3 = CLBLL_R_X73Y131_SLICE_X110Y131_AQ;
  assign CLBLM_L_X74Y132_SLICE_X112Y132_C4 = CLBLM_L_X70Y136_SLICE_X105Y136_A5Q;
  assign CLBLM_L_X74Y132_SLICE_X112Y132_C5 = 1'b1;
  assign CLBLM_L_X74Y132_SLICE_X112Y132_C6 = 1'b1;
  assign CLBLM_R_X103Y69_SLICE_X163Y69_B3 = 1'b1;
  assign CLBLM_L_X74Y132_SLICE_X112Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_X0Y85_OLOGIC_X0Y85_D1 = CLBLM_L_X60Y94_SLICE_X90Y94_BQ;
  assign CLBLM_L_X74Y132_SLICE_X112Y132_D1 = 1'b1;
  assign CLBLM_L_X74Y132_SLICE_X112Y132_D2 = 1'b1;
  assign CLBLM_L_X74Y132_SLICE_X112Y132_D3 = 1'b1;
  assign CLBLM_L_X74Y132_SLICE_X112Y132_D4 = 1'b1;
  assign CLBLM_L_X74Y132_SLICE_X112Y132_D5 = 1'b1;
  assign CLBLM_L_X74Y132_SLICE_X112Y132_D6 = 1'b1;
  assign CLBLM_L_X74Y132_SLICE_X112Y132_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_C5 = CLBLM_L_X74Y118_SLICE_X112Y118_BO5;
  assign CLBLM_R_X103Y69_SLICE_X163Y69_B4 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_C6 = CLBLL_R_X75Y124_SLICE_X115Y124_BQ;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X103Y69_SLICE_X163Y69_B5 = 1'b1;
  assign LIOI3_X0Y85_OLOGIC_X0Y85_T1 = 1'b1;
  assign RIOB33_X105Y117_IOB_X1Y118_O = CLBLM_L_X70Y136_SLICE_X105Y136_A5Q;
  assign RIOB33_X105Y117_IOB_X1Y117_O = CLBLL_R_X73Y118_SLICE_X111Y118_AQ;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_D4 = 1'b1;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_A4 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_D5 = 1'b1;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_A5 = 1'b1;
  assign CLBLM_L_X70Y108_SLICE_X104Y108_A1 = 1'b1;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_A6 = 1'b1;
  assign CLBLM_L_X70Y108_SLICE_X104Y108_A2 = 1'b1;
  assign CLBLM_L_X70Y108_SLICE_X104Y108_A3 = 1'b1;
  assign CLBLM_L_X70Y108_SLICE_X104Y108_A4 = 1'b1;
  assign CLBLM_L_X70Y108_SLICE_X104Y108_A5 = 1'b1;
  assign CLBLM_L_X70Y108_SLICE_X104Y108_A6 = 1'b1;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_C3 = CLBLL_R_X75Y122_SLICE_X114Y122_AQ;
  assign LIOB33_X0Y183_IOB_X0Y184_O = CLBLL_R_X73Y134_SLICE_X110Y134_AO5;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_C6 = CLBLM_L_X74Y109_SLICE_X113Y109_AQ;
  assign CLBLM_L_X70Y108_SLICE_X104Y108_B1 = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_D1 = CLBLM_L_X76Y118_SLICE_X117Y118_CQ;
  assign CLBLM_L_X70Y108_SLICE_X104Y108_B2 = 1'b1;
  assign CLBLM_L_X70Y108_SLICE_X104Y108_B3 = 1'b1;
  assign CLBLM_L_X70Y108_SLICE_X104Y108_B4 = 1'b1;
  assign RIOB33_X105Y165_IOB_X1Y166_O = 1'b1;
  assign CLBLM_L_X70Y108_SLICE_X104Y108_B5 = 1'b1;
  assign RIOB33_X105Y165_IOB_X1Y165_O = CLBLM_L_X70Y111_SLICE_X105Y111_DO6;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_C1 = 1'b1;
  assign CLBLM_L_X70Y108_SLICE_X104Y108_B6 = 1'b1;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_C2 = 1'b1;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_C5 = 1'b1;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_D1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign LIOB33_X0Y191_IOB_X0Y192_O = 1'b1;
  assign LIOB33_X0Y191_IOB_X0Y191_O = 1'b1;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_C6 = 1'b1;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_D2 = CLBLL_R_X77Y124_SLICE_X119Y124_CQ;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_D3 = CLBLL_R_X75Y122_SLICE_X114Y122_AQ;
  assign CLBLL_R_X71Y100_SLICE_X106Y100_A1 = CLBLL_R_X77Y108_SLICE_X118Y108_AQ;
  assign CLBLL_R_X71Y100_SLICE_X106Y100_A2 = CLBLL_R_X71Y100_SLICE_X106Y100_BQ;
  assign CLBLL_R_X71Y100_SLICE_X106Y100_A3 = CLBLM_L_X60Y99_SLICE_X90Y99_AQ;
  assign CLBLL_R_X71Y100_SLICE_X106Y100_A4 = CLBLM_L_X70Y100_SLICE_X105Y100_CQ;
  assign CLBLL_R_X71Y100_SLICE_X106Y100_A5 = CLBLL_R_X71Y98_SLICE_X106Y98_A5Q;
  assign CLBLL_R_X71Y100_SLICE_X106Y100_A6 = 1'b1;
  assign CLBLM_L_X70Y108_SLICE_X104Y108_C1 = 1'b1;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_D4 = CLBLM_L_X76Y125_SLICE_X117Y125_BQ;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_D5 = CLBLM_L_X76Y118_SLICE_X117Y118_CQ;
  assign CLBLL_R_X71Y100_SLICE_X106Y100_B1 = CLBLL_R_X77Y108_SLICE_X118Y108_AQ;
  assign CLBLL_R_X71Y100_SLICE_X106Y100_B2 = CLBLL_R_X71Y100_SLICE_X106Y100_BQ;
  assign CLBLL_R_X71Y100_SLICE_X106Y100_B3 = CLBLL_R_X71Y100_SLICE_X106Y100_DO6;
  assign CLBLL_R_X71Y100_SLICE_X106Y100_B4 = CLBLM_L_X60Y97_SLICE_X90Y97_BQ;
  assign CLBLL_R_X71Y100_SLICE_X106Y100_B5 = CLBLM_L_X70Y100_SLICE_X105Y100_CQ;
  assign CLBLL_R_X71Y100_SLICE_X106Y100_B6 = CLBLM_L_X60Y99_SLICE_X90Y99_AQ;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_D6 = 1'b1;
  assign CLBLM_R_X103Y69_SLICE_X163Y69_C2 = 1'b1;
  assign CLBLM_L_X74Y133_SLICE_X113Y133_A1 = CLBLM_L_X76Y133_SLICE_X116Y133_BQ;
  assign CLBLL_R_X71Y100_SLICE_X106Y100_C1 = CLBLM_L_X70Y100_SLICE_X105Y100_CQ;
  assign CLBLL_R_X71Y100_SLICE_X106Y100_C2 = CLBLL_R_X71Y101_SLICE_X106Y101_BQ;
  assign CLBLL_R_X71Y100_SLICE_X106Y100_C3 = CLBLM_L_X70Y100_SLICE_X105Y100_A5Q;
  assign CLBLL_R_X71Y100_SLICE_X106Y100_C4 = CLBLM_L_X60Y99_SLICE_X90Y99_AQ;
  assign CLBLL_R_X71Y100_SLICE_X106Y100_C5 = CLBLL_R_X71Y101_SLICE_X106Y101_CQ;
  assign CLBLL_R_X71Y100_SLICE_X106Y100_C6 = CLBLM_L_X70Y100_SLICE_X105Y100_AQ;
  assign CLBLM_L_X70Y108_SLICE_X104Y108_C6 = 1'b1;
  assign CLBLM_L_X74Y133_SLICE_X113Y133_A2 = CLBLL_R_X73Y133_SLICE_X110Y133_CQ;
  assign CLBLL_R_X71Y100_SLICE_X106Y100_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y133_SLICE_X113Y133_A3 = CLBLL_R_X75Y133_SLICE_X115Y133_AQ;
  assign CLBLM_L_X74Y133_SLICE_X113Y133_B2 = 1'b1;
  assign CLBLM_L_X74Y133_SLICE_X113Y133_B3 = 1'b1;
  assign CLBLM_L_X74Y133_SLICE_X113Y133_B4 = 1'b1;
  assign CLBLM_L_X74Y133_SLICE_X113Y133_B5 = 1'b1;
  assign CLBLL_R_X71Y100_SLICE_X106Y100_D1 = CLBLM_L_X70Y100_SLICE_X105Y100_CQ;
  assign CLBLL_R_X71Y100_SLICE_X106Y100_D2 = CLBLM_L_X70Y100_SLICE_X104Y100_A5Q;
  assign CLBLL_R_X71Y100_SLICE_X106Y100_D3 = CLBLL_R_X71Y100_SLICE_X106Y100_BQ;
  assign CLBLL_R_X71Y100_SLICE_X106Y100_D4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y100_SLICE_X106Y100_D5 = CLBLL_R_X77Y108_SLICE_X118Y108_AQ;
  assign CLBLL_R_X71Y100_SLICE_X106Y100_D6 = CLBLM_L_X60Y97_SLICE_X90Y97_BQ;
  assign CLBLM_L_X74Y133_SLICE_X113Y133_B6 = 1'b1;
  assign CLBLL_R_X71Y100_SLICE_X106Y100_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y133_SLICE_X113Y133_C1 = 1'b1;
  assign CLBLM_L_X74Y133_SLICE_X113Y133_C2 = 1'b1;
  assign CLBLM_L_X74Y133_SLICE_X113Y133_C3 = 1'b1;
  assign CLBLM_L_X74Y133_SLICE_X113Y133_C4 = 1'b1;
  assign CLBLM_L_X74Y133_SLICE_X113Y133_C5 = 1'b1;
  assign CLBLM_L_X74Y133_SLICE_X113Y133_C6 = 1'b1;
  assign CLBLM_L_X74Y133_SLICE_X113Y133_D1 = 1'b1;
  assign CLBLM_L_X74Y133_SLICE_X113Y133_D2 = 1'b1;
  assign CLBLM_L_X74Y133_SLICE_X113Y133_D3 = 1'b1;
  assign CLBLM_L_X74Y133_SLICE_X113Y133_D4 = 1'b1;
  assign CLBLM_L_X74Y133_SLICE_X113Y133_D5 = 1'b1;
  assign CLBLM_L_X74Y133_SLICE_X113Y133_D6 = 1'b1;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_A1 = CLBLL_R_X79Y127_SLICE_X122Y127_BQ;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X103Y69_SLICE_X163Y69_C4 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_D1 = CLBLM_R_X67Y116_SLICE_X100Y116_AQ;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_A3 = CLBLM_L_X76Y125_SLICE_X116Y125_AQ;
  assign CLBLM_L_X74Y133_SLICE_X112Y133_A1 = CLBLM_L_X74Y134_SLICE_X112Y134_AO5;
  assign CLBLM_L_X74Y133_SLICE_X112Y133_A2 = CLBLM_L_X74Y134_SLICE_X113Y134_BQ;
  assign CLBLM_L_X74Y133_SLICE_X112Y133_A3 = CLBLM_L_X74Y133_SLICE_X112Y133_AQ;
  assign CLBLL_R_X71Y100_SLICE_X107Y100_A1 = 1'b1;
  assign CLBLL_R_X71Y100_SLICE_X107Y100_A2 = 1'b1;
  assign CLBLL_R_X71Y100_SLICE_X107Y100_A3 = 1'b1;
  assign CLBLL_R_X71Y100_SLICE_X107Y100_A4 = 1'b1;
  assign CLBLL_R_X71Y100_SLICE_X107Y100_A5 = 1'b1;
  assign CLBLL_R_X71Y100_SLICE_X107Y100_A6 = 1'b1;
  assign CLBLM_L_X74Y133_SLICE_X112Y133_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y133_SLICE_X112Y133_A5 = CLBLM_L_X74Y132_SLICE_X112Y132_AQ;
  assign CLBLM_L_X74Y133_SLICE_X112Y133_A6 = CLBLL_R_X73Y133_SLICE_X111Y133_AQ;
  assign CLBLL_R_X71Y100_SLICE_X107Y100_B1 = 1'b1;
  assign CLBLL_R_X71Y100_SLICE_X107Y100_B2 = 1'b1;
  assign CLBLL_R_X71Y100_SLICE_X107Y100_B3 = 1'b1;
  assign CLBLL_R_X71Y100_SLICE_X107Y100_B4 = 1'b1;
  assign CLBLL_R_X71Y100_SLICE_X107Y100_B5 = 1'b1;
  assign CLBLL_R_X71Y100_SLICE_X107Y100_B6 = 1'b1;
  assign CLBLM_L_X74Y133_SLICE_X112Y133_B1 = CLBLM_L_X74Y133_SLICE_X112Y133_DO6;
  assign CLBLM_L_X74Y133_SLICE_X112Y133_B2 = CLBLM_L_X74Y133_SLICE_X112Y133_BQ;
  assign CLBLM_L_X74Y133_SLICE_X112Y133_B3 = CLBLM_L_X74Y133_SLICE_X112Y133_AQ;
  assign CLBLL_R_X71Y100_SLICE_X107Y100_C1 = 1'b1;
  assign CLBLL_R_X71Y100_SLICE_X107Y100_C2 = 1'b1;
  assign CLBLL_R_X71Y100_SLICE_X107Y100_C3 = 1'b1;
  assign CLBLL_R_X71Y100_SLICE_X107Y100_C4 = 1'b1;
  assign CLBLL_R_X71Y100_SLICE_X107Y100_C5 = 1'b1;
  assign CLBLL_R_X71Y100_SLICE_X107Y100_C6 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_A1 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_A2 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_A3 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_A4 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_A5 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_A6 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_AX = CLBLM_R_X65Y110_SLICE_X99Y110_B5Q;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_B4 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_B1 = 1'b1;
  assign CLBLL_R_X71Y100_SLICE_X107Y100_D1 = 1'b1;
  assign CLBLL_R_X71Y100_SLICE_X107Y100_D2 = 1'b1;
  assign CLBLL_R_X71Y100_SLICE_X107Y100_D3 = 1'b1;
  assign CLBLL_R_X71Y100_SLICE_X107Y100_D4 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_C1 = 1'b1;
  assign CLBLL_R_X71Y100_SLICE_X107Y100_D5 = 1'b1;
  assign CLBLL_R_X71Y100_SLICE_X107Y100_D6 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_B6 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X122Y96_A1 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X122Y96_A2 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X122Y96_A3 = CLBLM_R_X103Y69_SLICE_X162Y69_A5Q;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLL_R_X79Y96_SLICE_X122Y96_A4 = CLBLM_L_X82Y98_SLICE_X128Y98_A5Q;
  assign CLBLL_R_X79Y96_SLICE_X122Y96_A5 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X122Y96_A6 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_C4 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_C6 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X122Y96_B1 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X122Y96_B2 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_D3 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_D4 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_D5 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_D6 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X122Y96_B3 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X122Y96_B4 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X79Y96_SLICE_X122Y96_B5 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X122Y96_B6 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_A1 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_A2 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_A3 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_A4 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_A5 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_A6 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X122Y96_C1 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X122Y96_C2 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X122Y96_C3 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_AX = CLBLM_L_X62Y107_SLICE_X93Y107_A5Q;
  assign CLBLL_R_X79Y96_SLICE_X122Y96_C5 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_B1 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_B2 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_B3 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_B4 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_B5 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_B6 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X122Y96_D1 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X122Y96_D2 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_BX = CLBLM_L_X60Y99_SLICE_X90Y99_AQ;
  assign CLBLL_R_X79Y96_SLICE_X122Y96_D3 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_C2 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X122Y96_D4 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_C4 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_C5 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_C6 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_C1 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_C3 = 1'b1;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_C1 = CLBLM_R_X65Y105_SLICE_X99Y105_CQ;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_C2 = CLBLM_L_X76Y125_SLICE_X116Y125_CQ;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_A3 = CLBLM_L_X70Y129_SLICE_X105Y129_AQ;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_CX = CLBLM_R_X63Y98_SLICE_X94Y98_BQ;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_C3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_D1 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_D2 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_D3 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_D4 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_D5 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_D6 = 1'b1;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_A4 = CLBLM_L_X70Y130_SLICE_X105Y130_A5Q;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_C4 = CLBLL_R_X77Y127_SLICE_X119Y127_AO5;
  assign CLBLL_R_X79Y96_SLICE_X123Y96_A1 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X123Y96_A2 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X123Y96_A3 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X123Y96_A4 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X123Y96_A5 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X123Y96_A6 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_DX = CLBLM_L_X68Y97_SLICE_X103Y97_AQ;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_C6 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X123Y96_B1 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X123Y96_B2 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X123Y96_B3 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X123Y96_B4 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X123Y96_B5 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X123Y96_B6 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X123Y96_C1 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X123Y96_C2 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X123Y96_C3 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X123Y96_C4 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X123Y96_C5 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X123Y96_C6 = 1'b1;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X79Y96_SLICE_X123Y96_D1 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X123Y96_D2 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X123Y96_D3 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X123Y96_D4 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X123Y96_D5 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X123Y96_D6 = 1'b1;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_B4 = CLBLM_L_X72Y132_SLICE_X109Y132_AO6;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_B6 = CLBLM_L_X72Y133_SLICE_X109Y133_AO6;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_D1 = 1'b1;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_D2 = 1'b1;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_D3 = 1'b1;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_D4 = 1'b1;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_D5 = 1'b1;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_D6 = 1'b1;
  assign LIOB33_X0Y193_IOB_X0Y194_O = 1'b1;
  assign LIOB33_X0Y193_IOB_X0Y193_O = 1'b1;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X103Y75_SLICE_X163Y75_C6 = 1'b1;
  assign CLBLM_R_X67Y115_SLICE_X101Y115_B4 = 1'b1;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_D1 = 1'b1;
  assign CLBLL_R_X71Y101_SLICE_X106Y101_A1 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLL_R_X71Y101_SLICE_X106Y101_A2 = CLBLM_L_X70Y101_SLICE_X104Y101_CQ;
  assign CLBLL_R_X71Y101_SLICE_X106Y101_A3 = CLBLL_R_X71Y101_SLICE_X106Y101_AQ;
  assign CLBLL_R_X71Y101_SLICE_X106Y101_A4 = CLBLM_L_X70Y103_SLICE_X104Y103_DO5;
  assign CLBLL_R_X71Y101_SLICE_X106Y101_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y101_SLICE_X106Y101_A6 = CLBLM_L_X70Y103_SLICE_X105Y103_CO5;
  assign CLBLL_R_X71Y101_SLICE_X106Y101_B1 = CLBLM_L_X70Y103_SLICE_X105Y103_DO6;
  assign CLBLL_R_X71Y101_SLICE_X106Y101_B2 = CLBLL_R_X71Y101_SLICE_X106Y101_BQ;
  assign CLBLL_R_X71Y101_SLICE_X106Y101_B3 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLL_R_X71Y101_SLICE_X106Y101_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y101_SLICE_X106Y101_B5 = CLBLL_R_X71Y102_SLICE_X106Y102_BQ;
  assign CLBLL_R_X71Y101_SLICE_X106Y101_B6 = CLBLL_R_X71Y103_SLICE_X106Y103_BO6;
  assign CLBLM_L_X72Y130_SLICE_X108Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X71Y101_SLICE_X106Y101_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y101_SLICE_X106Y101_C2 = CLBLL_R_X71Y101_SLICE_X106Y101_CQ;
  assign CLBLL_R_X71Y101_SLICE_X106Y101_C3 = CLBLL_R_X71Y101_SLICE_X106Y101_BQ;
  assign CLBLL_R_X71Y101_SLICE_X106Y101_C4 = CLBLM_L_X70Y103_SLICE_X105Y103_DO5;
  assign CLBLL_R_X71Y101_SLICE_X106Y101_C5 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLL_R_X71Y101_SLICE_X106Y101_C6 = CLBLL_R_X71Y103_SLICE_X106Y103_BO6;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_D2 = 1'b1;
  assign CLBLM_L_X74Y134_SLICE_X113Y134_A1 = CLBLM_L_X74Y134_SLICE_X113Y134_AQ;
  assign CLBLL_R_X71Y101_SLICE_X106Y101_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y134_SLICE_X113Y134_A2 = CLBLM_L_X74Y134_SLICE_X113Y134_BQ;
  assign CLBLM_L_X74Y134_SLICE_X113Y134_A3 = CLBLM_L_X74Y134_SLICE_X112Y134_AO6;
  assign CLBLM_L_X74Y134_SLICE_X113Y134_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y134_SLICE_X113Y134_A5 = CLBLM_L_X74Y132_SLICE_X112Y132_AQ;
  assign CLBLM_L_X74Y134_SLICE_X113Y134_A6 = CLBLL_R_X73Y134_SLICE_X111Y134_AQ;
  assign CLBLL_R_X71Y101_SLICE_X106Y101_D1 = CLBLM_L_X70Y100_SLICE_X105Y100_AQ;
  assign CLBLL_R_X71Y101_SLICE_X106Y101_D2 = CLBLL_R_X71Y102_SLICE_X106Y102_AQ;
  assign CLBLL_R_X71Y101_SLICE_X106Y101_D3 = CLBLL_R_X71Y103_SLICE_X106Y103_AQ;
  assign CLBLL_R_X71Y101_SLICE_X106Y101_D4 = CLBLM_L_X70Y100_SLICE_X105Y100_A5Q;
  assign CLBLL_R_X71Y101_SLICE_X106Y101_D5 = CLBLM_L_X70Y101_SLICE_X104Y101_AQ;
  assign CLBLL_R_X71Y101_SLICE_X106Y101_D6 = CLBLM_L_X70Y100_SLICE_X104Y100_A5Q;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_D3 = CLBLM_L_X70Y129_SLICE_X105Y129_DQ;
  assign CLBLM_L_X74Y134_SLICE_X113Y134_B1 = CLBLM_L_X74Y134_SLICE_X113Y134_CQ;
  assign CLBLL_R_X71Y101_SLICE_X106Y101_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_D4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y134_SLICE_X113Y134_B4 = CLBLM_L_X74Y134_SLICE_X113Y134_A5Q;
  assign CLBLM_L_X74Y134_SLICE_X113Y134_B5 = CLBLM_L_X74Y129_SLICE_X112Y129_BQ;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_D3 = 1'b1;
  assign CLBLM_L_X74Y134_SLICE_X113Y134_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y134_SLICE_X113Y134_C2 = CLBLM_L_X74Y134_SLICE_X113Y134_CQ;
  assign CLBLM_L_X74Y134_SLICE_X113Y134_C3 = CLBLM_L_X74Y134_SLICE_X113Y134_A5Q;
  assign CLBLM_L_X74Y134_SLICE_X113Y134_C4 = CLBLL_R_X75Y133_SLICE_X114Y133_BQ;
  assign CLBLM_L_X74Y134_SLICE_X113Y134_C5 = CLBLL_R_X75Y134_SLICE_X115Y134_CO6;
  assign CLBLM_L_X74Y134_SLICE_X113Y134_C6 = CLBLM_L_X74Y135_SLICE_X113Y135_BQ;
  assign CLBLM_L_X74Y134_SLICE_X113Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y134_SLICE_X113Y134_D1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y134_SLICE_X113Y134_D2 = CLBLL_R_X75Y133_SLICE_X114Y133_BQ;
  assign CLBLM_L_X74Y134_SLICE_X113Y134_D3 = CLBLM_L_X74Y135_SLICE_X113Y135_DO6;
  assign CLBLM_L_X74Y134_SLICE_X113Y134_D4 = CLBLM_L_X74Y134_SLICE_X113Y134_A5Q;
  assign CLBLM_L_X74Y134_SLICE_X113Y134_D5 = CLBLM_L_X74Y134_SLICE_X113Y134_CQ;
  assign CLBLM_L_X74Y134_SLICE_X113Y134_D6 = 1'b1;
  assign CLBLM_L_X74Y134_SLICE_X113Y134_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X71Y101_SLICE_X107Y101_A1 = CLBLM_L_X70Y103_SLICE_X105Y103_DO6;
  assign CLBLL_R_X71Y101_SLICE_X107Y101_A2 = CLBLM_L_X70Y103_SLICE_X105Y103_CO5;
  assign CLBLL_R_X71Y101_SLICE_X107Y101_A3 = CLBLL_R_X71Y101_SLICE_X107Y101_AQ;
  assign CLBLL_R_X71Y101_SLICE_X107Y101_A4 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLL_R_X71Y101_SLICE_X107Y101_A5 = CLBLL_R_X71Y101_SLICE_X106Y101_AQ;
  assign CLBLL_R_X71Y101_SLICE_X107Y101_A6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_D4 = 1'b1;
  assign CLBLM_L_X74Y134_SLICE_X112Y134_A1 = CLBLM_L_X74Y134_SLICE_X113Y134_A5Q;
  assign CLBLM_L_X74Y134_SLICE_X112Y134_A2 = CLBLM_L_X74Y134_SLICE_X113Y134_CQ;
  assign CLBLL_R_X71Y101_SLICE_X107Y101_B1 = 1'b1;
  assign CLBLL_R_X71Y101_SLICE_X107Y101_B2 = 1'b1;
  assign CLBLL_R_X71Y101_SLICE_X107Y101_B3 = 1'b1;
  assign CLBLL_R_X71Y101_SLICE_X107Y101_B4 = 1'b1;
  assign CLBLL_R_X71Y101_SLICE_X107Y101_B5 = 1'b1;
  assign CLBLL_R_X71Y101_SLICE_X107Y101_B6 = 1'b1;
  assign CLBLM_L_X74Y134_SLICE_X112Y134_A6 = 1'b1;
  assign CLBLM_L_X74Y134_SLICE_X112Y134_B1 = CLBLM_L_X74Y132_SLICE_X112Y132_C5Q;
  assign CLBLL_R_X71Y101_SLICE_X107Y101_C1 = 1'b1;
  assign CLBLL_R_X71Y101_SLICE_X107Y101_C2 = 1'b1;
  assign CLBLL_R_X71Y101_SLICE_X107Y101_C3 = 1'b1;
  assign CLBLL_R_X71Y101_SLICE_X107Y101_C4 = 1'b1;
  assign CLBLL_R_X71Y101_SLICE_X107Y101_C5 = 1'b1;
  assign CLBLL_R_X71Y101_SLICE_X107Y101_C6 = 1'b1;
  assign CLBLM_L_X74Y134_SLICE_X112Y134_B5 = 1'b1;
  assign CLBLM_L_X74Y134_SLICE_X112Y134_B6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y101_SLICE_X107Y101_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_D5 = 1'b1;
  assign CLBLM_L_X74Y134_SLICE_X112Y134_C1 = 1'b1;
  assign CLBLM_L_X74Y134_SLICE_X112Y134_C2 = CLBLM_L_X74Y134_SLICE_X112Y134_CQ;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_A3 = CLBLM_L_X70Y129_SLICE_X104Y129_AQ;
  assign CLBLL_R_X71Y101_SLICE_X107Y101_D1 = 1'b1;
  assign CLBLL_R_X71Y101_SLICE_X107Y101_D2 = 1'b1;
  assign CLBLL_R_X71Y101_SLICE_X107Y101_D3 = 1'b1;
  assign CLBLL_R_X71Y101_SLICE_X107Y101_D4 = 1'b1;
  assign CLBLL_R_X71Y101_SLICE_X107Y101_D5 = 1'b1;
  assign CLBLL_R_X71Y101_SLICE_X107Y101_D6 = 1'b1;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_A4 = CLBLM_L_X70Y128_SLICE_X104Y128_AQ;
  assign CLBLL_R_X71Y101_SLICE_X107Y101_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y134_SLICE_X112Y134_D1 = CLBLM_L_X74Y134_SLICE_X113Y134_DO5;
  assign CLBLM_L_X74Y134_SLICE_X112Y134_D2 = CLBLM_L_X74Y132_SLICE_X112Y132_C5Q;
  assign CLBLM_L_X74Y134_SLICE_X112Y134_D3 = CLBLM_L_X74Y134_SLICE_X112Y134_DQ;
  assign CLBLM_L_X74Y134_SLICE_X112Y134_D4 = CLBLM_L_X74Y134_SLICE_X112Y134_BQ;
  assign CLBLM_L_X74Y134_SLICE_X112Y134_D5 = CLBLM_L_X74Y134_SLICE_X113Y134_A5Q;
  assign CLBLM_L_X74Y134_SLICE_X112Y134_D6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y134_SLICE_X112Y134_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_D6 = 1'b1;
  assign CLBLM_R_X67Y115_SLICE_X101Y115_B5 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1 = CLBLL_R_X77Y128_SLICE_X119Y128_BQ;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_B1 = CLBLL_R_X71Y130_SLICE_X106Y130_AO6;
  assign CLBLM_R_X53Y122_SLICE_X81Y122_A1 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X81Y122_A2 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X81Y122_A3 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X81Y122_A4 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X81Y122_A5 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X81Y122_A6 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X81Y122_B1 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X81Y122_B2 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X81Y122_B3 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X81Y122_B4 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X81Y122_B5 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X81Y122_B6 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X81Y122_C1 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X81Y122_C2 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X81Y122_C3 = 1'b1;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X53Y122_SLICE_X81Y122_C4 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X81Y122_C5 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X81Y122_C6 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X81Y122_D1 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X81Y122_D2 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X81Y122_D3 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X81Y122_D4 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X81Y122_D5 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X81Y122_D6 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X80Y122_A1 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X80Y122_A2 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X80Y122_A3 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X80Y122_A4 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X80Y122_A5 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X80Y122_A6 = 1'b1;
  assign CLBLM_R_X67Y109_SLICE_X101Y109_B1 = CLBLM_R_X65Y110_SLICE_X99Y110_AO5;
  assign CLBLM_R_X53Y122_SLICE_X80Y122_AX = CLBLM_R_X63Y122_SLICE_X95Y122_AQ;
  assign CLBLM_R_X67Y109_SLICE_X101Y109_B2 = CLBLM_R_X67Y109_SLICE_X101Y109_BQ;
  assign CLBLM_R_X53Y122_SLICE_X80Y122_B1 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X80Y122_B2 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X80Y122_B3 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X80Y122_B4 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X80Y122_B5 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X80Y122_B6 = 1'b1;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign LIOB33_X0Y195_IOB_X0Y195_O = 1'b1;
  assign LIOB33_X0Y195_IOB_X0Y196_O = CLBLM_L_X64Y105_SLICE_X97Y105_DO6;
  assign CLBLM_R_X53Y122_SLICE_X80Y122_C1 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X80Y122_C2 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X80Y122_C3 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X80Y122_C4 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X80Y122_C5 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X80Y122_C6 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X80Y122_CE = CLBLM_L_X76Y109_SLICE_X116Y109_AO6;
  assign CLBLM_R_X67Y109_SLICE_X101Y109_B5 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X78Y104_SLICE_X120Y104_B4 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X80Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X67Y109_SLICE_X101Y109_B6 = CLBLM_R_X67Y110_SLICE_X101Y110_CQ;
  assign CLBLM_R_X53Y122_SLICE_X80Y122_D1 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X80Y122_D2 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X80Y122_D3 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X80Y122_D4 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X80Y122_D5 = 1'b1;
  assign CLBLM_R_X53Y122_SLICE_X80Y122_D6 = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_D1 = CLBLM_L_X64Y99_SLICE_X97Y99_B5Q;
  assign CLBLM_R_X53Y122_SLICE_X80Y122_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X67Y109_SLICE_X101Y109_C1 = CLBLM_R_X65Y110_SLICE_X99Y110_CQ;
  assign CLBLM_R_X67Y109_SLICE_X101Y109_C2 = CLBLM_R_X67Y110_SLICE_X101Y110_CQ;
  assign CLBLM_R_X67Y109_SLICE_X101Y109_C3 = CLBLM_R_X67Y110_SLICE_X100Y110_CQ;
  assign CLBLM_R_X67Y109_SLICE_X101Y109_C4 = CLBLM_L_X60Y97_SLICE_X91Y97_AQ;
  assign CLBLM_R_X67Y109_SLICE_X101Y109_C5 = CLBLM_L_X68Y109_SLICE_X102Y109_A5Q;
  assign CLBLL_R_X71Y102_SLICE_X106Y102_A1 = CLBLL_R_X71Y103_SLICE_X106Y103_BO5;
  assign CLBLL_R_X71Y102_SLICE_X106Y102_A2 = CLBLM_L_X70Y103_SLICE_X104Y103_DO5;
  assign CLBLL_R_X71Y102_SLICE_X106Y102_A3 = CLBLL_R_X71Y102_SLICE_X106Y102_AQ;
  assign CLBLL_R_X71Y102_SLICE_X106Y102_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y102_SLICE_X106Y102_A5 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLL_R_X71Y102_SLICE_X106Y102_A6 = CLBLL_R_X71Y103_SLICE_X106Y103_AQ;
  assign CLBLM_R_X67Y109_SLICE_X101Y109_C6 = CLBLM_R_X65Y111_SLICE_X98Y111_AQ;
  assign CLBLL_R_X71Y102_SLICE_X106Y102_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y102_SLICE_X106Y102_B2 = CLBLL_R_X71Y102_SLICE_X106Y102_BQ;
  assign CLBLL_R_X71Y102_SLICE_X106Y102_B3 = CLBLL_R_X71Y103_SLICE_X106Y103_BO6;
  assign CLBLL_R_X71Y102_SLICE_X106Y102_B4 = CLBLM_L_X70Y103_SLICE_X104Y103_DO5;
  assign CLBLL_R_X71Y102_SLICE_X106Y102_B5 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLL_R_X71Y102_SLICE_X106Y102_B6 = CLBLM_L_X70Y102_SLICE_X105Y102_AQ;
  assign CLBLM_R_X67Y109_SLICE_X101Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X71Y102_SLICE_X106Y102_C1 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLL_R_X71Y102_SLICE_X106Y102_C2 = CLBLL_R_X71Y102_SLICE_X106Y102_CQ;
  assign CLBLL_R_X71Y102_SLICE_X106Y102_C3 = CLBLL_R_X71Y102_SLICE_X106Y102_AQ;
  assign CLBLL_R_X71Y102_SLICE_X106Y102_C4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y102_SLICE_X106Y102_C5 = CLBLM_L_X70Y103_SLICE_X105Y103_DO6;
  assign CLBLL_R_X71Y102_SLICE_X106Y102_C6 = CLBLL_R_X71Y103_SLICE_X106Y103_BO5;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_D3 = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_T1 = 1'b1;
  assign CLBLL_R_X71Y102_SLICE_X106Y102_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y135_SLICE_X113Y135_A1 = CLBLM_L_X74Y135_SLICE_X113Y135_DO6;
  assign CLBLM_L_X74Y135_SLICE_X113Y135_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y135_SLICE_X113Y135_A3 = CLBLM_L_X74Y135_SLICE_X113Y135_AQ;
  assign CLBLM_L_X74Y135_SLICE_X113Y135_A4 = 1'b1;
  assign CLBLM_L_X74Y135_SLICE_X113Y135_A5 = CLBLM_L_X74Y135_SLICE_X112Y135_AQ;
  assign CLBLL_R_X71Y102_SLICE_X106Y102_D1 = CLBLL_R_X71Y102_SLICE_X106Y102_BQ;
  assign CLBLL_R_X71Y102_SLICE_X106Y102_D2 = CLBLL_R_X71Y102_SLICE_X106Y102_CQ;
  assign CLBLL_R_X71Y102_SLICE_X106Y102_D3 = CLBLL_R_X77Y108_SLICE_X118Y108_AQ;
  assign CLBLL_R_X71Y102_SLICE_X106Y102_D4 = CLBLL_R_X71Y98_SLICE_X106Y98_A5Q;
  assign CLBLL_R_X71Y102_SLICE_X106Y102_D5 = CLBLM_L_X70Y101_SLICE_X105Y101_AQ;
  assign CLBLL_R_X71Y102_SLICE_X106Y102_D6 = CLBLL_R_X71Y100_SLICE_X106Y100_BQ;
  assign CLBLM_L_X74Y135_SLICE_X113Y135_A6 = CLBLM_L_X74Y135_SLICE_X113Y135_CO6;
  assign CLBLL_R_X71Y102_SLICE_X106Y102_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y135_SLICE_X113Y135_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y135_SLICE_X113Y135_B2 = CLBLM_L_X74Y135_SLICE_X112Y135_BO6;
  assign CLBLM_L_X74Y135_SLICE_X113Y135_B3 = CLBLM_L_X74Y135_SLICE_X113Y135_AQ;
  assign CLBLM_L_X74Y135_SLICE_X113Y135_B4 = CLBLL_R_X75Y134_SLICE_X115Y134_CO6;
  assign CLBLM_L_X74Y135_SLICE_X113Y135_B5 = CLBLM_L_X74Y134_SLICE_X112Y134_CQ;
  assign CLBLM_L_X74Y135_SLICE_X113Y135_C2 = CLBLM_L_X74Y134_SLICE_X113Y134_CQ;
  assign CLBLM_L_X74Y135_SLICE_X113Y135_C3 = CLBLM_L_X74Y132_SLICE_X112Y132_C5Q;
  assign CLBLM_L_X74Y135_SLICE_X113Y135_C4 = CLBLL_R_X75Y133_SLICE_X114Y133_BQ;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_A1 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_A2 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_A3 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_A4 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_A5 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_A6 = 1'b1;
  assign CLBLM_L_X74Y135_SLICE_X113Y135_C5 = CLBLM_L_X74Y134_SLICE_X112Y134_BQ;
  assign CLBLM_L_X74Y135_SLICE_X113Y135_C6 = CLBLM_L_X74Y134_SLICE_X112Y134_CQ;
  assign CLBLM_L_X74Y135_SLICE_X113Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_B1 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_B2 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_B3 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_B4 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_B5 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_B6 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_D4 = 1'b1;
  assign CLBLL_R_X71Y102_SLICE_X107Y102_A1 = 1'b1;
  assign CLBLL_R_X71Y102_SLICE_X107Y102_A2 = 1'b1;
  assign CLBLL_R_X71Y102_SLICE_X107Y102_A3 = 1'b1;
  assign CLBLL_R_X71Y102_SLICE_X107Y102_A4 = 1'b1;
  assign CLBLL_R_X71Y102_SLICE_X107Y102_A5 = 1'b1;
  assign CLBLL_R_X71Y102_SLICE_X107Y102_A6 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_C1 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_C2 = 1'b1;
  assign CLBLL_R_X71Y102_SLICE_X107Y102_B1 = 1'b1;
  assign CLBLL_R_X71Y102_SLICE_X107Y102_B2 = 1'b1;
  assign CLBLL_R_X71Y102_SLICE_X107Y102_B3 = 1'b1;
  assign CLBLL_R_X71Y102_SLICE_X107Y102_B4 = 1'b1;
  assign CLBLL_R_X71Y102_SLICE_X107Y102_B5 = 1'b1;
  assign CLBLL_R_X71Y102_SLICE_X107Y102_B6 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_C5 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_C6 = 1'b1;
  assign CLBLL_R_X71Y102_SLICE_X107Y102_C1 = 1'b1;
  assign CLBLL_R_X71Y102_SLICE_X107Y102_C2 = 1'b1;
  assign CLBLL_R_X71Y102_SLICE_X107Y102_C3 = 1'b1;
  assign CLBLL_R_X71Y102_SLICE_X107Y102_C4 = 1'b1;
  assign CLBLL_R_X71Y102_SLICE_X107Y102_C5 = 1'b1;
  assign CLBLL_R_X71Y102_SLICE_X107Y102_C6 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_D1 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_D2 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_D3 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_D4 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_D5 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_A1 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_A2 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_A3 = 1'b1;
  assign CLBLL_R_X71Y102_SLICE_X107Y102_D1 = 1'b1;
  assign CLBLL_R_X71Y102_SLICE_X107Y102_D2 = 1'b1;
  assign CLBLL_R_X71Y102_SLICE_X107Y102_D3 = 1'b1;
  assign CLBLL_R_X71Y102_SLICE_X107Y102_D4 = 1'b1;
  assign CLBLL_R_X71Y102_SLICE_X107Y102_D5 = 1'b1;
  assign CLBLL_R_X71Y102_SLICE_X107Y102_D6 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_A4 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_A5 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_A6 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_B1 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_B2 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_B3 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_B4 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_C1 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_C2 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_C3 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_C4 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_C5 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_C6 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_C1 = CLBLM_L_X70Y119_SLICE_X105Y119_AQ;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_C2 = CLBLM_L_X70Y123_SLICE_X104Y123_AQ;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_C3 = CLBLL_R_X71Y126_SLICE_X107Y126_BQ;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_C4 = CLBLM_L_X70Y123_SLICE_X104Y123_A5Q;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_C5 = CLBLM_L_X70Y123_SLICE_X104Y123_BQ;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_C6 = CLBLM_L_X70Y125_SLICE_X104Y125_AQ;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_D1 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_D2 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_D3 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_D4 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_D5 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_D6 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_D1 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_D2 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_D3 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_D4 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_D5 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_A1 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_A2 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_A3 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_A4 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_A5 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_A6 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_D3 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_AX = CLBLM_L_X70Y100_SLICE_X105Y100_CQ;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_B1 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_B2 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_B3 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_B4 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_B5 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_B6 = 1'b1;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_D4 = 1'b1;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_D5 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_BX = CLBLM_L_X60Y99_SLICE_X90Y99_DQ;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_D6 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_C1 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_C2 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_C3 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_C4 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_C5 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_C6 = 1'b1;
  assign CLBLM_R_X67Y109_SLICE_X101Y109_D6 = CLBLM_R_X67Y110_SLICE_X101Y110_BQ;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_CX = CLBLM_L_X60Y99_SLICE_X90Y99_BQ;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_D1 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_D2 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_D3 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_D4 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_D5 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_D6 = 1'b1;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X67Y109_SLICE_X100Y109_B5 = CLBLM_R_X67Y108_SLICE_X101Y108_AO6;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_D1 = RIOB33_X105Y51_IOB_X1Y52_I;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_DX = CLBLM_L_X62Y101_SLICE_X92Y101_AQ;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X67Y109_SLICE_X100Y109_B6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_T1 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_D1 = 1'b1;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_A1 = CLBLL_R_X73Y124_SLICE_X110Y124_A5Q;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_D1 = CLBLL_R_X73Y123_SLICE_X110Y123_AQ;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_T1 = 1'b1;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_A3 = CLBLM_L_X72Y124_SLICE_X108Y124_AQ;
  assign LIOB33_X0Y197_IOB_X0Y198_O = 1'b1;
  assign LIOB33_X0Y197_IOB_X0Y197_O = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_T1 = 1'b1;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_A4 = CLBLM_L_X72Y124_SLICE_X108Y124_BO6;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_D1 = CLBLM_L_X70Y111_SLICE_X105Y111_DO6;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_A5 = CLBLM_L_X72Y124_SLICE_X109Y124_AQ;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_A6 = CLBLM_L_X72Y125_SLICE_X108Y125_AQ;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_T1 = 1'b1;
  assign CLBLM_R_X67Y109_SLICE_X100Y109_C5 = CLBLM_R_X67Y108_SLICE_X100Y108_AQ;
  assign CLBLM_R_X67Y109_SLICE_X100Y109_C6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_B1 = CLBLL_R_X71Y126_SLICE_X107Y126_BQ;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_B2 = CLBLM_L_X70Y124_SLICE_X105Y124_BO6;
  assign CLBLM_R_X67Y109_SLICE_X100Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X67Y109_SLICE_X101Y109_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_B3 = CLBLL_R_X71Y126_SLICE_X107Y126_AQ;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_B4 = CLBLM_L_X70Y125_SLICE_X105Y125_AQ;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_B5 = CLBLM_L_X70Y123_SLICE_X104Y123_AQ;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_B6 = CLBLM_L_X70Y124_SLICE_X104Y124_BQ;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_A1 = 1'b1;
  assign CLBLL_R_X71Y103_SLICE_X106Y103_A1 = CLBLM_L_X70Y104_SLICE_X104Y104_A5Q;
  assign CLBLL_R_X71Y103_SLICE_X106Y103_A2 = CLBLM_L_X70Y103_SLICE_X104Y103_DO6;
  assign CLBLL_R_X71Y103_SLICE_X106Y103_A3 = CLBLL_R_X71Y103_SLICE_X106Y103_AQ;
  assign CLBLL_R_X71Y103_SLICE_X106Y103_A4 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLL_R_X71Y103_SLICE_X106Y103_A5 = CLBLM_L_X70Y103_SLICE_X104Y103_B5Q;
  assign CLBLL_R_X71Y103_SLICE_X106Y103_A6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y103_SLICE_X106Y103_B1 = CLBLM_L_X70Y104_SLICE_X104Y104_A5Q;
  assign CLBLL_R_X71Y103_SLICE_X106Y103_B2 = 1'b1;
  assign CLBLL_R_X71Y103_SLICE_X106Y103_B3 = CLBLM_L_X70Y103_SLICE_X104Y103_B5Q;
  assign CLBLL_R_X71Y103_SLICE_X106Y103_B4 = 1'b1;
  assign CLBLL_R_X71Y103_SLICE_X106Y103_B5 = 1'b1;
  assign CLBLL_R_X71Y103_SLICE_X106Y103_B6 = 1'b1;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_C1 = 1'b1;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_C2 = 1'b1;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_A2 = 1'b1;
  assign CLBLL_R_X71Y103_SLICE_X106Y103_C1 = 1'b1;
  assign CLBLL_R_X71Y103_SLICE_X106Y103_C2 = 1'b1;
  assign CLBLL_R_X71Y103_SLICE_X106Y103_C3 = 1'b1;
  assign CLBLL_R_X71Y103_SLICE_X106Y103_C4 = 1'b1;
  assign CLBLL_R_X71Y103_SLICE_X106Y103_C5 = 1'b1;
  assign CLBLL_R_X71Y103_SLICE_X106Y103_C6 = 1'b1;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_C3 = 1'b1;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_C4 = 1'b1;
  assign CLBLL_R_X71Y103_SLICE_X106Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_C5 = 1'b1;
  assign CLBLL_R_X71Y103_SLICE_X106Y103_D1 = 1'b1;
  assign CLBLL_R_X71Y103_SLICE_X106Y103_D2 = 1'b1;
  assign CLBLL_R_X71Y103_SLICE_X106Y103_D3 = 1'b1;
  assign CLBLL_R_X71Y103_SLICE_X106Y103_D4 = 1'b1;
  assign CLBLL_R_X71Y103_SLICE_X106Y103_D5 = 1'b1;
  assign CLBLL_R_X71Y103_SLICE_X106Y103_D6 = 1'b1;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_C6 = 1'b1;
  assign CLBLL_R_X71Y103_SLICE_X106Y103_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_A3 = CLBLM_R_X63Y102_SLICE_X95Y102_AQ;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_A1 = CLBLM_L_X70Y123_SLICE_X104Y123_AQ;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_A2 = CLBLL_R_X71Y126_SLICE_X107Y126_BQ;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_A3 = CLBLL_R_X71Y126_SLICE_X107Y126_AQ;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_A4 = CLBLM_L_X70Y124_SLICE_X105Y124_BO6;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_A5 = CLBLM_L_X70Y125_SLICE_X105Y125_AQ;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_A6 = CLBLM_L_X70Y125_SLICE_X104Y125_BQ;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_B1 = CLBLM_L_X70Y123_SLICE_X104Y123_AQ;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_B2 = CLBLM_L_X70Y123_SLICE_X104Y123_BQ;
  assign CLBLL_R_X71Y103_SLICE_X107Y103_A1 = 1'b1;
  assign CLBLL_R_X71Y103_SLICE_X107Y103_A2 = 1'b1;
  assign CLBLL_R_X71Y103_SLICE_X107Y103_A3 = 1'b1;
  assign CLBLL_R_X71Y103_SLICE_X107Y103_A4 = 1'b1;
  assign CLBLL_R_X71Y103_SLICE_X107Y103_A5 = 1'b1;
  assign CLBLL_R_X71Y103_SLICE_X107Y103_A6 = 1'b1;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_B3 = CLBLM_L_X70Y119_SLICE_X105Y119_AQ;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_B4 = CLBLL_R_X71Y126_SLICE_X107Y126_BQ;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_B5 = CLBLM_L_X70Y125_SLICE_X104Y125_AQ;
  assign CLBLL_R_X71Y103_SLICE_X107Y103_B1 = 1'b1;
  assign CLBLL_R_X71Y103_SLICE_X107Y103_B2 = 1'b1;
  assign CLBLL_R_X71Y103_SLICE_X107Y103_B3 = 1'b1;
  assign CLBLL_R_X71Y103_SLICE_X107Y103_B4 = 1'b1;
  assign CLBLL_R_X71Y103_SLICE_X107Y103_B5 = 1'b1;
  assign CLBLL_R_X71Y103_SLICE_X107Y103_B6 = 1'b1;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_C1 = CLBLM_L_X70Y119_SLICE_X105Y119_AQ;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_C2 = CLBLM_L_X70Y125_SLICE_X104Y125_AQ;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_C3 = CLBLM_L_X70Y123_SLICE_X104Y123_BQ;
  assign CLBLL_R_X71Y103_SLICE_X107Y103_C1 = 1'b1;
  assign CLBLL_R_X71Y103_SLICE_X107Y103_C2 = 1'b1;
  assign CLBLL_R_X71Y103_SLICE_X107Y103_C3 = 1'b1;
  assign CLBLL_R_X71Y103_SLICE_X107Y103_C4 = 1'b1;
  assign CLBLL_R_X71Y103_SLICE_X107Y103_C5 = 1'b1;
  assign CLBLL_R_X71Y103_SLICE_X107Y103_C6 = 1'b1;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_D1 = CLBLM_L_X70Y119_SLICE_X105Y119_AQ;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_D2 = CLBLM_L_X70Y125_SLICE_X104Y125_AQ;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_D3 = CLBLM_L_X70Y123_SLICE_X104Y123_BQ;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_D4 = CLBLM_L_X70Y123_SLICE_X104Y123_A5Q;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_D5 = CLBLM_L_X70Y123_SLICE_X104Y123_AQ;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_D6 = CLBLL_R_X71Y126_SLICE_X107Y126_BQ;
  assign CLBLL_R_X71Y103_SLICE_X107Y103_D1 = 1'b1;
  assign CLBLL_R_X71Y103_SLICE_X107Y103_D2 = 1'b1;
  assign CLBLL_R_X71Y103_SLICE_X107Y103_D3 = 1'b1;
  assign CLBLL_R_X71Y103_SLICE_X107Y103_D4 = 1'b1;
  assign CLBLL_R_X71Y103_SLICE_X107Y103_D5 = 1'b1;
  assign CLBLL_R_X71Y103_SLICE_X107Y103_D6 = 1'b1;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_A1 = CLBLM_L_X70Y125_SLICE_X105Y125_AO5;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_A2 = CLBLM_L_X70Y125_SLICE_X105Y125_BO6;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_A3 = CLBLM_L_X70Y124_SLICE_X104Y124_AQ;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_A4 = CLBLL_R_X71Y124_SLICE_X106Y124_AQ;
  assign CLBLL_R_X79Y99_SLICE_X122Y99_A1 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X122Y99_A2 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X122Y99_A3 = CLBLM_R_X103Y69_SLICE_X162Y69_A5Q;
  assign CLBLL_R_X79Y99_SLICE_X122Y99_A4 = CLBLM_L_X82Y98_SLICE_X128Y98_A5Q;
  assign CLBLL_R_X79Y99_SLICE_X122Y99_A5 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X122Y99_A6 = 1'b1;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_B1 = CLBLM_L_X70Y123_SLICE_X104Y123_CO6;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_B2 = CLBLM_L_X70Y124_SLICE_X104Y124_BQ;
  assign CLBLL_R_X79Y99_SLICE_X122Y99_B1 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X122Y99_B2 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X122Y99_B3 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X122Y99_B4 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X122Y99_B5 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X122Y99_B6 = 1'b1;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_C2 = CLBLM_L_X70Y124_SLICE_X104Y124_CQ;
  assign CLBLL_R_X79Y99_SLICE_X122Y99_C1 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X122Y99_C2 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X122Y99_C3 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X122Y99_C4 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X122Y99_C5 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X122Y99_C6 = 1'b1;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_C6 = CLBLM_L_X70Y125_SLICE_X105Y125_BO6;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_D1 = CLBLM_L_X70Y119_SLICE_X105Y119_AQ;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_D2 = CLBLM_L_X70Y123_SLICE_X104Y123_A5Q;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_D3 = CLBLM_L_X70Y123_SLICE_X104Y123_AQ;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_D4 = CLBLM_L_X70Y125_SLICE_X104Y125_AQ;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_D5 = CLBLM_L_X70Y123_SLICE_X104Y123_BQ;
  assign CLBLL_R_X79Y99_SLICE_X122Y99_D1 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X122Y99_D2 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X122Y99_D3 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X122Y99_D4 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X122Y99_D5 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X122Y99_D6 = 1'b1;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_D6 = CLBLL_R_X71Y126_SLICE_X107Y126_BQ;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X76Y134_SLICE_X117Y134_D3 = 1'b1;
  assign CLBLM_R_X67Y109_SLICE_X100Y109_A5 = CLBLM_R_X67Y108_SLICE_X101Y108_AO6;
  assign CLBLM_L_X76Y134_SLICE_X117Y134_D4 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X123Y99_A1 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X123Y99_A2 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X123Y99_A3 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X123Y99_A4 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X123Y99_A5 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X123Y99_A6 = 1'b1;
  assign CLBLM_R_X67Y109_SLICE_X100Y109_A6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X79Y99_SLICE_X123Y99_B1 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X123Y99_B2 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X123Y99_B3 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X123Y99_B4 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X123Y99_B5 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X123Y99_B6 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X123Y99_C1 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X123Y99_C2 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X123Y99_C3 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X123Y99_C4 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X123Y99_C5 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X123Y99_C6 = 1'b1;
  assign CLBLM_L_X76Y134_SLICE_X117Y134_D5 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X123Y99_D1 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X123Y99_D2 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X123Y99_D3 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X123Y99_D4 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X123Y99_D5 = 1'b1;
  assign CLBLL_R_X79Y99_SLICE_X123Y99_D6 = 1'b1;
  assign CLBLM_L_X76Y134_SLICE_X117Y134_D6 = 1'b1;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_D4 = 1'b1;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_D5 = 1'b1;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_D6 = 1'b1;
  assign CLBLM_L_X76Y134_SLICE_X117Y134_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign RIOI3_X105Y75_OLOGIC_X1Y76_D1 = CLBLM_R_X103Y75_SLICE_X163Y75_BQ;
  assign CLBLM_L_X70Y125_SLICE_X105Y125_A1 = 1'b1;
  assign CLBLM_L_X70Y125_SLICE_X105Y125_A2 = CLBLM_L_X70Y123_SLICE_X104Y123_A5Q;
  assign CLBLM_L_X70Y125_SLICE_X105Y125_A3 = CLBLM_L_X70Y119_SLICE_X105Y119_AQ;
  assign CLBLM_L_X70Y125_SLICE_X105Y125_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y125_SLICE_X105Y125_A5 = CLBLM_L_X70Y125_SLICE_X104Y125_AQ;
  assign CLBLM_L_X70Y125_SLICE_X105Y125_A6 = 1'b1;
  assign CLBLM_L_X70Y125_SLICE_X105Y125_AX = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y125_SLICE_X105Y125_B1 = 1'b1;
  assign CLBLM_L_X70Y125_SLICE_X105Y125_B2 = CLBLM_L_X70Y123_SLICE_X104Y123_BQ;
  assign CLBLM_L_X70Y125_SLICE_X105Y125_B3 = CLBLM_L_X70Y119_SLICE_X105Y119_AQ;
  assign CLBLM_L_X70Y125_SLICE_X105Y125_B4 = CLBLM_L_X70Y123_SLICE_X104Y123_A5Q;
  assign CLBLM_L_X70Y125_SLICE_X105Y125_B5 = CLBLM_L_X70Y125_SLICE_X104Y125_AQ;
  assign CLBLM_L_X70Y125_SLICE_X105Y125_B6 = 1'b1;
  assign CLBLM_L_X70Y125_SLICE_X105Y125_BX = CLBLM_L_X70Y125_SLICE_X105Y125_AO6;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_B3 = CLBLM_L_X76Y125_SLICE_X116Y125_C5Q;
  assign CLBLM_L_X70Y125_SLICE_X105Y125_C1 = CLBLM_L_X70Y125_SLICE_X105Y125_AQ;
  assign CLBLM_L_X70Y125_SLICE_X105Y125_C2 = CLBLL_R_X71Y126_SLICE_X107Y126_AQ;
  assign CLBLM_L_X70Y125_SLICE_X105Y125_C3 = CLBLM_L_X70Y126_SLICE_X105Y126_DO6;
  assign CLBLM_L_X70Y125_SLICE_X105Y125_C4 = CLBLM_L_X70Y125_SLICE_X104Y125_CQ;
  assign CLBLM_L_X70Y125_SLICE_X105Y125_C5 = CLBLM_L_X70Y125_SLICE_X105Y125_DO6;
  assign CLBLM_L_X70Y125_SLICE_X105Y125_C6 = CLBLM_L_X70Y125_SLICE_X104Y125_BQ;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_B4 = CLBLM_L_X76Y122_SLICE_X116Y122_CQ;
  assign RIOB33_X105Y147_IOB_X1Y147_O = CLBLL_R_X77Y108_SLICE_X118Y108_AQ;
  assign CLBLM_L_X70Y125_SLICE_X105Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_B5 = CLBLM_L_X72Y118_SLICE_X108Y118_CQ;
  assign CLBLM_L_X70Y109_SLICE_X105Y109_C1 = 1'b1;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_B6 = 1'b1;
  assign CLBLM_L_X70Y125_SLICE_X105Y125_D1 = CLBLM_L_X70Y124_SLICE_X105Y124_DO6;
  assign CLBLM_L_X70Y109_SLICE_X105Y109_C2 = 1'b1;
  assign CLBLM_L_X70Y125_SLICE_X105Y125_D2 = CLBLL_R_X71Y126_SLICE_X107Y126_AQ;
  assign CLBLM_L_X70Y125_SLICE_X105Y125_D4 = 1'b1;
  assign CLBLM_L_X70Y125_SLICE_X105Y125_D5 = CLBLM_L_X70Y125_SLICE_X105Y125_AQ;
  assign CLBLM_L_X70Y125_SLICE_X105Y125_D6 = CLBLL_R_X71Y125_SLICE_X106Y125_AQ;
  assign CLBLM_L_X70Y109_SLICE_X105Y109_C3 = 1'b1;
  assign CLBLM_L_X70Y125_SLICE_X105Y125_D3 = CLBLL_R_X71Y125_SLICE_X107Y125_AQ;
  assign CLBLM_L_X70Y125_SLICE_X105Y125_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X70Y109_SLICE_X105Y109_C4 = 1'b1;
  assign CLBLM_L_X70Y125_SLICE_X104Y125_A1 = 1'b1;
  assign CLBLM_L_X70Y125_SLICE_X104Y125_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_A1 = 1'b1;
  assign CLBLM_L_X70Y125_SLICE_X104Y125_A4 = CLBLM_L_X70Y125_SLICE_X105Y125_BQ;
  assign CLBLM_L_X70Y125_SLICE_X104Y125_A5 = CLBLM_L_X70Y123_SLICE_X104Y123_BQ;
  assign CLBLM_L_X70Y125_SLICE_X104Y125_A6 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_A2 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_A3 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_A4 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_A5 = 1'b1;
  assign CLBLM_L_X70Y125_SLICE_X104Y125_B1 = CLBLM_L_X70Y125_SLICE_X104Y125_CQ;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_A6 = 1'b1;
  assign CLBLM_L_X70Y125_SLICE_X104Y125_B3 = 1'b1;
  assign CLBLM_L_X70Y125_SLICE_X104Y125_B4 = CLBLM_L_X70Y123_SLICE_X104Y123_CO6;
  assign CLBLM_L_X70Y125_SLICE_X104Y125_B5 = CLBLM_L_X70Y126_SLICE_X104Y126_AQ;
  assign CLBLM_L_X70Y125_SLICE_X104Y125_B6 = CLBLM_L_X70Y125_SLICE_X104Y125_BQ;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_B1 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_B2 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_B3 = 1'b1;
  assign CLBLM_L_X70Y125_SLICE_X104Y125_C1 = 1'b1;
  assign CLBLM_L_X70Y125_SLICE_X104Y125_C2 = CLBLM_L_X70Y125_SLICE_X104Y125_CQ;
  assign CLBLM_L_X70Y125_SLICE_X104Y125_C3 = CLBLM_L_X70Y124_SLICE_X104Y124_DO6;
  assign CLBLM_L_X70Y125_SLICE_X104Y125_C4 = CLBLM_L_X70Y126_SLICE_X104Y126_BQ;
  assign CLBLM_L_X70Y125_SLICE_X104Y125_C5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y125_SLICE_X104Y125_C6 = CLBLL_R_X71Y125_SLICE_X106Y125_AQ;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_C4 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_C1 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_C2 = 1'b1;
  assign CLBLM_L_X70Y125_SLICE_X104Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_C5 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_C6 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_D1 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_D2 = 1'b1;
  assign CLBLM_L_X70Y125_SLICE_X104Y125_D1 = CLBLL_R_X71Y126_SLICE_X107Y126_BQ;
  assign CLBLM_L_X70Y125_SLICE_X104Y125_D2 = CLBLM_L_X70Y125_SLICE_X104Y125_CQ;
  assign CLBLM_L_X70Y125_SLICE_X104Y125_D3 = CLBLM_L_X70Y123_SLICE_X104Y123_AQ;
  assign CLBLM_L_X70Y125_SLICE_X104Y125_D4 = CLBLM_L_X70Y125_SLICE_X104Y125_BQ;
  assign CLBLM_L_X70Y125_SLICE_X104Y125_D5 = CLBLL_R_X71Y125_SLICE_X107Y125_AQ;
  assign CLBLM_L_X70Y125_SLICE_X104Y125_D6 = CLBLL_R_X71Y125_SLICE_X106Y125_AQ;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_D3 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_D4 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_D5 = 1'b1;
  assign CLBLM_L_X70Y125_SLICE_X104Y125_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_A1 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_A2 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_A3 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_A4 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_A5 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_A6 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_AX = CLBLM_L_X62Y95_SLICE_X92Y95_AQ;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_B1 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_B2 = 1'b1;
  assign CLBLM_L_X70Y109_SLICE_X105Y109_D1 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_B3 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_B5 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_B6 = 1'b1;
  assign CLBLM_L_X70Y109_SLICE_X105Y109_D2 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_B4 = 1'b1;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_BX = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_L_X70Y109_SLICE_X105Y109_D3 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_C1 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_C2 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_C3 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_C4 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_C5 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_C6 = 1'b1;
  assign CLBLM_L_X70Y109_SLICE_X105Y109_D4 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X70Y109_SLICE_X105Y109_D5 = 1'b1;
  assign CLBLM_L_X70Y109_SLICE_X105Y109_D6 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_D1 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_D2 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_D3 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_D4 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_D5 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_D6 = 1'b1;
  assign RIOI3_X105Y77_OLOGIC_X1Y77_D1 = CLBLM_R_X103Y76_SLICE_X163Y76_AQ;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_T1 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X70Y109_SLICE_X105Y109_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_D4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_D5 = CLBLM_L_X74Y119_SLICE_X112Y119_BO5;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_A5 = 1'b1;
  assign CLBLM_L_X70Y109_SLICE_X104Y109_A1 = CLBLM_L_X70Y112_SLICE_X105Y112_B5Q;
  assign CLBLM_L_X70Y109_SLICE_X104Y109_A2 = CLBLM_L_X70Y109_SLICE_X104Y109_BQ;
  assign CLBLM_L_X70Y109_SLICE_X104Y109_A3 = CLBLM_L_X70Y113_SLICE_X104Y113_B5Q;
  assign CLBLM_L_X70Y109_SLICE_X104Y109_A4 = CLBLM_L_X70Y107_SLICE_X104Y107_BQ;
  assign CLBLM_L_X70Y109_SLICE_X104Y109_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y109_SLICE_X104Y109_A6 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_D1 = 1'b1;
  assign CLBLM_L_X76Y126_SLICE_X117Y126_C3 = 1'b1;
  assign CLBLM_L_X76Y126_SLICE_X117Y126_C6 = 1'b1;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_B6 = 1'b1;
  assign CLBLM_L_X70Y109_SLICE_X104Y109_B1 = CLBLM_L_X70Y112_SLICE_X105Y112_B5Q;
  assign CLBLM_L_X70Y109_SLICE_X104Y109_B2 = CLBLM_L_X70Y109_SLICE_X104Y109_A5Q;
  assign CLBLM_L_X70Y109_SLICE_X104Y109_B3 = CLBLM_L_X70Y109_SLICE_X104Y109_AQ;
  assign CLBLM_L_X70Y109_SLICE_X104Y109_B5 = CLBLM_R_X65Y106_SLICE_X99Y106_AQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_D1 = CLBLL_L_X34Y123_SLICE_X50Y123_AO6;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_C1 = 1'b1;
  assign CLBLM_L_X70Y109_SLICE_X104Y109_B6 = 1'b1;
  assign CLBLM_L_X78Y104_SLICE_X121Y104_A1 = 1'b1;
  assign CLBLM_L_X78Y104_SLICE_X121Y104_A2 = 1'b1;
  assign CLBLM_L_X78Y104_SLICE_X121Y104_A3 = 1'b1;
  assign CLBLM_L_X78Y104_SLICE_X121Y104_A5 = 1'b1;
  assign CLBLM_L_X78Y104_SLICE_X121Y104_A6 = 1'b1;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_C4 = 1'b1;
  assign CLBLM_L_X78Y104_SLICE_X121Y104_A4 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_T1 = 1'b1;
  assign CLBLM_L_X78Y104_SLICE_X121Y104_B1 = 1'b1;
  assign CLBLM_L_X78Y104_SLICE_X121Y104_B2 = 1'b1;
  assign CLBLM_L_X76Y126_SLICE_X117Y126_D1 = 1'b1;
  assign CLBLM_L_X78Y104_SLICE_X121Y104_B3 = 1'b1;
  assign CLBLM_L_X78Y104_SLICE_X121Y104_B4 = 1'b1;
  assign CLBLM_L_X78Y104_SLICE_X121Y104_B5 = 1'b1;
  assign CLBLM_L_X76Y126_SLICE_X117Y126_D2 = 1'b1;
  assign CLBLM_L_X78Y104_SLICE_X121Y104_B6 = 1'b1;
  assign CLBLM_L_X78Y104_SLICE_X121Y104_C1 = 1'b1;
  assign CLBLM_L_X78Y104_SLICE_X121Y104_C2 = 1'b1;
  assign CLBLM_L_X76Y126_SLICE_X117Y126_D3 = 1'b1;
  assign CLBLM_L_X78Y104_SLICE_X121Y104_C3 = 1'b1;
  assign CLBLM_L_X78Y104_SLICE_X121Y104_C4 = 1'b1;
  assign CLBLM_L_X78Y104_SLICE_X121Y104_C5 = 1'b1;
  assign CLBLM_L_X78Y104_SLICE_X121Y104_C6 = 1'b1;
  assign CLBLM_L_X76Y126_SLICE_X117Y126_D4 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_T1 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_D1 = 1'b1;
  assign CLBLM_L_X76Y126_SLICE_X117Y126_D5 = 1'b1;
  assign CLBLM_L_X78Y104_SLICE_X121Y104_D1 = 1'b1;
  assign CLBLM_L_X78Y104_SLICE_X121Y104_D2 = 1'b1;
  assign CLBLM_L_X76Y126_SLICE_X117Y126_D6 = 1'b1;
  assign CLBLM_L_X78Y104_SLICE_X121Y104_D3 = 1'b1;
  assign CLBLM_L_X78Y104_SLICE_X121Y104_D4 = 1'b1;
  assign CLBLM_L_X78Y104_SLICE_X121Y104_D5 = 1'b1;
  assign CLBLM_L_X78Y104_SLICE_X121Y104_D6 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_T1 = 1'b1;
  assign CLBLM_L_X70Y109_SLICE_X104Y109_C5 = 1'b1;
  assign CLBLM_L_X78Y104_SLICE_X120Y104_A1 = CLBLM_L_X74Y121_SLICE_X113Y121_B5Q;
  assign CLBLM_L_X70Y109_SLICE_X104Y109_C6 = 1'b1;
  assign CLBLM_L_X78Y104_SLICE_X120Y104_A2 = CLBLM_L_X78Y104_SLICE_X120Y104_BQ;
  assign CLBLM_L_X78Y104_SLICE_X120Y104_A3 = CLBLM_L_X78Y104_SLICE_X120Y104_AQ;
  assign CLBLM_L_X78Y104_SLICE_X120Y104_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X78Y104_SLICE_X120Y104_A5 = CLBLM_L_X78Y104_SLICE_X120Y104_A5Q;
  assign CLBLM_L_X78Y104_SLICE_X120Y104_A6 = 1'b1;
  assign CLBLM_L_X70Y126_SLICE_X105Y126_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y126_SLICE_X105Y126_A2 = CLBLM_L_X70Y126_SLICE_X105Y126_BQ;
  assign CLBLM_L_X70Y126_SLICE_X105Y126_A3 = CLBLM_L_X70Y126_SLICE_X105Y126_AQ;
  assign CLBLM_L_X70Y126_SLICE_X105Y126_A4 = CLBLL_R_X71Y126_SLICE_X106Y126_AQ;
  assign CLBLM_L_X70Y126_SLICE_X105Y126_A5 = 1'b1;
  assign CLBLM_L_X70Y126_SLICE_X105Y126_A6 = CLBLM_L_X70Y124_SLICE_X105Y124_CO6;
  assign CLBLM_L_X76Y126_SLICE_X117Y126_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X78Y104_SLICE_X120Y104_B1 = 1'b1;
  assign CLBLM_L_X70Y126_SLICE_X105Y126_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y126_SLICE_X105Y126_B2 = CLBLM_L_X70Y126_SLICE_X105Y126_BQ;
  assign CLBLM_L_X70Y126_SLICE_X105Y126_B3 = CLBLM_L_X70Y125_SLICE_X105Y125_BO6;
  assign CLBLM_L_X70Y109_SLICE_X104Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X70Y126_SLICE_X105Y126_B4 = CLBLL_R_X73Y126_SLICE_X110Y126_BQ;
  assign CLBLM_L_X70Y126_SLICE_X105Y126_B5 = CLBLM_L_X70Y125_SLICE_X105Y125_AO5;
  assign CLBLM_L_X70Y126_SLICE_X105Y126_B6 = CLBLM_L_X70Y124_SLICE_X104Y124_CQ;
  assign CLBLM_L_X78Y104_SLICE_X120Y104_B6 = 1'b1;
  assign CLBLM_L_X78Y104_SLICE_X120Y104_BX = CLBLM_L_X78Y104_SLICE_X120Y104_A5Q;
  assign CLBLM_L_X70Y126_SLICE_X105Y126_C1 = CLBLM_L_X70Y125_SLICE_X104Y125_CQ;
  assign CLBLM_L_X70Y126_SLICE_X105Y126_C2 = CLBLM_L_X70Y123_SLICE_X104Y123_AQ;
  assign CLBLM_L_X70Y126_SLICE_X105Y126_C3 = CLBLL_R_X71Y126_SLICE_X107Y126_AQ;
  assign CLBLM_L_X70Y126_SLICE_X105Y126_C4 = CLBLL_R_X71Y126_SLICE_X107Y126_BQ;
  assign CLBLM_L_X70Y126_SLICE_X105Y126_C5 = CLBLM_L_X70Y125_SLICE_X105Y125_AQ;
  assign CLBLM_L_X70Y126_SLICE_X105Y126_C6 = CLBLM_L_X70Y124_SLICE_X105Y124_BO6;
  assign CLBLM_L_X76Y126_SLICE_X116Y126_A1 = CLBLM_L_X76Y126_SLICE_X116Y126_B5Q;
  assign CLBLM_L_X76Y126_SLICE_X116Y126_A2 = CLBLM_L_X76Y126_SLICE_X116Y126_DQ;
  assign CLBLM_L_X70Y126_SLICE_X105Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X78Y104_SLICE_X120Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X78Y104_SLICE_X120Y104_D1 = 1'b1;
  assign CLBLM_L_X76Y126_SLICE_X116Y126_A3 = CLBLM_L_X76Y125_SLICE_X116Y125_CQ;
  assign CLBLM_L_X78Y104_SLICE_X120Y104_D2 = 1'b1;
  assign CLBLM_L_X70Y126_SLICE_X105Y126_D1 = CLBLL_R_X71Y126_SLICE_X107Y126_AQ;
  assign CLBLM_L_X70Y126_SLICE_X105Y126_D2 = CLBLM_L_X70Y128_SLICE_X104Y128_CQ;
  assign CLBLM_L_X70Y126_SLICE_X105Y126_D3 = CLBLM_L_X70Y125_SLICE_X105Y125_AQ;
  assign CLBLM_L_X70Y126_SLICE_X105Y126_D4 = CLBLL_R_X71Y126_SLICE_X107Y126_AO5;
  assign CLBLM_L_X70Y126_SLICE_X105Y126_D5 = CLBLM_L_X70Y124_SLICE_X105Y124_DO6;
  assign CLBLM_L_X70Y126_SLICE_X105Y126_D6 = CLBLM_L_X70Y133_SLICE_X105Y133_BQ;
  assign CLBLM_L_X76Y126_SLICE_X116Y126_A4 = CLBLM_L_X76Y126_SLICE_X116Y126_CQ;
  assign CLBLM_L_X76Y126_SLICE_X116Y126_A5 = CLBLM_L_X76Y126_SLICE_X116Y126_BQ;
  assign CLBLM_L_X70Y126_SLICE_X105Y126_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X78Y104_SLICE_X120Y104_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X76Y126_SLICE_X116Y126_A6 = 1'b1;
  assign CLBLM_L_X70Y126_SLICE_X104Y126_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y126_SLICE_X104Y126_A2 = CLBLM_L_X70Y125_SLICE_X105Y125_AO5;
  assign CLBLM_L_X70Y126_SLICE_X104Y126_A3 = CLBLM_L_X70Y126_SLICE_X104Y126_AQ;
  assign CLBLM_L_X70Y126_SLICE_X104Y126_A4 = CLBLM_L_X70Y133_SLICE_X104Y133_BQ;
  assign CLBLM_L_X70Y126_SLICE_X104Y126_A5 = CLBLM_L_X70Y125_SLICE_X105Y125_BO6;
  assign CLBLM_L_X70Y126_SLICE_X104Y126_A6 = CLBLM_L_X70Y125_SLICE_X104Y125_A5Q;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_D1 = 1'b1;
  assign CLBLM_L_X70Y126_SLICE_X104Y126_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y126_SLICE_X104Y126_B2 = CLBLM_L_X70Y126_SLICE_X104Y126_BQ;
  assign CLBLM_L_X70Y126_SLICE_X104Y126_B3 = CLBLM_L_X70Y125_SLICE_X105Y125_AO5;
  assign CLBLM_L_X70Y126_SLICE_X104Y126_B4 = CLBLM_L_X70Y126_SLICE_X104Y126_AQ;
  assign CLBLM_L_X70Y126_SLICE_X104Y126_B5 = CLBLM_L_X70Y125_SLICE_X105Y125_BO6;
  assign CLBLM_L_X70Y109_SLICE_X104Y109_D4 = 1'b1;
  assign CLBLM_L_X70Y126_SLICE_X104Y126_B6 = CLBLM_L_X70Y129_SLICE_X104Y129_BQ;
  assign CLBLM_L_X70Y109_SLICE_X104Y109_D5 = 1'b1;
  assign CLBLM_L_X70Y126_SLICE_X104Y126_C1 = CLBLM_L_X70Y126_SLICE_X105Y126_AQ;
  assign CLBLM_L_X70Y126_SLICE_X104Y126_C2 = CLBLM_L_X70Y126_SLICE_X104Y126_CQ;
  assign CLBLM_L_X70Y126_SLICE_X104Y126_C3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y126_SLICE_X104Y126_C4 = CLBLM_L_X70Y124_SLICE_X104Y124_CQ;
  assign CLBLM_L_X70Y126_SLICE_X104Y126_C5 = CLBLM_L_X70Y124_SLICE_X104Y124_DO6;
  assign CLBLM_L_X70Y126_SLICE_X104Y126_C6 = 1'b1;
  assign CLBLM_L_X76Y126_SLICE_X116Y126_B1 = CLBLM_L_X76Y126_SLICE_X116Y126_B5Q;
  assign CLBLM_L_X70Y126_SLICE_X104Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X76Y126_SLICE_X116Y126_B2 = CLBLM_L_X76Y126_SLICE_X116Y126_BQ;
  assign CLBLM_L_X70Y126_SLICE_X104Y126_D1 = CLBLM_L_X70Y126_SLICE_X105Y126_AQ;
  assign CLBLM_L_X70Y126_SLICE_X104Y126_D2 = CLBLM_L_X70Y126_SLICE_X104Y126_CQ;
  assign CLBLM_L_X70Y126_SLICE_X104Y126_D3 = CLBLM_L_X70Y124_SLICE_X104Y124_BQ;
  assign CLBLM_L_X70Y126_SLICE_X104Y126_D4 = CLBLM_L_X70Y123_SLICE_X104Y123_AQ;
  assign CLBLM_L_X70Y126_SLICE_X104Y126_D5 = CLBLL_R_X71Y126_SLICE_X106Y126_AQ;
  assign CLBLM_L_X70Y126_SLICE_X104Y126_D6 = CLBLL_R_X71Y126_SLICE_X107Y126_BQ;
  assign CLBLM_L_X76Y126_SLICE_X116Y126_B3 = CLBLM_L_X76Y125_SLICE_X116Y125_CQ;
  assign CLBLM_L_X76Y126_SLICE_X116Y126_B4 = CLBLL_R_X77Y127_SLICE_X119Y127_AO5;
  assign CLBLM_L_X70Y126_SLICE_X104Y126_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X76Y126_SLICE_X116Y126_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X76Y126_SLICE_X116Y126_B6 = 1'b1;
  assign CLBLM_L_X76Y126_SLICE_X116Y126_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X76Y126_SLICE_X116Y126_C2 = CLBLM_L_X76Y125_SLICE_X116Y125_CQ;
  assign CLBLM_L_X76Y126_SLICE_X116Y126_C3 = CLBLM_L_X76Y126_SLICE_X116Y126_BQ;
  assign CLBLM_L_X78Y128_SLICE_X120Y128_A6 = 1'b1;
  assign CLBLM_L_X76Y126_SLICE_X116Y126_C4 = CLBLL_R_X77Y127_SLICE_X119Y127_AO5;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_B1 = 1'b1;
  assign CLBLM_L_X76Y126_SLICE_X116Y126_C5 = CLBLM_L_X76Y126_SLICE_X116Y126_B5Q;
  assign CLBLM_L_X76Y126_SLICE_X116Y126_C6 = CLBLM_L_X76Y126_SLICE_X116Y126_CQ;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_B4 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_B6 = 1'b1;
  assign CLBLM_L_X76Y126_SLICE_X116Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X83Y130_SLICE_X130Y130_A1 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X130Y130_A2 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X130Y130_A3 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X130Y130_A4 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X130Y130_A5 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X130Y130_A6 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_C1 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_C2 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X130Y130_AX = CLBLL_R_X83Y132_SLICE_X130Y132_AQ;
  assign CLBLM_L_X72Y130_SLICE_X108Y130_D6 = CLBLL_R_X71Y129_SLICE_X106Y129_AQ;
  assign CLBLL_R_X83Y130_SLICE_X130Y130_B1 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X130Y130_B2 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X130Y130_B3 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X130Y130_B4 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X130Y130_B5 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X130Y130_B6 = 1'b1;
  assign CLBLM_L_X76Y126_SLICE_X116Y126_D1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X83Y130_SLICE_X130Y130_BX = CLBLL_R_X83Y130_SLICE_X130Y130_AQ;
  assign CLBLL_R_X83Y130_SLICE_X130Y130_C1 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X130Y130_C2 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X130Y130_C3 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X130Y130_C4 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X130Y130_C5 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X130Y130_C6 = 1'b1;
  assign CLBLM_L_X76Y126_SLICE_X116Y126_D2 = CLBLM_L_X76Y126_SLICE_X116Y126_CQ;
  assign CLBLM_L_X76Y126_SLICE_X116Y126_D3 = CLBLM_L_X76Y126_SLICE_X116Y126_DQ;
  assign CLBLL_R_X83Y130_SLICE_X130Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X76Y126_SLICE_X116Y126_D4 = CLBLM_L_X76Y126_SLICE_X116Y126_AO5;
  assign CLBLL_R_X83Y130_SLICE_X130Y130_CX = CLBLL_R_X83Y130_SLICE_X130Y130_BQ;
  assign CLBLL_R_X83Y130_SLICE_X130Y130_D1 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X130Y130_D2 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X130Y130_D3 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X130Y130_D4 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X130Y130_D5 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X130Y130_D6 = 1'b1;
  assign CLBLM_L_X76Y126_SLICE_X116Y126_D5 = CLBLM_L_X76Y126_SLICE_X116Y126_B5Q;
  assign CLBLM_L_X76Y126_SLICE_X116Y126_D6 = CLBLL_R_X77Y127_SLICE_X119Y127_AO5;
  assign CLBLL_R_X83Y130_SLICE_X130Y130_DX = CLBLL_R_X83Y130_SLICE_X130Y130_CQ;
  assign CLBLL_R_X83Y130_SLICE_X130Y130_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y133_SLICE_X112Y133_D5 = 1'b1;
  assign CLBLM_L_X76Y126_SLICE_X116Y126_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X83Y130_SLICE_X131Y130_A1 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X131Y130_A2 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X131Y130_A3 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X131Y130_A4 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X131Y130_A5 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X131Y130_A6 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X131Y130_B1 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X131Y130_B2 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X131Y130_B3 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X131Y130_B4 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X131Y130_B5 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X131Y130_B6 = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_D1 = CLBLM_L_X62Y107_SLICE_X92Y107_AO5;
  assign CLBLL_R_X83Y130_SLICE_X131Y130_C1 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X131Y130_C2 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X131Y130_C3 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X131Y130_C4 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X131Y130_C5 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X131Y130_C6 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_D4 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X131Y130_D1 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X131Y130_D2 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X131Y130_D3 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X131Y130_D4 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X131Y130_D5 = 1'b1;
  assign CLBLL_R_X83Y130_SLICE_X131Y130_D6 = 1'b1;
  assign CLBLM_L_X70Y109_SLICE_X105Y109_C5 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X120Y128_B2 = 1'b1;
  assign CLBLM_L_X70Y109_SLICE_X105Y109_C6 = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_D1 = CLBLM_R_X67Y118_SLICE_X100Y118_A5Q;
  assign CLBLM_L_X74Y133_SLICE_X112Y133_D6 = 1'b1;
  assign CLBLM_L_X82Y130_SLICE_X129Y130_B5 = 1'b1;
  assign CLBLM_L_X70Y109_SLICE_X105Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X67Y109_SLICE_X100Y109_D4 = CLBLM_L_X60Y97_SLICE_X91Y97_AQ;
  assign CLBLM_R_X67Y109_SLICE_X100Y109_D5 = CLBLM_R_X65Y110_SLICE_X99Y110_B5Q;
  assign CLBLM_R_X67Y105_SLICE_X100Y105_A2 = CLBLM_L_X68Y103_SLICE_X102Y103_B5Q;
  assign CLBLM_R_X67Y110_SLICE_X101Y110_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y110_SLICE_X101Y110_A5 = CLBLM_R_X67Y109_SLICE_X101Y109_AQ;
  assign CLBLM_R_X67Y110_SLICE_X101Y110_A6 = CLBLM_R_X67Y111_SLICE_X101Y111_CO6;
  assign CLBLM_R_X67Y105_SLICE_X100Y105_A3 = CLBLM_L_X68Y103_SLICE_X102Y103_DQ;
  assign CLBLM_R_X67Y105_SLICE_X100Y105_A4 = CLBLM_L_X68Y105_SLICE_X102Y105_AO6;
  assign CLBLM_R_X67Y110_SLICE_X101Y110_B6 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLL_R_X71Y107_SLICE_X106Y107_A1 = 1'b1;
  assign CLBLL_R_X71Y107_SLICE_X106Y107_A2 = CLBLM_L_X72Y106_SLICE_X108Y106_CO6;
  assign CLBLL_R_X71Y107_SLICE_X106Y107_A3 = CLBLL_R_X71Y107_SLICE_X106Y107_AQ;
  assign CLBLL_R_X71Y107_SLICE_X106Y107_A4 = CLBLL_R_X71Y107_SLICE_X106Y107_BO6;
  assign CLBLL_R_X71Y107_SLICE_X106Y107_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y107_SLICE_X106Y107_A6 = CLBLL_R_X71Y108_SLICE_X106Y108_AQ;
  assign CLBLL_R_X71Y107_SLICE_X106Y107_B1 = CLBLL_R_X73Y108_SLICE_X110Y108_A5Q;
  assign CLBLL_R_X71Y107_SLICE_X106Y107_B2 = CLBLM_L_X62Y92_SLICE_X92Y92_AQ;
  assign CLBLL_R_X71Y107_SLICE_X106Y107_B3 = CLBLL_R_X71Y107_SLICE_X106Y107_CQ;
  assign CLBLL_R_X71Y107_SLICE_X106Y107_B4 = CLBLM_L_X70Y106_SLICE_X105Y106_CO6;
  assign CLBLL_R_X71Y107_SLICE_X106Y107_B5 = CLBLL_R_X71Y107_SLICE_X106Y107_C5Q;
  assign CLBLL_R_X71Y107_SLICE_X106Y107_B6 = 1'b1;
  assign CLBLM_R_X67Y110_SLICE_X101Y110_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y110_SLICE_X101Y110_C2 = CLBLM_R_X67Y110_SLICE_X101Y110_CQ;
  assign CLBLL_R_X71Y107_SLICE_X106Y107_C1 = CLBLL_R_X71Y107_SLICE_X106Y107_C5Q;
  assign CLBLL_R_X71Y107_SLICE_X106Y107_C2 = CLBLL_R_X71Y107_SLICE_X107Y107_C5Q;
  assign CLBLL_R_X71Y107_SLICE_X106Y107_C3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y107_SLICE_X106Y107_C4 = CLBLM_L_X70Y106_SLICE_X105Y106_CO6;
  assign CLBLL_R_X71Y107_SLICE_X106Y107_C5 = CLBLL_R_X71Y107_SLICE_X106Y107_CQ;
  assign CLBLL_R_X71Y107_SLICE_X106Y107_C6 = 1'b1;
  assign CLBLM_L_X78Y106_SLICE_X121Y106_A1 = 1'b1;
  assign CLBLM_L_X78Y106_SLICE_X121Y106_A2 = 1'b1;
  assign CLBLL_R_X71Y107_SLICE_X106Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X78Y106_SLICE_X121Y106_A3 = 1'b1;
  assign CLBLM_L_X78Y106_SLICE_X121Y106_A4 = 1'b1;
  assign CLBLM_L_X78Y106_SLICE_X121Y106_A5 = 1'b1;
  assign CLBLM_L_X78Y106_SLICE_X121Y106_A6 = 1'b1;
  assign CLBLL_R_X71Y107_SLICE_X106Y107_D1 = CLBLL_R_X71Y107_SLICE_X106Y107_C5Q;
  assign CLBLL_R_X71Y107_SLICE_X106Y107_D2 = CLBLM_L_X70Y107_SLICE_X105Y107_BQ;
  assign CLBLL_R_X71Y107_SLICE_X106Y107_D3 = CLBLL_R_X71Y107_SLICE_X107Y107_C5Q;
  assign CLBLL_R_X71Y107_SLICE_X106Y107_D4 = CLBLL_R_X71Y107_SLICE_X107Y107_CQ;
  assign CLBLL_R_X71Y107_SLICE_X106Y107_D5 = CLBLL_R_X71Y107_SLICE_X106Y107_CQ;
  assign CLBLL_R_X71Y107_SLICE_X106Y107_D6 = CLBLM_L_X70Y106_SLICE_X105Y106_CO6;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_C6 = CLBLL_R_X75Y124_SLICE_X115Y124_BQ;
  assign CLBLM_L_X78Y106_SLICE_X121Y106_B5 = 1'b1;
  assign CLBLL_R_X71Y107_SLICE_X106Y107_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X78Y106_SLICE_X121Y106_B6 = 1'b1;
  assign CLBLM_L_X78Y106_SLICE_X121Y106_C1 = 1'b1;
  assign CLBLM_L_X78Y106_SLICE_X121Y106_C2 = 1'b1;
  assign CLBLM_L_X78Y106_SLICE_X121Y106_C3 = 1'b1;
  assign CLBLM_L_X78Y106_SLICE_X121Y106_C4 = 1'b1;
  assign CLBLM_L_X78Y106_SLICE_X121Y106_C5 = 1'b1;
  assign CLBLM_L_X78Y106_SLICE_X121Y106_C6 = 1'b1;
  assign CLBLM_R_X67Y110_SLICE_X101Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X78Y106_SLICE_X121Y106_D1 = 1'b1;
  assign CLBLM_L_X78Y106_SLICE_X121Y106_D2 = 1'b1;
  assign CLBLM_L_X78Y106_SLICE_X121Y106_D3 = 1'b1;
  assign CLBLM_L_X78Y106_SLICE_X121Y106_D4 = 1'b1;
  assign CLBLM_L_X78Y106_SLICE_X121Y106_D5 = 1'b1;
  assign CLBLM_L_X78Y106_SLICE_X121Y106_D6 = 1'b1;
  assign CLBLL_R_X71Y107_SLICE_X107Y107_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y107_SLICE_X107Y107_A2 = CLBLM_L_X72Y108_SLICE_X109Y108_BO6;
  assign CLBLL_R_X71Y107_SLICE_X107Y107_A3 = CLBLL_R_X71Y107_SLICE_X107Y107_AQ;
  assign CLBLL_R_X71Y107_SLICE_X107Y107_A4 = CLBLM_L_X72Y108_SLICE_X108Y108_AQ;
  assign CLBLL_R_X71Y107_SLICE_X107Y107_A5 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLL_R_X71Y107_SLICE_X107Y107_A6 = CLBLL_R_X71Y109_SLICE_X106Y109_CO6;
  assign CLBLM_L_X78Y106_SLICE_X120Y106_A1 = 1'b1;
  assign CLBLM_L_X78Y106_SLICE_X120Y106_A2 = 1'b1;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_A2 = CLBLM_L_X70Y130_SLICE_X104Y130_BQ;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_A1 = CLBLM_L_X70Y128_SLICE_X105Y128_BO6;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_A4 = CLBLM_L_X70Y128_SLICE_X104Y128_BQ;
  assign CLBLL_R_X71Y107_SLICE_X107Y107_B1 = CLBLL_R_X71Y109_SLICE_X106Y109_CO6;
  assign CLBLL_R_X71Y107_SLICE_X107Y107_B2 = CLBLL_R_X71Y107_SLICE_X107Y107_BQ;
  assign CLBLL_R_X71Y107_SLICE_X107Y107_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y107_SLICE_X107Y107_B4 = CLBLL_R_X71Y107_SLICE_X107Y107_AQ;
  assign CLBLL_R_X71Y107_SLICE_X107Y107_B5 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLL_R_X71Y107_SLICE_X107Y107_B6 = CLBLM_L_X72Y108_SLICE_X109Y108_BO5;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_B1 = 1'b1;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_B2 = CLBLM_L_X70Y130_SLICE_X105Y130_BQ;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_B3 = CLBLM_L_X70Y129_SLICE_X104Y129_AQ;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_B4 = CLBLM_L_X70Y128_SLICE_X104Y128_BQ;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_B5 = CLBLM_L_X70Y128_SLICE_X104Y128_AQ;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_B6 = CLBLM_L_X70Y129_SLICE_X105Y129_CQ;
  assign CLBLL_R_X71Y107_SLICE_X107Y107_C1 = CLBLL_R_X71Y107_SLICE_X107Y107_C5Q;
  assign CLBLL_R_X71Y107_SLICE_X107Y107_C2 = CLBLL_R_X71Y107_SLICE_X107Y107_CQ;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_C1 = CLBLM_L_X70Y129_SLICE_X104Y129_AQ;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_C2 = 1'b1;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_C3 = CLBLM_L_X70Y130_SLICE_X105Y130_CQ;
  assign CLBLL_R_X71Y107_SLICE_X107Y107_C3 = CLBLL_R_X73Y108_SLICE_X110Y108_A5Q;
  assign CLBLL_R_X71Y107_SLICE_X107Y107_C4 = CLBLM_L_X72Y107_SLICE_X109Y107_DO6;
  assign CLBLL_R_X71Y107_SLICE_X107Y107_C5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y107_SLICE_X107Y107_C6 = 1'b1;
  assign CLBLL_R_X71Y107_SLICE_X107Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X71Y107_SLICE_X107Y107_D1 = CLBLM_L_X72Y107_SLICE_X108Y107_BQ;
  assign CLBLL_R_X71Y107_SLICE_X107Y107_D2 = CLBLM_L_X72Y107_SLICE_X109Y107_BQ;
  assign CLBLL_R_X71Y107_SLICE_X107Y107_D3 = CLBLM_L_X72Y108_SLICE_X108Y108_CQ;
  assign CLBLL_R_X71Y107_SLICE_X107Y107_D4 = CLBLL_R_X71Y107_SLICE_X106Y107_CQ;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_D1 = 1'b1;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_D2 = 1'b1;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_D3 = 1'b1;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_D4 = 1'b1;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_D5 = 1'b1;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_D6 = 1'b1;
  assign CLBLL_R_X71Y107_SLICE_X107Y107_D6 = CLBLL_R_X71Y107_SLICE_X107Y107_AQ;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X71Y107_SLICE_X107Y107_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X78Y106_SLICE_X120Y106_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_A1 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_A2 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_A3 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_A4 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_A5 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_A6 = 1'b1;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_A2 = CLBLM_L_X70Y128_SLICE_X104Y128_BQ;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_AX = CLBLM_L_X70Y128_SLICE_X104Y128_BO6;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_B1 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_B2 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_B3 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_B4 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_B5 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_B6 = 1'b1;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_B2 = 1'b1;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_B6 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_C1 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_C2 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_C3 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_C4 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_C5 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_C6 = 1'b1;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_BX = CLBLM_L_X70Y128_SLICE_X104Y128_AO5;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_C1 = CLBLM_L_X70Y128_SLICE_X104Y128_BQ;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_C2 = CLBLM_L_X70Y128_SLICE_X104Y128_CQ;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_C3 = CLBLM_L_X70Y128_SLICE_X105Y128_AO6;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_C4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_C5 = 1'b1;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_C6 = CLBLM_L_X70Y126_SLICE_X105Y126_CO6;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_D1 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_D2 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_D3 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_D4 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_D5 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_D6 = 1'b1;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_D1 = CLBLM_L_X70Y129_SLICE_X104Y129_AQ;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_D2 = CLBLM_L_X70Y128_SLICE_X104Y128_CQ;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_D3 = CLBLM_L_X70Y128_SLICE_X104Y128_DQ;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_D4 = CLBLM_L_X70Y128_SLICE_X104Y128_AQ;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_D5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_D6 = CLBLM_L_X70Y126_SLICE_X105Y126_CO6;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_A1 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_A2 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_A3 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_A4 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_A5 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_A6 = 1'b1;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_AX = CLBLL_R_X75Y127_SLICE_X115Y127_AQ;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_A4 = CLBLL_R_X79Y127_SLICE_X122Y127_CQ;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_B1 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_B2 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_B3 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_B4 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_B5 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_B6 = 1'b1;
  assign RIOI3_X105Y103_OLOGIC_X1Y103_D1 = CLBLL_R_X77Y128_SLICE_X119Y128_DQ;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_C1 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_C2 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_C3 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_C4 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_C5 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_C6 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X67Y110_SLICE_X100Y110_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_D1 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_D2 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_D3 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_D4 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_D5 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_D6 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X67Y110_SLICE_X100Y110_B5 = CLBLM_R_X65Y110_SLICE_X99Y110_AO6;
  assign CLBLM_R_X67Y110_SLICE_X100Y110_B6 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X76Y134_SLICE_X116Y134_D5 = CLBLL_R_X75Y134_SLICE_X115Y134_AO5;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_A5 = CLBLM_L_X72Y124_SLICE_X108Y124_BO6;
  assign CLBLL_R_X83Y132_SLICE_X130Y132_A1 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X130Y132_A2 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X130Y132_A3 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X130Y132_A4 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X130Y132_A5 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X130Y132_A6 = 1'b1;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_A6 = CLBLL_R_X73Y124_SLICE_X110Y124_BQ;
  assign CLBLM_R_X67Y110_SLICE_X100Y110_C3 = CLBLM_R_X65Y111_SLICE_X99Y111_AO5;
  assign CLBLL_R_X83Y132_SLICE_X130Y132_AX = CLBLM_L_X82Y130_SLICE_X128Y130_AQ;
  assign CLBLL_R_X83Y132_SLICE_X130Y132_B1 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X130Y132_B2 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X130Y132_B3 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X130Y132_B4 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X130Y132_B5 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X130Y132_B6 = 1'b1;
  assign CLBLM_R_X67Y110_SLICE_X100Y110_C5 = CLBLM_R_X65Y110_SLICE_X98Y110_DQ;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_T1 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X130Y132_C1 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X130Y132_C2 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X130Y132_C3 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X130Y132_C4 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X130Y132_C5 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X130Y132_C6 = 1'b1;
  assign CLBLM_R_X67Y110_SLICE_X100Y110_C6 = CLBLM_R_X67Y111_SLICE_X101Y111_DO5;
  assign CLBLL_R_X83Y132_SLICE_X130Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X83Y132_SLICE_X130Y132_D1 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X130Y132_D2 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X130Y132_D3 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X130Y132_D4 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X130Y132_D5 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X130Y132_D6 = 1'b1;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_A5 = CLBLM_L_X76Y123_SLICE_X116Y123_AQ;
  assign CLBLM_R_X67Y110_SLICE_X100Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X71Y108_SLICE_X106Y108_A1 = CLBLL_R_X71Y109_SLICE_X106Y109_B5Q;
  assign CLBLL_R_X71Y108_SLICE_X106Y108_A2 = CLBLL_R_X71Y109_SLICE_X106Y109_BQ;
  assign CLBLL_R_X71Y108_SLICE_X106Y108_A3 = CLBLL_R_X71Y108_SLICE_X106Y108_AQ;
  assign CLBLL_R_X71Y108_SLICE_X106Y108_A4 = CLBLM_L_X72Y108_SLICE_X109Y108_A5Q;
  assign CLBLL_R_X71Y108_SLICE_X106Y108_A5 = CLBLL_R_X71Y108_SLICE_X107Y108_AQ;
  assign CLBLL_R_X71Y108_SLICE_X106Y108_A6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X83Y132_SLICE_X130Y132_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_B3 = CLBLM_L_X72Y124_SLICE_X109Y124_AQ;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y108_SLICE_X106Y108_B1 = 1'b1;
  assign CLBLL_R_X71Y108_SLICE_X106Y108_B2 = CLBLL_R_X71Y108_SLICE_X106Y108_BQ;
  assign CLBLL_R_X71Y108_SLICE_X106Y108_B3 = CLBLL_R_X71Y108_SLICE_X106Y108_AQ;
  assign CLBLL_R_X71Y108_SLICE_X106Y108_B4 = CLBLL_R_X71Y107_SLICE_X106Y107_BO6;
  assign CLBLL_R_X71Y108_SLICE_X106Y108_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y108_SLICE_X106Y108_B6 = CLBLL_R_X71Y107_SLICE_X106Y107_AQ;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_B5 = CLBLM_L_X72Y124_SLICE_X108Y124_BO6;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_B6 = CLBLL_R_X73Y124_SLICE_X110Y124_BQ;
  assign CLBLL_R_X71Y108_SLICE_X106Y108_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y108_SLICE_X106Y108_C2 = CLBLL_R_X71Y108_SLICE_X106Y108_CQ;
  assign CLBLL_R_X71Y108_SLICE_X106Y108_C3 = CLBLM_L_X72Y108_SLICE_X109Y108_A5Q;
  assign CLBLL_R_X71Y108_SLICE_X106Y108_C4 = CLBLL_R_X71Y108_SLICE_X106Y108_BQ;
  assign CLBLL_R_X71Y108_SLICE_X106Y108_C5 = CLBLL_R_X71Y109_SLICE_X106Y109_B5Q;
  assign CLBLL_R_X71Y108_SLICE_X106Y108_C6 = CLBLL_R_X71Y109_SLICE_X106Y109_BQ;
  assign CLBLL_R_X83Y132_SLICE_X131Y132_A1 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X131Y132_A2 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X131Y132_A3 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X131Y132_A4 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X131Y132_A5 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X131Y132_A6 = 1'b1;
  assign CLBLL_R_X71Y108_SLICE_X106Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X71Y108_SLICE_X106Y108_D1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X83Y132_SLICE_X131Y132_B1 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X131Y132_B2 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X131Y132_B3 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X131Y132_B4 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X131Y132_B5 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X131Y132_B6 = 1'b1;
  assign CLBLL_R_X71Y108_SLICE_X106Y108_D2 = CLBLL_R_X71Y108_SLICE_X106Y108_CQ;
  assign CLBLL_R_X71Y108_SLICE_X106Y108_D3 = CLBLL_R_X71Y108_SLICE_X106Y108_DQ;
  assign CLBLL_R_X71Y108_SLICE_X106Y108_D4 = CLBLL_R_X71Y107_SLICE_X106Y107_BO6;
  assign CLBLL_R_X71Y108_SLICE_X106Y108_D5 = CLBLL_R_X71Y108_SLICE_X106Y108_D5Q;
  assign CLBLL_R_X71Y108_SLICE_X106Y108_D6 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X131Y132_C2 = 1'b1;
  assign CLBLL_R_X71Y108_SLICE_X106Y108_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X83Y132_SLICE_X131Y132_C1 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X131Y132_C3 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X131Y132_C4 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X131Y132_C5 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X131Y132_C6 = 1'b1;
  assign CLBLM_R_X67Y110_SLICE_X100Y110_D4 = CLBLM_R_X67Y110_SLICE_X100Y110_BQ;
  assign CLBLM_R_X67Y110_SLICE_X100Y110_D5 = CLBLM_R_X65Y110_SLICE_X99Y110_B5Q;
  assign CLBLM_R_X67Y110_SLICE_X100Y110_D6 = CLBLM_L_X60Y97_SLICE_X91Y97_AQ;
  assign CLBLL_R_X83Y132_SLICE_X131Y132_D1 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X131Y132_D2 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X131Y132_D3 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X131Y132_D4 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X131Y132_D5 = 1'b1;
  assign CLBLL_R_X83Y132_SLICE_X131Y132_D6 = 1'b1;
  assign CLBLL_R_X71Y108_SLICE_X107Y108_A1 = CLBLL_R_X71Y109_SLICE_X106Y109_B5Q;
  assign CLBLL_R_X71Y108_SLICE_X107Y108_A2 = CLBLM_L_X72Y108_SLICE_X109Y108_A5Q;
  assign CLBLL_R_X71Y108_SLICE_X107Y108_A3 = CLBLL_R_X71Y108_SLICE_X107Y108_AQ;
  assign CLBLL_R_X71Y108_SLICE_X107Y108_A4 = CLBLL_R_X71Y109_SLICE_X106Y109_BQ;
  assign CLBLL_R_X71Y108_SLICE_X107Y108_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y108_SLICE_X107Y108_A6 = CLBLL_R_X79Y99_SLICE_X122Y99_AO6;
  assign CLBLL_R_X71Y108_SLICE_X107Y108_AX = CLBLM_L_X72Y109_SLICE_X109Y109_DQ;
  assign CLBLL_R_X71Y108_SLICE_X107Y108_B1 = 1'b1;
  assign CLBLL_R_X71Y108_SLICE_X107Y108_B2 = 1'b1;
  assign CLBLL_R_X71Y108_SLICE_X107Y108_B3 = 1'b1;
  assign CLBLL_R_X71Y108_SLICE_X107Y108_B4 = 1'b1;
  assign CLBLL_R_X71Y108_SLICE_X107Y108_B5 = 1'b1;
  assign CLBLL_R_X71Y108_SLICE_X107Y108_B6 = 1'b1;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_A1 = CLBLM_L_X70Y130_SLICE_X104Y130_AO6;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_A2 = CLBLM_L_X70Y129_SLICE_X105Y129_BQ;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_A6 = CLBLM_L_X72Y133_SLICE_X109Y133_AO6;
  assign CLBLL_R_X71Y108_SLICE_X107Y108_C1 = 1'b1;
  assign CLBLL_R_X71Y108_SLICE_X107Y108_C2 = 1'b1;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_B1 = CLBLM_L_X70Y129_SLICE_X105Y129_CQ;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_B2 = CLBLM_L_X70Y129_SLICE_X105Y129_BQ;
  assign CLBLL_R_X71Y108_SLICE_X107Y108_C3 = 1'b1;
  assign CLBLL_R_X71Y108_SLICE_X107Y108_C4 = 1'b1;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_B5 = CLBLL_R_X71Y130_SLICE_X106Y130_AO6;
  assign CLBLL_R_X71Y108_SLICE_X107Y108_C5 = 1'b1;
  assign CLBLL_R_X71Y108_SLICE_X107Y108_C6 = 1'b1;
  assign CLBLL_R_X71Y108_SLICE_X107Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_C2 = CLBLM_L_X70Y129_SLICE_X105Y129_CQ;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_C3 = CLBLM_L_X70Y130_SLICE_X105Y130_CQ;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_C4 = CLBLM_L_X72Y133_SLICE_X109Y133_AO6;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_C5 = CLBLM_L_X72Y132_SLICE_X109Y132_AO6;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_C6 = CLBLM_L_X70Y130_SLICE_X105Y130_DO5;
  assign CLBLL_R_X71Y108_SLICE_X107Y108_D1 = 1'b1;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X71Y108_SLICE_X107Y108_D2 = 1'b1;
  assign CLBLL_R_X71Y108_SLICE_X107Y108_D3 = 1'b1;
  assign CLBLL_R_X71Y108_SLICE_X107Y108_D4 = 1'b1;
  assign CLBLL_R_X71Y108_SLICE_X107Y108_D5 = 1'b1;
  assign CLBLL_R_X71Y108_SLICE_X107Y108_D6 = 1'b1;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_D1 = CLBLM_L_X70Y130_SLICE_X105Y130_A5Q;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_D2 = CLBLM_L_X70Y130_SLICE_X105Y130_AQ;
  assign CLBLL_R_X71Y108_SLICE_X107Y108_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_D5 = CLBLM_L_X70Y130_SLICE_X104Y130_DQ;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_D6 = CLBLM_L_X72Y132_SLICE_X109Y132_AO6;
  assign CLBLL_R_X79Y104_SLICE_X122Y104_A1 = CLBLM_L_X72Y118_SLICE_X108Y118_A5Q;
  assign CLBLL_R_X79Y104_SLICE_X122Y104_A2 = 1'b1;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X79Y104_SLICE_X122Y104_A4 = CLBLL_R_X75Y124_SLICE_X115Y124_BQ;
  assign CLBLL_R_X79Y104_SLICE_X122Y104_A5 = CLBLM_R_X103Y69_SLICE_X162Y69_A5Q;
  assign CLBLL_R_X79Y104_SLICE_X122Y104_A6 = CLBLL_R_X77Y104_SLICE_X118Y104_CQ;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_A1 = CLBLM_L_X70Y128_SLICE_X104Y128_BQ;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_A2 = CLBLM_L_X70Y129_SLICE_X104Y129_BQ;
  assign CLBLL_R_X79Y104_SLICE_X122Y104_AX = CLBLL_R_X75Y103_SLICE_X115Y103_AQ;
  assign CLBLL_R_X79Y104_SLICE_X122Y104_B1 = CLBLM_L_X72Y118_SLICE_X108Y118_A5Q;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_A6 = CLBLM_L_X70Y126_SLICE_X105Y126_CO6;
  assign CLBLL_R_X79Y104_SLICE_X122Y104_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X79Y104_SLICE_X122Y104_B4 = CLBLM_R_X103Y76_SLICE_X162Y76_AO6;
  assign CLBLL_R_X79Y104_SLICE_X122Y104_B5 = CLBLM_R_X103Y76_SLICE_X162Y76_BQ;
  assign CLBLL_R_X79Y104_SLICE_X122Y104_B6 = CLBLL_R_X77Y104_SLICE_X118Y104_CQ;
  assign CLBLL_R_X79Y104_SLICE_X122Y104_C1 = 1'b1;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_B2 = CLBLM_L_X70Y129_SLICE_X104Y129_BQ;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_B3 = CLBLM_L_X70Y128_SLICE_X104Y128_AO6;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_B5 = CLBLM_L_X70Y129_SLICE_X105Y129_AQ;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_B6 = CLBLM_L_X70Y126_SLICE_X105Y126_CO6;
  assign CLBLL_R_X79Y104_SLICE_X122Y104_C4 = 1'b1;
  assign CLBLL_R_X79Y104_SLICE_X122Y104_C5 = 1'b1;
  assign CLBLL_R_X79Y104_SLICE_X122Y104_C6 = 1'b1;
  assign CLBLL_R_X79Y104_SLICE_X122Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X79Y104_SLICE_X122Y104_D1 = 1'b1;
  assign CLBLL_R_X79Y104_SLICE_X122Y104_D2 = 1'b1;
  assign CLBLL_R_X79Y104_SLICE_X122Y104_D3 = 1'b1;
  assign CLBLL_R_X79Y104_SLICE_X122Y104_D4 = 1'b1;
  assign CLBLL_R_X79Y104_SLICE_X122Y104_D5 = 1'b1;
  assign CLBLL_R_X79Y104_SLICE_X122Y104_D6 = 1'b1;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_A6 = CLBLM_L_X62Y106_SLICE_X93Y106_CQ;
  assign CLBLL_R_X79Y104_SLICE_X122Y104_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_C2 = CLBLM_L_X70Y129_SLICE_X104Y129_CQ;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_C3 = 1'b1;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_C4 = CLBLM_L_X70Y128_SLICE_X104Y128_DQ;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_C5 = CLBLM_L_X70Y128_SLICE_X104Y128_BO5;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_C6 = CLBLM_L_X70Y131_SLICE_X104Y131_BQ;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_D1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_D2 = CLBLM_L_X70Y129_SLICE_X104Y129_CQ;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_AX = CLBLM_L_X60Y104_SLICE_X90Y104_AQ;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_D3 = CLBLM_L_X70Y129_SLICE_X104Y129_DQ;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_D4 = CLBLM_L_X70Y126_SLICE_X105Y126_CO6;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_D5 = CLBLM_L_X70Y129_SLICE_X104Y129_AQ;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_D6 = CLBLM_L_X70Y128_SLICE_X104Y128_BQ;
  assign CLBLM_L_X78Y104_SLICE_X120Y104_C2 = 1'b1;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X78Y104_SLICE_X120Y104_C3 = 1'b1;
  assign CLBLM_L_X78Y104_SLICE_X120Y104_C4 = 1'b1;
  assign CLBLL_R_X79Y104_SLICE_X123Y104_A1 = 1'b1;
  assign CLBLL_R_X79Y104_SLICE_X123Y104_A2 = 1'b1;
  assign CLBLL_R_X79Y104_SLICE_X123Y104_A3 = 1'b1;
  assign CLBLL_R_X79Y104_SLICE_X123Y104_A4 = 1'b1;
  assign CLBLL_R_X79Y104_SLICE_X123Y104_A5 = 1'b1;
  assign CLBLL_R_X79Y104_SLICE_X123Y104_A6 = 1'b1;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_B3 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X78Y104_SLICE_X120Y104_C5 = 1'b1;
  assign CLBLM_L_X78Y104_SLICE_X120Y104_C6 = 1'b1;
  assign CLBLL_R_X79Y104_SLICE_X123Y104_B1 = 1'b1;
  assign CLBLL_R_X79Y104_SLICE_X123Y104_B2 = 1'b1;
  assign CLBLL_R_X79Y104_SLICE_X123Y104_B3 = 1'b1;
  assign CLBLL_R_X79Y104_SLICE_X123Y104_B4 = 1'b1;
  assign CLBLL_R_X79Y104_SLICE_X123Y104_B5 = 1'b1;
  assign CLBLL_R_X79Y104_SLICE_X123Y104_B6 = 1'b1;
  assign CLBLM_R_X67Y110_SLICE_X101Y110_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X79Y104_SLICE_X123Y104_C1 = 1'b1;
  assign CLBLL_R_X79Y104_SLICE_X123Y104_C2 = 1'b1;
  assign CLBLL_R_X79Y104_SLICE_X123Y104_C3 = 1'b1;
  assign CLBLL_R_X79Y104_SLICE_X123Y104_C4 = 1'b1;
  assign CLBLL_R_X79Y104_SLICE_X123Y104_C5 = 1'b1;
  assign CLBLL_R_X79Y104_SLICE_X123Y104_C6 = 1'b1;
  assign CLBLL_R_X79Y104_SLICE_X123Y104_D1 = 1'b1;
  assign CLBLL_R_X79Y104_SLICE_X123Y104_D2 = 1'b1;
  assign CLBLL_R_X79Y104_SLICE_X123Y104_D3 = 1'b1;
  assign CLBLL_R_X79Y104_SLICE_X123Y104_D4 = 1'b1;
  assign CLBLL_R_X79Y104_SLICE_X123Y104_D5 = 1'b1;
  assign CLBLL_R_X79Y104_SLICE_X123Y104_D6 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_C1 = 1'b1;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_C2 = CLBLM_L_X62Y105_SLICE_X93Y105_CQ;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_C4 = 1'b1;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_C3 = CLBLM_L_X64Y105_SLICE_X96Y105_BO5;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_C4 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_C6 = 1'b1;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_C5 = CLBLM_L_X62Y105_SLICE_X93Y105_AQ;
  assign CLBLM_L_X78Y104_SLICE_X120Y104_D3 = 1'b1;
  assign CLBLM_L_X78Y104_SLICE_X120Y104_D4 = 1'b1;
  assign CLBLM_L_X78Y104_SLICE_X120Y104_D5 = 1'b1;
  assign CLBLM_L_X78Y104_SLICE_X120Y104_D6 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_D3 = 1'b1;
  assign CLBLL_R_X71Y109_SLICE_X106Y109_A1 = 1'b1;
  assign CLBLL_R_X71Y109_SLICE_X106Y109_A2 = CLBLL_R_X71Y110_SLICE_X106Y110_BQ;
  assign CLBLL_R_X71Y109_SLICE_X106Y109_A3 = CLBLL_R_X71Y109_SLICE_X106Y109_AQ;
  assign CLBLL_R_X71Y109_SLICE_X106Y109_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y109_SLICE_X106Y109_A5 = CLBLL_R_X71Y109_SLICE_X106Y109_CO5;
  assign CLBLL_R_X71Y109_SLICE_X106Y109_A6 = CLBLL_R_X71Y110_SLICE_X106Y110_AQ;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_D4 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_D5 = 1'b1;
  assign LIOB33_X0Y187_IOB_X0Y187_O = 1'b1;
  assign CLBLL_R_X71Y109_SLICE_X106Y109_B1 = CLBLL_R_X71Y109_SLICE_X106Y109_B5Q;
  assign CLBLL_R_X71Y109_SLICE_X106Y109_B2 = 1'b1;
  assign CLBLL_R_X71Y109_SLICE_X106Y109_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y109_SLICE_X106Y109_B4 = CLBLM_L_X72Y108_SLICE_X109Y108_A5Q;
  assign CLBLL_R_X71Y109_SLICE_X106Y109_B5 = CLBLL_R_X71Y109_SLICE_X106Y109_BQ;
  assign CLBLL_R_X71Y109_SLICE_X106Y109_B6 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_D6 = 1'b1;
  assign CLBLL_R_X71Y109_SLICE_X106Y109_C1 = CLBLL_R_X71Y109_SLICE_X106Y109_BQ;
  assign CLBLL_R_X71Y109_SLICE_X106Y109_C2 = 1'b1;
  assign CLBLL_R_X71Y109_SLICE_X106Y109_C3 = 1'b1;
  assign CLBLL_R_X71Y109_SLICE_X106Y109_C4 = CLBLM_L_X72Y108_SLICE_X109Y108_A5Q;
  assign CLBLL_R_X71Y109_SLICE_X106Y109_C5 = CLBLL_R_X71Y109_SLICE_X106Y109_B5Q;
  assign CLBLL_R_X71Y109_SLICE_X106Y109_C6 = 1'b1;
  assign CLBLL_R_X71Y109_SLICE_X106Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOB33_X105Y169_IOB_X1Y170_O = 1'b1;
  assign RIOB33_X105Y169_IOB_X1Y169_O = 1'b1;
  assign CLBLL_R_X71Y109_SLICE_X106Y109_D1 = 1'b1;
  assign CLBLL_R_X71Y109_SLICE_X106Y109_D2 = 1'b1;
  assign CLBLL_R_X71Y109_SLICE_X106Y109_D3 = 1'b1;
  assign CLBLL_R_X71Y109_SLICE_X106Y109_D4 = 1'b1;
  assign CLBLL_R_X71Y109_SLICE_X106Y109_D5 = 1'b1;
  assign CLBLL_R_X71Y109_SLICE_X106Y109_D6 = 1'b1;
  assign CLBLL_R_X71Y109_SLICE_X106Y109_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_A1 = CLBLM_R_X65Y105_SLICE_X99Y105_CQ;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_A2 = CLBLM_L_X74Y119_SLICE_X112Y119_CQ;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_A3 = CLBLM_L_X72Y118_SLICE_X108Y118_CQ;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_A4 = CLBLM_L_X74Y120_SLICE_X112Y120_BO6;
  assign CLBLL_R_X71Y109_SLICE_X107Y109_A1 = 1'b1;
  assign CLBLL_R_X71Y109_SLICE_X107Y109_A2 = 1'b1;
  assign CLBLL_R_X71Y109_SLICE_X107Y109_A3 = 1'b1;
  assign CLBLL_R_X71Y109_SLICE_X107Y109_A4 = 1'b1;
  assign CLBLL_R_X71Y109_SLICE_X107Y109_A5 = 1'b1;
  assign CLBLL_R_X71Y109_SLICE_X107Y109_A6 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_A5 = CLBLM_L_X74Y121_SLICE_X113Y121_AQ;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_A6 = CLBLM_L_X74Y120_SLICE_X112Y120_CO6;
  assign CLBLL_R_X71Y109_SLICE_X107Y109_B1 = 1'b1;
  assign CLBLL_R_X71Y109_SLICE_X107Y109_B2 = 1'b1;
  assign CLBLL_R_X71Y109_SLICE_X107Y109_B3 = 1'b1;
  assign CLBLL_R_X71Y109_SLICE_X107Y109_B4 = 1'b1;
  assign CLBLL_R_X71Y109_SLICE_X107Y109_B5 = 1'b1;
  assign CLBLL_R_X71Y109_SLICE_X107Y109_B6 = 1'b1;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_A5 = 1'b1;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_A6 = 1'b1;
  assign CLBLM_L_X70Y130_SLICE_X105Y130_A1 = CLBLM_L_X72Y132_SLICE_X109Y132_AO6;
  assign CLBLM_L_X70Y130_SLICE_X105Y130_A2 = CLBLM_L_X70Y130_SLICE_X105Y130_A5Q;
  assign CLBLM_L_X70Y130_SLICE_X105Y130_A3 = CLBLM_L_X70Y130_SLICE_X105Y130_AQ;
  assign CLBLM_L_X70Y130_SLICE_X105Y130_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y130_SLICE_X105Y130_A5 = CLBLL_R_X71Y130_SLICE_X106Y130_AQ;
  assign CLBLM_L_X70Y130_SLICE_X105Y130_A6 = 1'b1;
  assign CLBLL_R_X71Y109_SLICE_X107Y109_C1 = 1'b1;
  assign CLBLL_R_X71Y109_SLICE_X107Y109_C2 = 1'b1;
  assign CLBLM_L_X70Y130_SLICE_X105Y130_B1 = CLBLM_L_X72Y133_SLICE_X109Y133_AO6;
  assign CLBLM_L_X70Y130_SLICE_X105Y130_B2 = CLBLM_L_X70Y130_SLICE_X105Y130_BQ;
  assign CLBLM_L_X70Y130_SLICE_X105Y130_B3 = CLBLM_L_X70Y130_SLICE_X104Y130_AO6;
  assign CLBLM_L_X70Y130_SLICE_X105Y130_B4 = CLBLM_L_X70Y130_SLICE_X104Y130_BQ;
  assign CLBLM_L_X70Y130_SLICE_X105Y130_B5 = CLBLL_R_X71Y130_SLICE_X106Y130_AQ;
  assign CLBLM_L_X70Y130_SLICE_X105Y130_B6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y109_SLICE_X107Y109_C6 = 1'b1;
  assign CLBLL_R_X71Y109_SLICE_X107Y109_D1 = 1'b1;
  assign CLBLM_L_X70Y130_SLICE_X105Y130_C1 = CLBLM_L_X70Y130_SLICE_X105Y130_BQ;
  assign CLBLM_L_X70Y130_SLICE_X105Y130_C2 = CLBLM_L_X70Y130_SLICE_X105Y130_CQ;
  assign CLBLM_L_X70Y130_SLICE_X105Y130_C3 = CLBLL_R_X71Y130_SLICE_X106Y130_AQ;
  assign CLBLM_L_X70Y130_SLICE_X105Y130_C4 = CLBLM_L_X72Y133_SLICE_X109Y133_AO6;
  assign CLBLM_L_X70Y130_SLICE_X105Y130_C5 = CLBLM_L_X70Y130_SLICE_X105Y130_DO6;
  assign CLBLM_L_X70Y130_SLICE_X105Y130_C6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y109_SLICE_X107Y109_D2 = 1'b1;
  assign CLBLL_R_X71Y109_SLICE_X107Y109_D3 = 1'b1;
  assign CLBLM_L_X70Y130_SLICE_X105Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X71Y109_SLICE_X107Y109_D4 = 1'b1;
  assign CLBLL_R_X71Y109_SLICE_X107Y109_D5 = 1'b1;
  assign CLBLL_R_X71Y109_SLICE_X107Y109_D6 = 1'b1;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_B1 = 1'b1;
  assign CLBLM_L_X70Y130_SLICE_X105Y130_D1 = 1'b1;
  assign CLBLM_L_X70Y130_SLICE_X105Y130_D2 = CLBLM_L_X72Y132_SLICE_X109Y132_AO6;
  assign CLBLM_L_X70Y130_SLICE_X105Y130_D3 = CLBLL_R_X71Y130_SLICE_X106Y130_AQ;
  assign CLBLM_L_X70Y130_SLICE_X105Y130_D4 = CLBLM_L_X70Y130_SLICE_X105Y130_A5Q;
  assign CLBLM_L_X70Y130_SLICE_X105Y130_D5 = 1'b1;
  assign CLBLM_L_X70Y130_SLICE_X105Y130_D6 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_B4 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_B5 = 1'b1;
  assign CLBLM_L_X70Y130_SLICE_X105Y130_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_B6 = CLBLL_R_X75Y122_SLICE_X115Y122_AQ;
  assign CLBLM_L_X70Y130_SLICE_X104Y130_A1 = CLBLM_L_X70Y130_SLICE_X105Y130_A5Q;
  assign CLBLM_L_X70Y130_SLICE_X104Y130_A2 = CLBLM_L_X72Y132_SLICE_X109Y132_AO6;
  assign CLBLM_L_X70Y130_SLICE_X104Y130_A3 = 1'b1;
  assign CLBLM_L_X70Y130_SLICE_X104Y130_A4 = 1'b1;
  assign CLBLM_L_X70Y130_SLICE_X104Y130_A5 = CLBLM_L_X70Y130_SLICE_X105Y130_AQ;
  assign CLBLM_L_X70Y130_SLICE_X104Y130_A6 = 1'b1;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_B5 = 1'b1;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_B6 = 1'b1;
  assign CLBLM_L_X70Y110_SLICE_X105Y110_C3 = 1'b1;
  assign CLBLM_L_X70Y110_SLICE_X105Y110_C4 = 1'b1;
  assign CLBLM_L_X70Y130_SLICE_X104Y130_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y130_SLICE_X104Y130_B2 = CLBLM_L_X70Y130_SLICE_X104Y130_BQ;
  assign CLBLM_L_X70Y130_SLICE_X104Y130_B3 = 1'b1;
  assign CLBLM_L_X70Y130_SLICE_X104Y130_B4 = CLBLM_L_X70Y131_SLICE_X104Y131_BQ;
  assign CLBLM_L_X70Y130_SLICE_X104Y130_B5 = CLBLM_L_X72Y133_SLICE_X109Y133_AO6;
  assign CLBLM_L_X70Y130_SLICE_X104Y130_B6 = CLBLM_L_X70Y130_SLICE_X104Y130_AO5;
  assign CLBLM_L_X70Y110_SLICE_X105Y110_C5 = 1'b1;
  assign CLBLM_L_X70Y110_SLICE_X105Y110_C6 = 1'b1;
  assign CLBLM_L_X70Y130_SLICE_X104Y130_C1 = CLBLM_L_X70Y130_SLICE_X105Y130_AQ;
  assign CLBLM_L_X70Y130_SLICE_X104Y130_C2 = CLBLM_L_X70Y130_SLICE_X104Y130_CQ;
  assign CLBLM_L_X70Y130_SLICE_X104Y130_C3 = CLBLM_L_X72Y132_SLICE_X109Y132_AO6;
  assign CLBLM_L_X70Y130_SLICE_X104Y130_C4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y130_SLICE_X104Y130_C5 = CLBLM_L_X70Y130_SLICE_X105Y130_A5Q;
  assign CLBLM_L_X70Y130_SLICE_X104Y130_C6 = CLBLM_L_X70Y129_SLICE_X104Y129_DQ;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_C1 = 1'b1;
  assign CLBLM_L_X70Y130_SLICE_X104Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_C2 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_C3 = 1'b1;
  assign CLBLM_L_X70Y130_SLICE_X104Y130_D1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y130_SLICE_X104Y130_D2 = CLBLM_L_X70Y130_SLICE_X104Y130_CQ;
  assign CLBLM_L_X70Y130_SLICE_X104Y130_D3 = CLBLM_L_X70Y130_SLICE_X104Y130_DQ;
  assign CLBLM_L_X70Y130_SLICE_X104Y130_D4 = CLBLM_L_X70Y130_SLICE_X104Y130_AO5;
  assign CLBLM_L_X70Y130_SLICE_X104Y130_D5 = 1'b1;
  assign CLBLM_L_X70Y130_SLICE_X104Y130_D6 = CLBLM_L_X70Y129_SLICE_X104Y129_DQ;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_C4 = CLBLM_L_X76Y125_SLICE_X116Y125_C5Q;
  assign CLBLM_L_X70Y130_SLICE_X104Y130_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_C5 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_C6 = CLBLM_L_X76Y122_SLICE_X116Y122_CQ;
  assign CLBLM_L_X70Y110_SLICE_X105Y110_D1 = 1'b1;
  assign CLBLM_R_X67Y97_SLICE_X101Y97_A1 = CLBLM_R_X67Y97_SLICE_X101Y97_AQ;
  assign CLBLM_L_X70Y110_SLICE_X105Y110_D2 = 1'b1;
  assign CLBLM_L_X70Y110_SLICE_X105Y110_D3 = 1'b1;
  assign CLBLM_L_X70Y110_SLICE_X105Y110_D4 = 1'b1;
  assign CLBLM_L_X70Y110_SLICE_X105Y110_D5 = 1'b1;
  assign CLBLM_L_X70Y110_SLICE_X105Y110_D6 = 1'b1;
  assign CLBLM_R_X67Y97_SLICE_X101Y97_A2 = CLBLM_R_X67Y98_SLICE_X101Y98_AO6;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_D1 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_D2 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_D1 = CLBLL_R_X73Y131_SLICE_X110Y131_AQ;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_D3 = 1'b1;
  assign CLBLM_R_X67Y97_SLICE_X101Y97_A3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_D4 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_T1 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_D5 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_D1 = CLBLM_L_X70Y111_SLICE_X105Y111_DO6;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_D6 = 1'b1;
  assign CLBLM_L_X70Y110_SLICE_X104Y110_A1 = CLBLM_L_X70Y110_SLICE_X104Y110_B5Q;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_D1 = CLBLL_L_X34Y126_SLICE_X50Y126_AO6;
  assign CLBLM_L_X70Y110_SLICE_X104Y110_A2 = CLBLM_L_X70Y110_SLICE_X104Y110_BQ;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_T1 = 1'b1;
  assign CLBLM_L_X70Y110_SLICE_X104Y110_A3 = CLBLM_L_X70Y110_SLICE_X104Y110_AQ;
  assign CLBLM_R_X67Y97_SLICE_X101Y97_A4 = CLBLM_R_X67Y96_SLICE_X101Y96_AQ;
  assign CLBLM_L_X70Y110_SLICE_X104Y110_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_T1 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_D1 = 1'b1;
  assign CLBLM_L_X70Y110_SLICE_X104Y110_A5 = CLBLM_L_X70Y111_SLICE_X104Y111_CO6;
  assign CLBLM_L_X70Y110_SLICE_X104Y110_A6 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_T1 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_B2 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_C3 = 1'b1;
  assign CLBLM_R_X67Y97_SLICE_X101Y97_A5 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_C4 = 1'b1;
  assign CLBLL_R_X71Y110_SLICE_X106Y110_A1 = CLBLL_R_X71Y108_SLICE_X106Y108_D5Q;
  assign CLBLL_R_X71Y110_SLICE_X106Y110_A2 = CLBLL_R_X71Y114_SLICE_X106Y114_AQ;
  assign CLBLL_R_X71Y110_SLICE_X106Y110_A3 = CLBLL_R_X71Y110_SLICE_X106Y110_AQ;
  assign CLBLL_R_X71Y110_SLICE_X106Y110_A4 = CLBLL_R_X71Y107_SLICE_X106Y107_BO6;
  assign CLBLL_R_X71Y110_SLICE_X106Y110_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y110_SLICE_X106Y110_A6 = 1'b1;
  assign LIOB33_SING_X0Y199_IOB_X0Y199_O = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_B5 = 1'b1;
  assign CLBLL_R_X71Y110_SLICE_X106Y110_B1 = CLBLL_R_X71Y109_SLICE_X106Y109_B5Q;
  assign CLBLL_R_X71Y110_SLICE_X106Y110_B2 = CLBLL_R_X71Y110_SLICE_X106Y110_BQ;
  assign CLBLL_R_X71Y110_SLICE_X106Y110_B3 = CLBLL_R_X71Y110_SLICE_X106Y110_AQ;
  assign CLBLL_R_X71Y110_SLICE_X106Y110_B4 = CLBLM_L_X72Y108_SLICE_X109Y108_A5Q;
  assign CLBLL_R_X71Y110_SLICE_X106Y110_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y110_SLICE_X106Y110_B6 = CLBLL_R_X71Y109_SLICE_X106Y109_BQ;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_C6 = 1'b1;
  assign CLBLL_R_X71Y110_SLICE_X106Y110_C1 = 1'b1;
  assign CLBLL_R_X71Y110_SLICE_X106Y110_C2 = 1'b1;
  assign CLBLL_R_X71Y110_SLICE_X106Y110_C3 = 1'b1;
  assign CLBLL_R_X71Y110_SLICE_X106Y110_C4 = 1'b1;
  assign CLBLL_R_X71Y110_SLICE_X106Y110_C5 = 1'b1;
  assign CLBLL_R_X71Y110_SLICE_X106Y110_C6 = 1'b1;
  assign CLBLM_L_X70Y110_SLICE_X104Y110_B3 = CLBLM_L_X70Y110_SLICE_X104Y110_AQ;
  assign CLBLM_R_X67Y97_SLICE_X101Y97_A6 = CLBLM_R_X67Y98_SLICE_X101Y98_CO6;
  assign CLBLL_R_X71Y110_SLICE_X106Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X71Y110_SLICE_X106Y110_D1 = 1'b1;
  assign CLBLL_R_X71Y110_SLICE_X106Y110_D2 = 1'b1;
  assign CLBLL_R_X71Y110_SLICE_X106Y110_D3 = 1'b1;
  assign CLBLL_R_X71Y110_SLICE_X106Y110_D4 = 1'b1;
  assign CLBLL_R_X71Y110_SLICE_X106Y110_D5 = 1'b1;
  assign CLBLL_R_X71Y110_SLICE_X106Y110_D6 = 1'b1;
  assign CLBLM_L_X70Y110_SLICE_X104Y110_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y110_SLICE_X106Y110_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_D1 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_D2 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_D3 = 1'b1;
  assign CLBLL_R_X71Y110_SLICE_X107Y110_A1 = 1'b1;
  assign CLBLL_R_X71Y110_SLICE_X107Y110_A2 = 1'b1;
  assign CLBLL_R_X71Y110_SLICE_X107Y110_A3 = 1'b1;
  assign CLBLL_R_X71Y110_SLICE_X107Y110_A4 = 1'b1;
  assign CLBLL_R_X71Y110_SLICE_X107Y110_A5 = 1'b1;
  assign CLBLL_R_X71Y110_SLICE_X107Y110_A6 = 1'b1;
  assign CLBLM_L_X70Y110_SLICE_X104Y110_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_D4 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_D5 = 1'b1;
  assign CLBLL_R_X71Y110_SLICE_X107Y110_B1 = 1'b1;
  assign CLBLL_R_X71Y110_SLICE_X107Y110_B2 = 1'b1;
  assign CLBLL_R_X71Y110_SLICE_X107Y110_B3 = 1'b1;
  assign CLBLL_R_X71Y110_SLICE_X107Y110_B4 = 1'b1;
  assign CLBLL_R_X71Y110_SLICE_X107Y110_B5 = 1'b1;
  assign CLBLL_R_X71Y110_SLICE_X107Y110_B6 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_D6 = 1'b1;
  assign CLBLL_R_X71Y110_SLICE_X107Y110_C1 = 1'b1;
  assign CLBLL_R_X71Y110_SLICE_X107Y110_C2 = 1'b1;
  assign CLBLL_R_X71Y110_SLICE_X107Y110_C3 = 1'b1;
  assign CLBLL_R_X71Y110_SLICE_X107Y110_C4 = 1'b1;
  assign CLBLL_R_X71Y110_SLICE_X107Y110_C5 = 1'b1;
  assign CLBLL_R_X71Y110_SLICE_X107Y110_C6 = 1'b1;
  assign CLBLM_L_X70Y131_SLICE_X105Y131_A1 = 1'b1;
  assign CLBLM_L_X70Y131_SLICE_X105Y131_A2 = 1'b1;
  assign CLBLM_L_X70Y131_SLICE_X105Y131_A3 = 1'b1;
  assign CLBLM_L_X70Y131_SLICE_X105Y131_A4 = 1'b1;
  assign CLBLM_L_X70Y131_SLICE_X105Y131_A5 = 1'b1;
  assign CLBLM_L_X70Y131_SLICE_X105Y131_A6 = 1'b1;
  assign CLBLM_L_X70Y131_SLICE_X105Y131_B1 = 1'b1;
  assign CLBLL_R_X71Y110_SLICE_X107Y110_D1 = 1'b1;
  assign CLBLL_R_X71Y110_SLICE_X107Y110_D2 = 1'b1;
  assign CLBLL_R_X71Y110_SLICE_X107Y110_D3 = 1'b1;
  assign CLBLL_R_X71Y110_SLICE_X107Y110_D4 = 1'b1;
  assign CLBLL_R_X71Y110_SLICE_X107Y110_D5 = 1'b1;
  assign CLBLL_R_X71Y110_SLICE_X107Y110_D6 = 1'b1;
  assign CLBLM_L_X70Y131_SLICE_X105Y131_B2 = 1'b1;
  assign CLBLM_L_X70Y131_SLICE_X105Y131_B3 = 1'b1;
  assign CLBLM_L_X70Y131_SLICE_X105Y131_B4 = 1'b1;
  assign CLBLM_L_X70Y110_SLICE_X104Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X70Y131_SLICE_X105Y131_B6 = 1'b1;
  assign CLBLM_L_X70Y131_SLICE_X105Y131_C1 = 1'b1;
  assign CLBLM_L_X70Y131_SLICE_X105Y131_C2 = 1'b1;
  assign CLBLM_L_X70Y131_SLICE_X105Y131_C3 = 1'b1;
  assign CLBLM_L_X70Y131_SLICE_X105Y131_C4 = 1'b1;
  assign CLBLM_L_X70Y131_SLICE_X105Y131_C5 = 1'b1;
  assign CLBLM_L_X70Y131_SLICE_X105Y131_C6 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_A1 = 1'b1;
  assign CLBLM_L_X70Y131_SLICE_X105Y131_D1 = 1'b1;
  assign CLBLM_L_X70Y131_SLICE_X105Y131_D2 = 1'b1;
  assign CLBLM_L_X70Y131_SLICE_X105Y131_D3 = 1'b1;
  assign CLBLM_L_X70Y131_SLICE_X105Y131_D4 = 1'b1;
  assign CLBLM_L_X70Y131_SLICE_X105Y131_D5 = 1'b1;
  assign CLBLM_L_X70Y131_SLICE_X105Y131_D6 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_A2 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_A3 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_A4 = 1'b1;
  assign LIOI3_SING_X0Y50_OLOGIC_X0Y50_T1 = 1'b1;
  assign CLBLM_L_X70Y131_SLICE_X104Y131_A1 = CLBLM_L_X72Y133_SLICE_X109Y133_AO5;
  assign CLBLM_L_X70Y131_SLICE_X104Y131_A2 = CLBLM_L_X72Y132_SLICE_X109Y132_AO6;
  assign CLBLM_L_X70Y131_SLICE_X104Y131_A3 = CLBLM_L_X70Y131_SLICE_X104Y131_AQ;
  assign CLBLM_L_X70Y131_SLICE_X104Y131_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y131_SLICE_X104Y131_A5 = CLBLM_L_X70Y130_SLICE_X105Y130_AQ;
  assign CLBLM_L_X70Y131_SLICE_X104Y131_A6 = CLBLM_L_X70Y130_SLICE_X105Y130_A5Q;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_A5 = 1'b1;
  assign CLBLM_R_X67Y97_SLICE_X101Y97_B1 = CLBLM_R_X67Y98_SLICE_X101Y98_AO6;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_A6 = 1'b1;
  assign CLBLM_L_X70Y131_SLICE_X104Y131_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y131_SLICE_X104Y131_B2 = CLBLM_L_X70Y131_SLICE_X104Y131_BQ;
  assign CLBLM_L_X70Y131_SLICE_X104Y131_B3 = CLBLM_L_X70Y131_SLICE_X104Y131_AQ;
  assign CLBLM_L_X70Y131_SLICE_X104Y131_B4 = CLBLM_L_X72Y132_SLICE_X109Y132_AO6;
  assign CLBLM_L_X70Y131_SLICE_X104Y131_B5 = CLBLM_L_X70Y130_SLICE_X105Y130_AQ;
  assign CLBLM_L_X70Y131_SLICE_X104Y131_B6 = CLBLM_L_X70Y130_SLICE_X105Y130_A5Q;
  assign RIOB33_X105Y63_IOB_X1Y63_O = CLBLM_R_X103Y67_SLICE_X162Y67_AQ;
  assign CLBLM_L_X70Y131_SLICE_X104Y131_C1 = 1'b1;
  assign CLBLM_L_X70Y131_SLICE_X104Y131_C2 = 1'b1;
  assign CLBLM_L_X70Y131_SLICE_X104Y131_C3 = 1'b1;
  assign CLBLM_L_X70Y110_SLICE_X104Y110_D4 = 1'b1;
  assign CLBLM_L_X70Y131_SLICE_X104Y131_C4 = 1'b1;
  assign CLBLM_L_X70Y131_SLICE_X104Y131_C5 = 1'b1;
  assign CLBLM_L_X70Y131_SLICE_X104Y131_C6 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_AX = CLBLL_R_X77Y129_SLICE_X118Y129_AQ;
  assign CLBLM_L_X70Y110_SLICE_X104Y110_D5 = 1'b1;
  assign CLBLM_L_X70Y131_SLICE_X104Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X67Y97_SLICE_X101Y97_B2 = CLBLM_R_X67Y97_SLICE_X101Y97_BQ;
  assign CLBLM_L_X70Y131_SLICE_X104Y131_D1 = 1'b1;
  assign CLBLM_L_X70Y131_SLICE_X104Y131_D2 = 1'b1;
  assign CLBLM_L_X70Y131_SLICE_X104Y131_D3 = 1'b1;
  assign CLBLM_L_X70Y131_SLICE_X104Y131_D4 = 1'b1;
  assign CLBLM_L_X70Y131_SLICE_X104Y131_D5 = 1'b1;
  assign CLBLM_L_X70Y131_SLICE_X104Y131_D6 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_B1 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_B2 = 1'b1;
  assign CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_CE = 1'b1;
  assign CLBLM_L_X70Y131_SLICE_X104Y131_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_B3 = 1'b1;
  assign RIOI3_X105Y51_ILOGIC_X1Y52_D = RIOB33_X105Y51_IOB_X1Y52_I;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_B4 = 1'b1;
  assign CLBLM_R_X67Y97_SLICE_X101Y97_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign RIOI3_X105Y51_ILOGIC_X1Y51_D = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_B5 = 1'b1;
  assign CLBLM_R_X67Y115_SLICE_X101Y115_D3 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_B6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y57_ILOGIC_X1Y58_D = RIOB33_X105Y57_IOB_X1Y58_I;
  assign CLBLM_R_X67Y97_SLICE_X101Y97_B4 = CLBLM_R_X67Y98_SLICE_X101Y98_CO5;
  assign RIOI3_TBYTESRC_X105Y57_ILOGIC_X1Y57_D = RIOB33_X105Y57_IOB_X1Y57_I;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_C1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_T1 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_C2 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_C3 = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_D1 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_C4 = 1'b1;
  assign CLBLM_R_X67Y97_SLICE_X101Y97_B5 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_C5 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_C6 = 1'b1;
  assign CLBLM_R_X67Y97_SLICE_X101Y97_B6 = CLBLM_R_X67Y96_SLICE_X101Y96_BQ;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_D1 = CLBLL_R_X71Y110_SLICE_X106Y110_A5Q;
  assign CLBLM_L_X70Y131_SLICE_X105Y131_B5 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_T1 = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_T1 = 1'b1;
  assign CLBLL_R_X71Y111_SLICE_X106Y111_A1 = CLBLL_R_X71Y111_SLICE_X106Y111_DO6;
  assign CLBLL_R_X71Y111_SLICE_X106Y111_A2 = CLBLM_L_X72Y108_SLICE_X109Y108_A5Q;
  assign CLBLL_R_X71Y111_SLICE_X106Y111_A3 = CLBLL_R_X71Y111_SLICE_X106Y111_AQ;
  assign CLBLL_R_X71Y111_SLICE_X106Y111_A4 = CLBLL_R_X71Y112_SLICE_X106Y112_AQ;
  assign CLBLL_R_X71Y111_SLICE_X106Y111_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y111_SLICE_X106Y111_A6 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_D1 = 1'b1;
  assign CLBLM_L_X82Y130_SLICE_X129Y130_A1 = 1'b1;
  assign CLBLM_L_X82Y130_SLICE_X129Y130_A2 = 1'b1;
  assign CLBLL_R_X71Y111_SLICE_X106Y111_B1 = CLBLM_L_X70Y111_SLICE_X104Y111_AQ;
  assign CLBLL_R_X71Y111_SLICE_X106Y111_B2 = CLBLL_R_X71Y111_SLICE_X106Y111_BQ;
  assign CLBLL_R_X71Y111_SLICE_X106Y111_B3 = 1'b1;
  assign CLBLL_R_X71Y111_SLICE_X106Y111_B4 = CLBLM_L_X70Y111_SLICE_X104Y111_BO5;
  assign CLBLL_R_X71Y111_SLICE_X106Y111_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y111_SLICE_X106Y111_B6 = CLBLM_L_X70Y111_SLICE_X105Y111_BQ;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_D2 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_D3 = 1'b1;
  assign CLBLL_R_X71Y111_SLICE_X106Y111_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y111_SLICE_X106Y111_C2 = CLBLL_R_X71Y111_SLICE_X106Y111_CQ;
  assign CLBLL_R_X71Y111_SLICE_X106Y111_C3 = CLBLM_L_X70Y111_SLICE_X105Y111_BQ;
  assign CLBLL_R_X71Y111_SLICE_X106Y111_C4 = CLBLL_R_X71Y111_SLICE_X106Y111_BQ;
  assign CLBLL_R_X71Y111_SLICE_X106Y111_C5 = 1'b1;
  assign CLBLL_R_X71Y111_SLICE_X106Y111_C6 = CLBLM_L_X70Y111_SLICE_X104Y111_BO5;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_D4 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_D5 = 1'b1;
  assign CLBLL_R_X71Y111_SLICE_X106Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X82Y130_SLICE_X129Y130_C1 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_D6 = 1'b1;
  assign CLBLM_L_X82Y130_SLICE_X129Y130_C2 = 1'b1;
  assign CLBLM_L_X82Y130_SLICE_X129Y130_C4 = 1'b1;
  assign CLBLL_R_X71Y111_SLICE_X106Y111_D1 = CLBLL_R_X71Y111_SLICE_X107Y111_AQ;
  assign CLBLL_R_X71Y111_SLICE_X106Y111_D2 = CLBLL_R_X71Y111_SLICE_X107Y111_CO6;
  assign CLBLL_R_X71Y111_SLICE_X106Y111_D3 = CLBLM_L_X70Y112_SLICE_X104Y112_AQ;
  assign CLBLL_R_X71Y111_SLICE_X106Y111_D4 = CLBLM_L_X70Y111_SLICE_X104Y111_DO6;
  assign CLBLL_R_X71Y111_SLICE_X106Y111_D5 = CLBLM_L_X70Y112_SLICE_X104Y112_A5Q;
  assign CLBLL_R_X71Y111_SLICE_X106Y111_D6 = 1'b1;
  assign CLBLM_L_X82Y130_SLICE_X129Y130_D1 = 1'b1;
  assign CLBLL_R_X71Y111_SLICE_X106Y111_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X82Y130_SLICE_X129Y130_D2 = 1'b1;
  assign CLBLM_L_X82Y130_SLICE_X129Y130_D3 = 1'b1;
  assign CLBLM_L_X82Y130_SLICE_X129Y130_D4 = 1'b1;
  assign CLBLM_L_X82Y130_SLICE_X129Y130_D5 = 1'b1;
  assign CLBLM_L_X82Y130_SLICE_X129Y130_D6 = 1'b1;
  assign CLBLM_L_X82Y130_SLICE_X128Y130_A1 = 1'b1;
  assign CLBLM_L_X82Y130_SLICE_X128Y130_A2 = 1'b1;
  assign CLBLM_L_X82Y130_SLICE_X128Y130_A3 = 1'b1;
  assign CLBLM_L_X82Y130_SLICE_X128Y130_A4 = 1'b1;
  assign CLBLM_L_X82Y130_SLICE_X128Y130_A5 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X82Y130_SLICE_X128Y130_A6 = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_D1 = 1'b1;
  assign CLBLM_L_X82Y130_SLICE_X128Y130_AX = CLBLL_R_X77Y125_SLICE_X118Y125_AQ;
  assign CLBLM_L_X82Y130_SLICE_X128Y130_B1 = 1'b1;
  assign CLBLM_L_X82Y130_SLICE_X128Y130_B2 = 1'b1;
  assign CLBLM_L_X82Y130_SLICE_X128Y130_B3 = 1'b1;
  assign CLBLM_L_X82Y130_SLICE_X128Y130_B4 = 1'b1;
  assign CLBLM_L_X82Y130_SLICE_X128Y130_B5 = 1'b1;
  assign CLBLM_L_X82Y130_SLICE_X128Y130_B6 = 1'b1;
  assign CLBLL_R_X71Y111_SLICE_X107Y111_A1 = CLBLM_L_X72Y111_SLICE_X109Y111_CQ;
  assign CLBLL_R_X71Y111_SLICE_X107Y111_A2 = CLBLM_L_X72Y111_SLICE_X109Y111_A5Q;
  assign CLBLL_R_X71Y111_SLICE_X107Y111_A3 = CLBLM_L_X72Y111_SLICE_X109Y111_AQ;
  assign CLBLL_R_X71Y111_SLICE_X107Y111_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y111_SLICE_X107Y111_A5 = CLBLM_L_X70Y111_SLICE_X104Y111_BQ;
  assign CLBLL_R_X71Y111_SLICE_X107Y111_A6 = CLBLL_R_X71Y111_SLICE_X107Y111_AQ;
  assign CLBLM_L_X82Y130_SLICE_X128Y130_C5 = 1'b1;
  assign CLBLM_L_X82Y130_SLICE_X128Y130_C6 = 1'b1;
  assign CLBLL_R_X71Y111_SLICE_X107Y111_B1 = CLBLL_R_X71Y111_SLICE_X107Y111_DO6;
  assign CLBLL_R_X71Y111_SLICE_X107Y111_B2 = CLBLM_L_X70Y111_SLICE_X105Y111_AQ;
  assign CLBLL_R_X71Y111_SLICE_X107Y111_B3 = CLBLL_R_X71Y111_SLICE_X107Y111_AQ;
  assign CLBLL_R_X71Y111_SLICE_X107Y111_B4 = CLBLL_R_X71Y111_SLICE_X106Y111_BQ;
  assign CLBLL_R_X71Y111_SLICE_X107Y111_B5 = CLBLM_L_X72Y111_SLICE_X108Y111_AO6;
  assign CLBLL_R_X71Y111_SLICE_X107Y111_B6 = CLBLM_L_X70Y111_SLICE_X104Y111_AQ;
  assign CLBLM_L_X82Y130_SLICE_X128Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X82Y130_SLICE_X128Y130_D1 = 1'b1;
  assign CLBLL_R_X71Y111_SLICE_X107Y111_C1 = CLBLL_R_X71Y111_SLICE_X106Y111_CQ;
  assign CLBLL_R_X71Y111_SLICE_X107Y111_C2 = CLBLM_L_X70Y111_SLICE_X105Y111_AQ;
  assign CLBLL_R_X71Y111_SLICE_X107Y111_C3 = CLBLM_L_X70Y111_SLICE_X104Y111_AQ;
  assign CLBLL_R_X71Y111_SLICE_X107Y111_C4 = CLBLM_L_X70Y111_SLICE_X105Y111_BQ;
  assign CLBLL_R_X71Y111_SLICE_X107Y111_C5 = 1'b1;
  assign CLBLL_R_X71Y111_SLICE_X107Y111_C6 = CLBLL_R_X71Y111_SLICE_X106Y111_BQ;
  assign CLBLM_L_X82Y130_SLICE_X128Y130_D2 = 1'b1;
  assign CLBLM_L_X82Y130_SLICE_X128Y130_D3 = 1'b1;
  assign CLBLL_R_X71Y111_SLICE_X107Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X70Y132_SLICE_X105Y132_A1 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X105Y132_A2 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X105Y132_A3 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X105Y132_A4 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X105Y132_A5 = 1'b1;
  assign CLBLL_R_X71Y111_SLICE_X107Y111_D1 = 1'b1;
  assign CLBLL_R_X71Y111_SLICE_X107Y111_D2 = CLBLM_L_X70Y111_SLICE_X105Y111_BQ;
  assign CLBLL_R_X71Y111_SLICE_X107Y111_D3 = CLBLM_L_X70Y112_SLICE_X104Y112_A5Q;
  assign CLBLL_R_X71Y111_SLICE_X107Y111_D4 = CLBLL_R_X71Y111_SLICE_X106Y111_CQ;
  assign CLBLL_R_X71Y111_SLICE_X107Y111_D5 = CLBLM_L_X70Y112_SLICE_X104Y112_AQ;
  assign CLBLL_R_X71Y111_SLICE_X107Y111_D6 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X105Y132_A6 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X105Y132_AX = CLBLM_L_X70Y135_SLICE_X105Y135_AQ;
  assign CLBLL_R_X71Y111_SLICE_X107Y111_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X70Y132_SLICE_X105Y132_B1 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X105Y132_B2 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X105Y132_B3 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X105Y132_B4 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X105Y132_B5 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X105Y132_B6 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X105Y132_BX = CLBLM_L_X70Y133_SLICE_X104Y133_A5Q;
  assign CLBLM_L_X70Y132_SLICE_X105Y132_C1 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X105Y132_C2 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X105Y132_C3 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X105Y132_C4 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X105Y132_C5 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X105Y132_C6 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X105Y132_CE = CLBLM_L_X76Y109_SLICE_X116Y109_AO6;
  assign CLBLM_L_X70Y132_SLICE_X105Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X70Y132_SLICE_X105Y132_D1 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X105Y132_D2 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X105Y132_D3 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X105Y132_D4 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X105Y132_D5 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X105Y132_D6 = 1'b1;
  assign RIOB33_X105Y65_IOB_X1Y65_O = CLBLM_R_X103Y67_SLICE_X162Y67_BQ;
  assign RIOB33_X105Y65_IOB_X1Y66_O = CLBLM_R_X103Y67_SLICE_X162Y67_CQ;
  assign CLBLM_L_X70Y132_SLICE_X105Y132_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X70Y132_SLICE_X104Y132_A1 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X104Y132_A2 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X104Y132_A3 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X104Y132_A4 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X104Y132_A5 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X104Y132_A6 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X104Y132_B1 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X104Y132_B2 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X104Y132_B3 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X104Y132_B4 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X104Y132_B5 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X104Y132_B6 = 1'b1;
  assign CLBLM_R_X67Y115_SLICE_X101Y115_D5 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X104Y132_C1 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X104Y132_C2 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X104Y132_C3 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X104Y132_C4 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X104Y132_C5 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X104Y132_C6 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_B3 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X104Y132_D1 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X104Y132_D2 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X104Y132_D3 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X104Y132_D4 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X104Y132_D5 = 1'b1;
  assign CLBLM_L_X70Y132_SLICE_X104Y132_D6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1 = 1'b1;
  assign CLBLM_R_X67Y115_SLICE_X101Y115_D6 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_B4 = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_T1 = 1'b1;
  assign CLBLL_R_X71Y112_SLICE_X106Y112_A1 = CLBLL_R_X71Y111_SLICE_X107Y111_CO6;
  assign CLBLL_R_X71Y112_SLICE_X106Y112_A2 = CLBLM_L_X70Y112_SLICE_X104Y112_A5Q;
  assign CLBLL_R_X71Y112_SLICE_X106Y112_A3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y112_SLICE_X106Y112_A4 = CLBLM_L_X70Y112_SLICE_X104Y112_AQ;
  assign CLBLL_R_X71Y112_SLICE_X106Y112_A5 = CLBLM_L_X72Y111_SLICE_X108Y111_AO6;
  assign CLBLL_R_X71Y112_SLICE_X106Y112_A6 = CLBLL_R_X71Y111_SLICE_X107Y111_AQ;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_B4 = CLBLM_L_X76Y126_SLICE_X117Y126_AQ;
  assign CLBLM_R_X67Y111_SLICE_X101Y111_B4 = CLBLM_R_X67Y111_SLICE_X101Y111_B5Q;
  assign CLBLL_R_X71Y112_SLICE_X106Y112_B1 = CLBLM_L_X70Y112_SLICE_X105Y112_A5Q;
  assign CLBLL_R_X71Y112_SLICE_X106Y112_B2 = CLBLL_R_X71Y112_SLICE_X106Y112_BQ;
  assign CLBLL_R_X71Y112_SLICE_X106Y112_B3 = CLBLL_R_X71Y112_SLICE_X106Y112_B5Q;
  assign CLBLL_R_X71Y112_SLICE_X106Y112_B4 = CLBLM_L_X72Y111_SLICE_X109Y111_CQ;
  assign CLBLL_R_X71Y112_SLICE_X106Y112_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y112_SLICE_X106Y112_B6 = 1'b1;
  assign CLBLM_R_X67Y111_SLICE_X101Y111_B5 = 1'b1;
  assign CLBLM_R_X67Y111_SLICE_X101Y111_B6 = 1'b1;
  assign CLBLL_R_X71Y112_SLICE_X106Y112_C1 = 1'b1;
  assign CLBLL_R_X71Y112_SLICE_X106Y112_C2 = 1'b1;
  assign CLBLL_R_X71Y112_SLICE_X106Y112_C3 = 1'b1;
  assign CLBLL_R_X71Y112_SLICE_X106Y112_C4 = 1'b1;
  assign CLBLL_R_X71Y112_SLICE_X106Y112_C5 = 1'b1;
  assign CLBLL_R_X71Y112_SLICE_X106Y112_C6 = 1'b1;
  assign CLBLL_R_X71Y112_SLICE_X106Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X71Y112_SLICE_X106Y112_D1 = 1'b1;
  assign CLBLL_R_X71Y112_SLICE_X106Y112_D2 = 1'b1;
  assign CLBLL_R_X71Y112_SLICE_X106Y112_D3 = 1'b1;
  assign CLBLL_R_X71Y112_SLICE_X106Y112_D4 = 1'b1;
  assign CLBLL_R_X71Y112_SLICE_X106Y112_D5 = 1'b1;
  assign CLBLL_R_X71Y112_SLICE_X106Y112_D6 = 1'b1;
  assign CLBLL_R_X71Y112_SLICE_X106Y112_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X67Y111_SLICE_X101Y111_C1 = CLBLM_R_X67Y111_SLICE_X101Y111_B5Q;
  assign CLBLM_R_X67Y111_SLICE_X101Y111_C2 = 1'b1;
  assign CLBLM_R_X67Y111_SLICE_X101Y111_C3 = CLBLM_R_X67Y111_SLICE_X101Y111_BQ;
  assign CLBLM_R_X67Y111_SLICE_X101Y111_C4 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_D1 = 1'b1;
  assign CLBLM_R_X67Y111_SLICE_X101Y111_C5 = CLBLM_R_X67Y111_SLICE_X101Y111_AQ;
  assign CLBLL_R_X71Y112_SLICE_X107Y112_A1 = 1'b1;
  assign CLBLL_R_X71Y112_SLICE_X107Y112_A2 = 1'b1;
  assign CLBLL_R_X71Y112_SLICE_X107Y112_A3 = 1'b1;
  assign CLBLL_R_X71Y112_SLICE_X107Y112_A4 = 1'b1;
  assign CLBLL_R_X71Y112_SLICE_X107Y112_A5 = 1'b1;
  assign CLBLL_R_X71Y112_SLICE_X107Y112_A6 = 1'b1;
  assign CLBLM_R_X67Y111_SLICE_X101Y111_C6 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_T1 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_D1 = CLBLL_R_X73Y119_SLICE_X110Y119_AQ;
  assign CLBLL_R_X71Y112_SLICE_X107Y112_B1 = 1'b1;
  assign CLBLL_R_X71Y112_SLICE_X107Y112_B2 = 1'b1;
  assign CLBLL_R_X71Y112_SLICE_X107Y112_B3 = 1'b1;
  assign CLBLL_R_X71Y112_SLICE_X107Y112_B4 = 1'b1;
  assign CLBLL_R_X71Y112_SLICE_X107Y112_B5 = 1'b1;
  assign CLBLL_R_X71Y112_SLICE_X107Y112_B6 = 1'b1;
  assign CLBLM_R_X67Y111_SLICE_X101Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_D1 = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign CLBLL_R_X71Y112_SLICE_X107Y112_C1 = 1'b1;
  assign CLBLL_R_X71Y112_SLICE_X107Y112_C2 = 1'b1;
  assign CLBLL_R_X71Y112_SLICE_X107Y112_C3 = 1'b1;
  assign CLBLL_R_X71Y112_SLICE_X107Y112_C4 = 1'b1;
  assign CLBLL_R_X71Y112_SLICE_X107Y112_C5 = 1'b1;
  assign CLBLL_R_X71Y112_SLICE_X107Y112_C6 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_T1 = 1'b1;
  assign CLBLM_L_X70Y133_SLICE_X105Y133_A1 = CLBLM_L_X70Y133_SLICE_X104Y133_A5Q;
  assign CLBLL_R_X71Y112_SLICE_X107Y112_D1 = 1'b1;
  assign CLBLL_R_X71Y112_SLICE_X107Y112_D2 = 1'b1;
  assign CLBLL_R_X71Y112_SLICE_X107Y112_D3 = 1'b1;
  assign CLBLL_R_X71Y112_SLICE_X107Y112_D4 = 1'b1;
  assign CLBLL_R_X71Y112_SLICE_X107Y112_D5 = 1'b1;
  assign CLBLL_R_X71Y112_SLICE_X107Y112_D6 = 1'b1;
  assign CLBLM_L_X70Y133_SLICE_X105Y133_A4 = CLBLM_L_X70Y132_SLICE_X105Y132_BQ;
  assign CLBLM_L_X70Y133_SLICE_X105Y133_A5 = CLBLM_L_X70Y124_SLICE_X105Y124_AO6;
  assign CLBLM_L_X70Y133_SLICE_X105Y133_A6 = 1'b1;
  assign CLBLM_L_X70Y133_SLICE_X105Y133_B1 = 1'b1;
  assign CLBLM_L_X70Y133_SLICE_X105Y133_B2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y133_SLICE_X105Y133_B3 = CLBLM_L_X70Y133_SLICE_X105Y133_AQ;
  assign CLBLM_L_X70Y133_SLICE_X105Y133_B4 = CLBLM_L_X70Y133_SLICE_X104Y133_DO6;
  assign CLBLM_L_X70Y133_SLICE_X105Y133_B5 = CLBLM_L_X70Y124_SLICE_X105Y124_AO6;
  assign CLBLM_L_X70Y133_SLICE_X105Y133_B6 = CLBLM_L_X70Y133_SLICE_X105Y133_BQ;
  assign CLBLM_L_X70Y133_SLICE_X105Y133_C1 = CLBLM_L_X70Y124_SLICE_X105Y124_AO6;
  assign CLBLM_L_X70Y133_SLICE_X105Y133_C2 = CLBLM_L_X70Y133_SLICE_X105Y133_CQ;
  assign CLBLM_L_X70Y133_SLICE_X105Y133_C3 = CLBLM_L_X70Y133_SLICE_X105Y133_BQ;
  assign CLBLM_L_X70Y133_SLICE_X105Y133_C4 = CLBLM_L_X70Y133_SLICE_X104Y133_AQ;
  assign CLBLM_L_X70Y133_SLICE_X105Y133_C5 = CLBLM_L_X70Y133_SLICE_X104Y133_A5Q;
  assign CLBLM_L_X70Y133_SLICE_X105Y133_C6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_B5 = 1'b1;
  assign CLBLM_R_X67Y111_SLICE_X101Y111_D2 = 1'b1;
  assign CLBLM_L_X70Y133_SLICE_X105Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X67Y111_SLICE_X101Y111_D3 = CLBLM_R_X67Y111_SLICE_X101Y111_BQ;
  assign CLBLM_R_X67Y111_SLICE_X101Y111_D4 = CLBLM_R_X67Y111_SLICE_X101Y111_AQ;
  assign CLBLM_L_X70Y133_SLICE_X105Y133_D1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y133_SLICE_X105Y133_D2 = CLBLM_L_X70Y133_SLICE_X105Y133_CQ;
  assign CLBLM_L_X70Y133_SLICE_X105Y133_D3 = CLBLM_L_X70Y133_SLICE_X105Y133_DQ;
  assign CLBLM_L_X70Y133_SLICE_X105Y133_D4 = CLBLM_L_X70Y133_SLICE_X104Y133_CO5;
  assign CLBLM_L_X70Y133_SLICE_X105Y133_D5 = 1'b1;
  assign CLBLM_L_X70Y133_SLICE_X105Y133_D6 = CLBLM_L_X70Y134_SLICE_X105Y134_CQ;
  assign CLBLM_R_X67Y111_SLICE_X101Y111_D5 = 1'b1;
  assign CLBLM_R_X67Y111_SLICE_X101Y111_D6 = 1'b1;
  assign CLBLM_L_X70Y133_SLICE_X105Y133_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_D1 = CLBLM_L_X82Y98_SLICE_X128Y98_AQ;
  assign CLBLM_L_X70Y133_SLICE_X104Y133_A1 = CLBLM_L_X70Y133_SLICE_X104Y133_AQ;
  assign CLBLM_L_X70Y133_SLICE_X104Y133_A2 = CLBLM_L_X70Y133_SLICE_X104Y133_BQ;
  assign CLBLM_L_X70Y133_SLICE_X104Y133_A3 = CLBLM_L_X70Y124_SLICE_X105Y124_AO6;
  assign CLBLM_L_X70Y133_SLICE_X104Y133_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y133_SLICE_X104Y133_A5 = CLBLM_L_X70Y133_SLICE_X105Y133_AQ;
  assign CLBLM_L_X70Y133_SLICE_X104Y133_A6 = CLBLM_L_X70Y133_SLICE_X104Y133_A5Q;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_T1 = 1'b1;
  assign CLBLM_L_X70Y133_SLICE_X104Y133_AX = CLBLM_L_X70Y133_SLICE_X104Y133_CO6;
  assign CLBLM_L_X70Y133_SLICE_X104Y133_B1 = CLBLL_R_X71Y133_SLICE_X106Y133_AO6;
  assign CLBLM_L_X70Y133_SLICE_X104Y133_B2 = CLBLM_L_X70Y133_SLICE_X104Y133_BQ;
  assign CLBLM_L_X70Y133_SLICE_X104Y133_B3 = CLBLM_L_X70Y124_SLICE_X105Y124_AO6;
  assign CLBLM_L_X70Y133_SLICE_X104Y133_B4 = CLBLM_L_X70Y134_SLICE_X104Y134_CO5;
  assign CLBLM_L_X70Y133_SLICE_X104Y133_B5 = CLBLM_L_X70Y134_SLICE_X104Y134_AQ;
  assign CLBLM_L_X70Y133_SLICE_X104Y133_B6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y111_SLICE_X101Y111_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_D1 = CLBLM_R_X103Y69_SLICE_X163Y69_AQ;
  assign CLBLM_L_X70Y133_SLICE_X104Y133_C1 = CLBLM_L_X70Y124_SLICE_X105Y124_AO6;
  assign CLBLM_L_X70Y133_SLICE_X104Y133_C2 = CLBLM_L_X70Y133_SLICE_X104Y133_AQ;
  assign CLBLM_L_X70Y133_SLICE_X104Y133_C3 = CLBLM_L_X70Y133_SLICE_X104Y133_A5Q;
  assign CLBLM_L_X70Y133_SLICE_X104Y133_C4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y133_SLICE_X104Y133_C5 = 1'b1;
  assign CLBLM_L_X70Y133_SLICE_X104Y133_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_T1 = 1'b1;
  assign CLBLM_L_X70Y133_SLICE_X104Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X70Y133_SLICE_X104Y133_D1 = CLBLM_L_X70Y133_SLICE_X105Y133_AQ;
  assign CLBLM_L_X70Y133_SLICE_X104Y133_D2 = CLBLM_L_X70Y133_SLICE_X104Y133_AQ;
  assign CLBLM_L_X70Y133_SLICE_X104Y133_D3 = CLBLM_L_X70Y134_SLICE_X104Y134_DO6;
  assign CLBLM_L_X70Y133_SLICE_X104Y133_D4 = CLBLM_L_X70Y134_SLICE_X104Y134_CO6;
  assign CLBLM_L_X70Y133_SLICE_X104Y133_D5 = CLBLM_L_X70Y134_SLICE_X104Y134_AQ;
  assign CLBLM_L_X70Y133_SLICE_X104Y133_D6 = CLBLM_L_X70Y134_SLICE_X105Y134_BQ;
  assign CLBLM_L_X70Y133_SLICE_X104Y133_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_A2 = CLBLM_R_X67Y100_SLICE_X100Y100_BQ;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_A3 = 1'b1;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_A4 = CLBLM_R_X67Y99_SLICE_X100Y99_AQ;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_A5 = CLBLM_R_X67Y99_SLICE_X100Y99_BQ;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_A6 = CLBLM_R_X67Y100_SLICE_X100Y100_CQ;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_B1 = CLBLM_R_X67Y100_SLICE_X100Y100_CQ;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_B2 = CLBLM_R_X67Y103_SLICE_X100Y103_BQ;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_B3 = CLBLM_R_X65Y99_SLICE_X99Y99_AQ;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_B4 = CLBLM_R_X67Y99_SLICE_X100Y99_AQ;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_B5 = CLBLM_R_X67Y99_SLICE_X100Y99_BQ;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_B6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_C2 = CLBLM_R_X65Y99_SLICE_X99Y99_CQ;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_C3 = CLBLM_R_X65Y99_SLICE_X99Y99_DQ;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_C4 = CLBLM_R_X65Y99_SLICE_X99Y99_BQ;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_C5 = CLBLM_R_X65Y99_SLICE_X99Y99_AQ;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_C6 = 1'b1;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_D1 = CLBLM_R_X65Y99_SLICE_X99Y99_C5Q;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_D2 = CLBLM_R_X65Y99_SLICE_X99Y99_CQ;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_D3 = CLBLM_R_X65Y99_SLICE_X99Y99_DQ;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_D4 = CLBLM_R_X65Y99_SLICE_X99Y99_BQ;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_D5 = CLBLM_R_X65Y99_SLICE_X99Y99_AQ;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_D6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_A1 = CLBLM_R_X63Y98_SLICE_X95Y98_AO6;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_B6 = CLBLL_R_X77Y127_SLICE_X119Y127_AO5;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_A2 = CLBLM_R_X65Y99_SLICE_X98Y99_BQ;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_A3 = CLBLM_R_X65Y99_SLICE_X98Y99_AQ;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_A5 = 1'b1;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_A6 = CLBLM_R_X63Y99_SLICE_X95Y99_AO5;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_B1 = CLBLM_L_X64Y99_SLICE_X96Y99_A5Q;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_B2 = CLBLM_R_X65Y99_SLICE_X98Y99_BQ;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_B3 = CLBLM_R_X65Y99_SLICE_X98Y99_CQ;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_B4 = CLBLM_R_X63Y99_SLICE_X94Y99_A5Q;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_B5 = CLBLM_L_X64Y99_SLICE_X96Y99_BQ;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_B6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y111_SLICE_X100Y111_B6 = CLBLM_R_X67Y111_SLICE_X100Y111_A5Q;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_C1 = CLBLM_L_X64Y99_SLICE_X96Y99_BQ;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_C2 = CLBLM_R_X65Y99_SLICE_X98Y99_CQ;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_C3 = CLBLL_R_X79Y99_SLICE_X122Y99_AO6;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_C4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_C5 = CLBLM_L_X64Y99_SLICE_X96Y99_A5Q;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_C6 = CLBLM_R_X63Y99_SLICE_X94Y99_A5Q;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_D1 = 1'b1;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_D2 = 1'b1;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_D3 = 1'b1;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_D4 = 1'b1;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_D5 = 1'b1;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_D6 = 1'b1;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_A5 = CLBLM_L_X72Y127_SLICE_X108Y127_AQ;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_A6 = CLBLM_L_X72Y127_SLICE_X108Y127_A5Q;
  assign RIOI3_X105Y53_ILOGIC_X1Y54_D = RIOB33_X105Y53_IOB_X1Y54_I;
  assign CLBLM_R_X67Y111_SLICE_X100Y111_C5 = 1'b1;
  assign RIOI3_X105Y53_ILOGIC_X1Y53_D = RIOB33_X105Y53_IOB_X1Y53_I;
  assign CLBLM_R_X67Y111_SLICE_X100Y111_C6 = 1'b1;
  assign CLBLM_R_X67Y111_SLICE_X100Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_B4 = CLBLL_R_X75Y127_SLICE_X115Y127_DQ;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_B5 = 1'b1;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_B6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_D1 = 1'b1;
  assign CLBLM_R_X67Y111_SLICE_X100Y111_D4 = 1'b1;
  assign RIOB33_X105Y69_IOB_X1Y70_O = CLBLM_L_X82Y98_SLICE_X128Y98_AQ;
  assign RIOB33_X105Y69_IOB_X1Y69_O = CLBLM_R_X103Y69_SLICE_X163Y69_AQ;
  assign CLBLM_R_X67Y111_SLICE_X100Y111_D5 = 1'b1;
  assign CLBLM_L_X70Y134_SLICE_X105Y134_A1 = CLBLL_R_X71Y133_SLICE_X106Y133_AQ;
  assign CLBLM_L_X70Y134_SLICE_X105Y134_A2 = CLBLM_L_X70Y134_SLICE_X105Y134_BQ;
  assign CLBLM_L_X70Y134_SLICE_X105Y134_A3 = CLBLM_L_X70Y134_SLICE_X105Y134_AQ;
  assign CLBLM_L_X70Y134_SLICE_X105Y134_A4 = CLBLM_L_X70Y134_SLICE_X105Y134_DO5;
  assign CLBLM_L_X70Y134_SLICE_X105Y134_A5 = CLBLM_L_X72Y134_SLICE_X109Y134_AO6;
  assign CLBLM_L_X70Y134_SLICE_X105Y134_A6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_T1 = 1'b1;
  assign CLBLM_L_X70Y134_SLICE_X105Y134_B1 = CLBLM_L_X70Y134_SLICE_X105Y134_DO6;
  assign CLBLM_L_X70Y134_SLICE_X105Y134_B2 = CLBLM_L_X70Y134_SLICE_X105Y134_BQ;
  assign CLBLM_L_X70Y134_SLICE_X105Y134_B3 = CLBLM_L_X70Y134_SLICE_X105Y134_CQ;
  assign CLBLM_L_X70Y134_SLICE_X105Y134_B4 = CLBLM_L_X72Y134_SLICE_X109Y134_AO6;
  assign CLBLM_L_X70Y134_SLICE_X105Y134_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y134_SLICE_X105Y134_B6 = 1'b1;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X70Y134_SLICE_X105Y134_C1 = CLBLM_L_X70Y135_SLICE_X105Y135_AQ;
  assign CLBLM_L_X70Y134_SLICE_X105Y134_C2 = CLBLM_L_X70Y135_SLICE_X105Y135_A5Q;
  assign CLBLM_L_X70Y134_SLICE_X105Y134_C3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y134_SLICE_X105Y134_C4 = CLBLL_R_X71Y134_SLICE_X106Y134_BQ;
  assign CLBLM_L_X64Y122_SLICE_X97Y122_A1 = 1'b1;
  assign CLBLM_L_X64Y122_SLICE_X97Y122_A2 = 1'b1;
  assign CLBLM_L_X64Y122_SLICE_X97Y122_A3 = 1'b1;
  assign CLBLM_L_X64Y122_SLICE_X97Y122_A4 = 1'b1;
  assign CLBLM_L_X64Y122_SLICE_X97Y122_A5 = 1'b1;
  assign CLBLM_L_X64Y122_SLICE_X97Y122_A6 = 1'b1;
  assign CLBLM_L_X70Y134_SLICE_X105Y134_C5 = CLBLM_L_X72Y133_SLICE_X109Y133_CO6;
  assign CLBLM_L_X70Y134_SLICE_X105Y134_C6 = CLBLM_L_X70Y134_SLICE_X105Y134_CQ;
  assign CLBLM_L_X70Y134_SLICE_X105Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X64Y122_SLICE_X97Y122_B1 = 1'b1;
  assign CLBLM_L_X64Y122_SLICE_X97Y122_B2 = 1'b1;
  assign CLBLM_L_X70Y134_SLICE_X105Y134_D2 = CLBLM_L_X70Y135_SLICE_X105Y135_A5Q;
  assign CLBLM_L_X70Y134_SLICE_X105Y134_D3 = 1'b1;
  assign CLBLM_L_X64Y122_SLICE_X97Y122_B4 = 1'b1;
  assign CLBLM_L_X64Y122_SLICE_X97Y122_B5 = 1'b1;
  assign CLBLM_L_X64Y122_SLICE_X97Y122_B3 = 1'b1;
  assign CLBLM_L_X64Y122_SLICE_X97Y122_B6 = 1'b1;
  assign CLBLM_L_X70Y134_SLICE_X105Y134_D1 = CLBLM_L_X70Y135_SLICE_X105Y135_AQ;
  assign CLBLM_L_X64Y122_SLICE_X97Y122_C1 = 1'b1;
  assign CLBLM_L_X64Y122_SLICE_X97Y122_C2 = 1'b1;
  assign CLBLM_L_X64Y122_SLICE_X97Y122_C3 = 1'b1;
  assign CLBLM_L_X64Y122_SLICE_X97Y122_C4 = 1'b1;
  assign CLBLM_L_X64Y122_SLICE_X97Y122_C5 = 1'b1;
  assign CLBLM_L_X70Y134_SLICE_X104Y134_A2 = CLBLM_L_X70Y134_SLICE_X105Y134_DO5;
  assign CLBLM_L_X64Y122_SLICE_X97Y122_C6 = 1'b1;
  assign CLBLM_L_X70Y134_SLICE_X104Y134_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y134_SLICE_X105Y134_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X70Y134_SLICE_X104Y134_A1 = CLBLM_L_X70Y134_SLICE_X104Y134_BQ;
  assign CLBLM_L_X70Y134_SLICE_X104Y134_A3 = CLBLM_L_X70Y134_SLICE_X104Y134_AQ;
  assign CLBLM_L_X70Y134_SLICE_X104Y134_A5 = CLBLM_L_X72Y134_SLICE_X109Y134_AO6;
  assign CLBLM_L_X70Y134_SLICE_X104Y134_A6 = CLBLM_L_X70Y135_SLICE_X105Y135_A5Q;
  assign CLBLM_L_X64Y122_SLICE_X97Y122_D1 = 1'b1;
  assign CLBLM_L_X64Y122_SLICE_X97Y122_D2 = 1'b1;
  assign CLBLM_L_X64Y122_SLICE_X97Y122_D3 = 1'b1;
  assign CLBLM_L_X64Y122_SLICE_X97Y122_D4 = 1'b1;
  assign CLBLM_L_X70Y134_SLICE_X104Y134_B5 = CLBLL_R_X71Y133_SLICE_X106Y133_AO6;
  assign CLBLM_L_X70Y134_SLICE_X104Y134_B6 = CLBLM_L_X72Y133_SLICE_X109Y133_CO6;
  assign CLBLM_L_X64Y122_SLICE_X97Y122_D5 = 1'b1;
  assign CLBLM_L_X64Y122_SLICE_X97Y122_D6 = 1'b1;
  assign CLBLM_L_X70Y134_SLICE_X104Y134_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y134_SLICE_X104Y134_B2 = CLBLM_L_X70Y134_SLICE_X104Y134_BQ;
  assign CLBLM_L_X70Y134_SLICE_X104Y134_C1 = CLBLM_L_X70Y134_SLICE_X105Y134_AQ;
  assign CLBLM_L_X70Y134_SLICE_X104Y134_B4 = CLBLM_L_X70Y135_SLICE_X104Y135_BQ;
  assign CLBLM_L_X64Y122_SLICE_X96Y122_A1 = 1'b1;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_A4 = CLBLM_L_X62Y107_SLICE_X93Y107_BQ;
  assign CLBLM_L_X64Y122_SLICE_X96Y122_A2 = 1'b1;
  assign CLBLM_L_X64Y122_SLICE_X96Y122_A3 = 1'b1;
  assign CLBLM_L_X64Y122_SLICE_X96Y122_A4 = 1'b1;
  assign CLBLM_L_X64Y122_SLICE_X96Y122_A5 = 1'b1;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_A5 = CLBLM_R_X63Y106_SLICE_X95Y106_BQ;
  assign CLBLM_L_X64Y122_SLICE_X96Y122_A6 = 1'b1;
  assign CLBLM_L_X70Y134_SLICE_X104Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X64Y122_SLICE_X96Y122_AX = CLBLM_L_X68Y121_SLICE_X102Y121_AQ;
  assign CLBLM_L_X70Y134_SLICE_X104Y134_C4 = CLBLM_L_X70Y133_SLICE_X104Y133_AQ;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_A6 = 1'b1;
  assign CLBLM_L_X64Y122_SLICE_X96Y122_B1 = 1'b1;
  assign CLBLM_L_X64Y122_SLICE_X96Y122_B2 = 1'b1;
  assign CLBLM_L_X64Y122_SLICE_X96Y122_B3 = 1'b1;
  assign CLBLM_L_X64Y122_SLICE_X96Y122_B4 = 1'b1;
  assign CLBLM_L_X64Y122_SLICE_X96Y122_B5 = 1'b1;
  assign CLBLM_L_X64Y122_SLICE_X96Y122_B6 = 1'b1;
  assign CLBLM_L_X70Y134_SLICE_X104Y134_D1 = CLBLM_L_X70Y133_SLICE_X104Y133_A5Q;
  assign CLBLM_L_X70Y134_SLICE_X104Y134_D2 = CLBLM_L_X70Y133_SLICE_X105Y133_AQ;
  assign CLBLM_L_X64Y122_SLICE_X96Y122_C1 = 1'b1;
  assign CLBLM_L_X64Y122_SLICE_X96Y122_C2 = 1'b1;
  assign CLBLM_L_X64Y122_SLICE_X96Y122_C3 = 1'b1;
  assign CLBLM_L_X64Y122_SLICE_X96Y122_C4 = 1'b1;
  assign CLBLM_L_X64Y122_SLICE_X96Y122_C5 = 1'b1;
  assign CLBLM_L_X64Y122_SLICE_X96Y122_C6 = 1'b1;
  assign CLBLM_L_X64Y122_SLICE_X96Y122_CE = CLBLM_L_X76Y109_SLICE_X116Y109_AO6;
  assign CLBLM_L_X70Y134_SLICE_X104Y134_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X64Y122_SLICE_X96Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_A1 = CLBLM_R_X63Y99_SLICE_X95Y99_AO5;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_A3 = CLBLM_R_X65Y100_SLICE_X99Y100_AQ;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_A4 = CLBLM_R_X65Y100_SLICE_X98Y100_BQ;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_A5 = CLBLM_R_X65Y100_SLICE_X99Y100_A5Q;
  assign CLBLM_L_X64Y122_SLICE_X96Y122_D1 = 1'b1;
  assign CLBLM_L_X64Y122_SLICE_X96Y122_D2 = 1'b1;
  assign CLBLM_L_X64Y122_SLICE_X96Y122_D3 = 1'b1;
  assign CLBLM_L_X64Y122_SLICE_X96Y122_D4 = 1'b1;
  assign CLBLM_L_X64Y122_SLICE_X96Y122_D5 = 1'b1;
  assign CLBLM_L_X64Y122_SLICE_X96Y122_D6 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_B5 = CLBLM_R_X63Y99_SLICE_X94Y99_A5Q;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_B6 = CLBLM_R_X65Y100_SLICE_X99Y100_BQ;
  assign CLBLM_L_X64Y122_SLICE_X96Y122_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_C1 = CLBLM_R_X65Y101_SLICE_X99Y101_AQ;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_C2 = CLBLM_R_X65Y100_SLICE_X99Y100_CQ;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_C3 = CLBLM_L_X64Y99_SLICE_X96Y99_BO5;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_C4 = CLBLM_R_X65Y100_SLICE_X99Y100_BQ;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_C5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_C6 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_T1 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_B6 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_D1 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_D2 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_D3 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_D4 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_D5 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_D6 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_C1 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_A1 = CLBLM_R_X63Y99_SLICE_X95Y99_AO5;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_A2 = CLBLM_R_X65Y99_SLICE_X98Y99_AQ;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_A3 = CLBLM_R_X65Y100_SLICE_X98Y100_AQ;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_C2 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_A5 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_A6 = CLBLM_R_X65Y99_SLICE_X98Y99_BQ;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_B2 = CLBLM_R_X65Y100_SLICE_X98Y100_BQ;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_C4 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_B3 = CLBLM_R_X65Y100_SLICE_X98Y100_AQ;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_B4 = CLBLM_L_X64Y99_SLICE_X96Y99_A5Q;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_B5 = CLBLM_R_X63Y99_SLICE_X94Y99_A5Q;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_B6 = CLBLM_L_X64Y99_SLICE_X96Y99_BQ;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_C3 = CLBLM_L_X64Y106_SLICE_X96Y106_BO5;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_C5 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_C1 = 1'b1;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_C4 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_C6 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_C2 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_C3 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_C4 = 1'b1;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_C5 = CLBLM_L_X64Y105_SLICE_X96Y105_BO5;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_C5 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_C6 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_D1 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_D2 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_D3 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_D4 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_D5 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_D6 = 1'b1;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X71Y114_SLICE_X106Y114_A1 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X106Y114_A2 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X106Y114_A3 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X106Y114_A4 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X106Y114_A5 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X106Y114_A6 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X106Y114_AX = CLBLL_R_X71Y110_SLICE_X106Y110_A5Q;
  assign CLBLL_R_X71Y114_SLICE_X106Y114_B1 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X106Y114_B2 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X106Y114_B3 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X106Y114_B4 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X106Y114_B5 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X106Y114_B6 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X106Y114_C1 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X106Y114_C2 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X106Y114_C3 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X106Y114_C4 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X106Y114_C5 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X106Y114_C6 = 1'b1;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_D1 = 1'b1;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_D2 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X106Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_D3 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X106Y114_D1 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X106Y114_D2 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X106Y114_D3 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X106Y114_D4 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X106Y114_D5 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X106Y114_D6 = 1'b1;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_D4 = 1'b1;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_D5 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X106Y114_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_D6 = 1'b1;
  assign RIOB33_X105Y71_IOB_X1Y72_O = CLBLM_R_X103Y76_SLICE_X162Y76_AQ;
  assign RIOB33_X105Y71_IOB_X1Y71_O = CLBLM_R_X103Y75_SLICE_X162Y75_BQ;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X71Y114_SLICE_X107Y114_A1 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X107Y114_A2 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X107Y114_A3 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X107Y114_A4 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X107Y114_A5 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X107Y114_A6 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X107Y114_B1 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X107Y114_B2 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X107Y114_B3 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X107Y114_B4 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X107Y114_B5 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X107Y114_B6 = 1'b1;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_A1 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X107Y114_C1 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X107Y114_C2 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X107Y114_C3 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X107Y114_C4 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X107Y114_C5 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X107Y114_C6 = 1'b1;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_A2 = 1'b1;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_A3 = 1'b1;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_A4 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X107Y114_D1 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X107Y114_D2 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X107Y114_D3 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X107Y114_D4 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X107Y114_D5 = 1'b1;
  assign CLBLL_R_X71Y114_SLICE_X107Y114_D6 = 1'b1;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_A5 = 1'b1;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_A6 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X114Y107_A6 = 1'b1;
  assign CLBLM_L_X70Y135_SLICE_X105Y135_A1 = CLBLM_L_X72Y133_SLICE_X109Y133_CO6;
  assign CLBLM_L_X70Y135_SLICE_X105Y135_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y135_SLICE_X105Y135_A3 = CLBLM_L_X70Y135_SLICE_X105Y135_AQ;
  assign CLBLM_L_X70Y135_SLICE_X105Y135_A4 = CLBLL_R_X71Y133_SLICE_X106Y133_AQ;
  assign CLBLM_L_X70Y135_SLICE_X105Y135_A5 = CLBLM_L_X70Y135_SLICE_X105Y135_A5Q;
  assign CLBLM_L_X70Y135_SLICE_X105Y135_A6 = 1'b1;
  assign CLBLM_R_X63Y122_SLICE_X95Y122_B3 = 1'b1;
  assign CLBLM_L_X70Y135_SLICE_X105Y135_B1 = 1'b1;
  assign CLBLM_L_X70Y111_SLICE_X105Y111_B3 = CLBLM_L_X70Y111_SLICE_X105Y111_AQ;
  assign CLBLM_L_X70Y135_SLICE_X105Y135_B2 = 1'b1;
  assign CLBLM_L_X70Y135_SLICE_X105Y135_B3 = 1'b1;
  assign CLBLM_L_X70Y135_SLICE_X105Y135_B4 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X114Y107_AX = CLBLM_L_X62Y107_SLICE_X93Y107_BQ;
  assign CLBLM_L_X70Y111_SLICE_X105Y111_B4 = CLBLM_L_X70Y111_SLICE_X104Y111_BO5;
  assign CLBLM_L_X70Y135_SLICE_X105Y135_B5 = 1'b1;
  assign CLBLM_L_X70Y135_SLICE_X105Y135_B6 = 1'b1;
  assign CLBLM_L_X70Y135_SLICE_X105Y135_C1 = 1'b1;
  assign CLBLM_L_X70Y111_SLICE_X105Y111_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y135_SLICE_X105Y135_C2 = 1'b1;
  assign CLBLM_L_X70Y135_SLICE_X105Y135_C3 = 1'b1;
  assign CLBLM_L_X70Y135_SLICE_X105Y135_C4 = 1'b1;
  assign CLBLM_L_X70Y135_SLICE_X105Y135_C5 = 1'b1;
  assign CLBLM_L_X70Y111_SLICE_X105Y111_B6 = CLBLM_L_X70Y111_SLICE_X105Y111_CO6;
  assign CLBLM_L_X70Y135_SLICE_X105Y135_C6 = 1'b1;
  assign CLBLM_L_X70Y135_SLICE_X105Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_B1 = 1'b1;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_B2 = 1'b1;
  assign CLBLM_L_X70Y135_SLICE_X105Y135_D1 = 1'b1;
  assign CLBLM_L_X70Y135_SLICE_X105Y135_D2 = 1'b1;
  assign CLBLM_L_X70Y135_SLICE_X105Y135_D3 = 1'b1;
  assign CLBLM_L_X70Y135_SLICE_X105Y135_D4 = 1'b1;
  assign CLBLM_L_X70Y135_SLICE_X105Y135_D5 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X114Y107_B4 = 1'b1;
  assign CLBLM_L_X70Y135_SLICE_X105Y135_D6 = 1'b1;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_B3 = 1'b1;
  assign CLBLM_L_X70Y135_SLICE_X105Y135_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X75Y107_SLICE_X114Y107_B5 = 1'b1;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_B4 = 1'b1;
  assign CLBLM_L_X70Y135_SLICE_X104Y135_A1 = CLBLM_L_X70Y134_SLICE_X105Y134_AQ;
  assign CLBLM_L_X70Y135_SLICE_X104Y135_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y107_SLICE_X114Y107_B6 = 1'b1;
  assign CLBLM_L_X70Y111_SLICE_X105Y111_C1 = CLBLM_L_X70Y111_SLICE_X104Y111_AQ;
  assign CLBLM_L_X70Y135_SLICE_X104Y135_A3 = CLBLM_L_X70Y135_SLICE_X104Y135_AQ;
  assign CLBLM_L_X70Y135_SLICE_X104Y135_A4 = CLBLL_R_X71Y133_SLICE_X106Y133_AQ;
  assign CLBLM_L_X70Y135_SLICE_X104Y135_A5 = CLBLM_L_X70Y135_SLICE_X104Y135_CO5;
  assign CLBLM_L_X70Y135_SLICE_X104Y135_A6 = CLBLM_L_X72Y134_SLICE_X109Y134_AO6;
  assign CLBLM_L_X70Y111_SLICE_X105Y111_C2 = CLBLM_L_X70Y111_SLICE_X104Y111_CO6;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_B5 = 1'b1;
  assign CLBLM_L_X70Y135_SLICE_X104Y135_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y135_SLICE_X104Y135_B2 = CLBLM_L_X70Y135_SLICE_X104Y135_BQ;
  assign CLBLM_L_X70Y111_SLICE_X105Y111_C3 = CLBLM_L_X70Y110_SLICE_X104Y110_BQ;
  assign CLBLM_L_X70Y135_SLICE_X104Y135_B3 = CLBLM_L_X70Y135_SLICE_X104Y135_AQ;
  assign CLBLM_L_X70Y135_SLICE_X104Y135_B4 = CLBLM_L_X72Y134_SLICE_X109Y134_AO6;
  assign CLBLM_L_X70Y135_SLICE_X104Y135_B6 = CLBLM_L_X70Y135_SLICE_X104Y135_CO6;
  assign CLBLM_L_X70Y135_SLICE_X104Y135_B5 = CLBLM_L_X72Y133_SLICE_X109Y133_CO6;
  assign CLBLM_L_X70Y111_SLICE_X105Y111_C4 = CLBLL_R_X71Y111_SLICE_X106Y111_BQ;
  assign CLBLM_L_X70Y135_SLICE_X104Y135_C1 = CLBLL_R_X71Y133_SLICE_X106Y133_AQ;
  assign CLBLM_L_X70Y111_SLICE_X105Y111_C5 = CLBLM_L_X70Y110_SLICE_X104Y110_B5Q;
  assign CLBLM_L_X70Y135_SLICE_X104Y135_C2 = CLBLM_L_X70Y135_SLICE_X105Y135_A5Q;
  assign CLBLM_L_X70Y135_SLICE_X104Y135_C3 = CLBLM_L_X72Y133_SLICE_X109Y133_CO6;
  assign CLBLM_L_X70Y135_SLICE_X104Y135_C4 = 1'b1;
  assign CLBLM_L_X70Y135_SLICE_X104Y135_C5 = 1'b1;
  assign CLBLM_L_X70Y111_SLICE_X105Y111_C6 = CLBLL_R_X71Y111_SLICE_X106Y111_CQ;
  assign CLBLM_L_X70Y135_SLICE_X104Y135_C6 = 1'b1;
  assign CLBLM_L_X70Y135_SLICE_X104Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X67Y97_SLICE_X100Y97_B3 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_D1 = CLBLM_L_X70Y135_SLICE_X104Y135_CO6;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_C1 = 1'b1;
  assign CLBLM_L_X70Y135_SLICE_X104Y135_D1 = 1'b1;
  assign CLBLM_L_X70Y135_SLICE_X104Y135_D2 = 1'b1;
  assign CLBLM_L_X70Y135_SLICE_X104Y135_D3 = 1'b1;
  assign CLBLM_L_X70Y135_SLICE_X104Y135_D4 = 1'b1;
  assign CLBLM_L_X70Y135_SLICE_X104Y135_D5 = 1'b1;
  assign CLBLM_L_X70Y111_SLICE_X105Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X70Y135_SLICE_X104Y135_D6 = 1'b1;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_C2 = 1'b1;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_C3 = 1'b1;
  assign CLBLM_L_X70Y135_SLICE_X104Y135_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_D1 = CLBLL_R_X73Y119_SLICE_X110Y119_BQ;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_C4 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_D1 = CLBLM_R_X63Y105_SLICE_X95Y105_A5Q;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_A1 = CLBLM_R_X65Y100_SLICE_X99Y100_CQ;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_A2 = CLBLM_R_X63Y99_SLICE_X95Y99_AO5;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_C5 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_A3 = CLBLM_R_X65Y101_SLICE_X99Y101_AQ;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_A5 = CLBLM_R_X65Y100_SLICE_X99Y100_A5Q;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_A6 = 1'b1;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_C6 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_T1 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_B1 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_B2 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_B3 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_B4 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_B5 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_B6 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_D1 = CLBLM_L_X72Y119_SLICE_X109Y119_BQ;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_C1 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_C2 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_C3 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_C4 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_C5 = 1'b1;
  assign CLBLM_L_X70Y111_SLICE_X105Y111_D1 = CLBLM_L_X70Y112_SLICE_X105Y112_AQ;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_C6 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_T1 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X70Y111_SLICE_X105Y111_D2 = CLBLM_L_X70Y110_SLICE_X104Y110_B5Q;
  assign CLBLM_L_X70Y111_SLICE_X105Y111_D3 = CLBLL_R_X71Y112_SLICE_X106Y112_AQ;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_D1 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_D2 = 1'b1;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_A6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_D3 = 1'b1;
  assign CLBLM_L_X70Y111_SLICE_X105Y111_D4 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_D4 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_D5 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_D6 = 1'b1;
  assign CLBLM_L_X70Y111_SLICE_X105Y111_D5 = CLBLM_L_X70Y110_SLICE_X104Y110_AQ;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_A1 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_A2 = 1'b1;
  assign CLBLM_L_X70Y111_SLICE_X105Y111_D6 = CLBLM_L_X70Y110_SLICE_X104Y110_BQ;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_A3 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_A4 = 1'b1;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_AX = CLBLM_L_X76Y128_SLICE_X117Y128_CO5;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_A5 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_A6 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_B1 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_B2 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_B3 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_B4 = 1'b1;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_D1 = 1'b1;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_B1 = CLBLM_L_X76Y128_SLICE_X117Y128_B5Q;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_B5 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_B6 = 1'b1;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_D2 = 1'b1;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_B2 = CLBLM_L_X76Y128_SLICE_X117Y128_BQ;
  assign CLBLM_L_X70Y111_SLICE_X105Y111_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_C1 = 1'b1;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_D3 = 1'b1;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_C2 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_C3 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_C4 = 1'b1;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_D4 = 1'b1;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_B4 = CLBLL_R_X77Y128_SLICE_X118Y128_CO6;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_C5 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_C6 = 1'b1;
  assign CLBLM_L_X74Y107_SLICE_X113Y107_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_D5 = 1'b1;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_B5 = CLBLL_R_X77Y128_SLICE_X118Y128_AQ;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_D1 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_D2 = 1'b1;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_D6 = 1'b1;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_B6 = 1'b1;
  assign CLBLM_L_X70Y111_SLICE_X104Y111_A1 = CLBLM_L_X72Y111_SLICE_X109Y111_A5Q;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_D3 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_D4 = 1'b1;
  assign CLBLM_L_X76Y122_SLICE_X116Y122_A4 = CLBLL_R_X75Y123_SLICE_X114Y123_AO6;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_D5 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_T1 = 1'b1;
  assign CLBLM_L_X70Y111_SLICE_X104Y111_A3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y111_SLICE_X104Y111_A4 = CLBLM_L_X72Y111_SLICE_X109Y111_CQ;
  assign CLBLM_L_X72Y108_SLICE_X108Y108_D4 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X70Y111_SLICE_X104Y111_A5 = CLBLM_L_X70Y111_SLICE_X104Y111_BQ;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_C1 = CLBLL_R_X77Y126_SLICE_X118Y126_AQ;
  assign CLBLM_L_X70Y111_SLICE_X104Y111_A6 = 1'b1;
  assign CLBLM_L_X76Y122_SLICE_X116Y122_A5 = CLBLM_L_X76Y122_SLICE_X116Y122_A5Q;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_C2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_C3 = CLBLM_L_X76Y128_SLICE_X116Y128_AQ;
  assign RIOB33_X105Y73_IOB_X1Y74_O = CLBLM_R_X103Y75_SLICE_X162Y75_AQ;
  assign RIOB33_X105Y73_IOB_X1Y73_O = CLBLM_R_X103Y75_SLICE_X163Y75_AQ;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_C4 = CLBLM_L_X76Y128_SLICE_X117Y128_A5Q;
  assign CLBLM_L_X72Y108_SLICE_X108Y108_D5 = CLBLM_L_X72Y108_SLICE_X109Y108_DQ;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_C5 = CLBLL_R_X77Y126_SLICE_X118Y126_BQ;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_C6 = 1'b1;
  assign CLBLM_L_X76Y122_SLICE_X116Y122_A6 = 1'b1;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X72Y108_SLICE_X108Y108_D6 = 1'b1;
  assign CLBLM_L_X70Y111_SLICE_X104Y111_B4 = CLBLM_L_X70Y110_SLICE_X104Y110_B5Q;
  assign CLBLM_L_X70Y111_SLICE_X104Y111_B5 = CLBLM_L_X70Y111_SLICE_X104Y111_CO6;
  assign CLBLM_L_X70Y111_SLICE_X104Y111_B6 = 1'b1;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_D1 = 1'b1;
  assign CLBLM_L_X70Y111_SLICE_X104Y111_BX = CLBLM_L_X70Y111_SLICE_X104Y111_AO5;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_D2 = 1'b1;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_D3 = 1'b1;
  assign CLBLM_R_X67Y97_SLICE_X100Y97_C1 = 1'b1;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_D4 = 1'b1;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_D5 = 1'b1;
  assign CLBLM_L_X70Y136_SLICE_X105Y136_A1 = CLBLM_L_X76Y125_SLICE_X116Y125_AQ;
  assign CLBLM_L_X70Y136_SLICE_X105Y136_A2 = CLBLL_R_X73Y133_SLICE_X111Y133_A5Q;
  assign CLBLM_L_X70Y136_SLICE_X105Y136_A3 = CLBLM_L_X70Y136_SLICE_X105Y136_AQ;
  assign CLBLM_L_X70Y136_SLICE_X105Y136_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y136_SLICE_X105Y136_A5 = CLBLM_L_X70Y136_SLICE_X104Y136_AQ;
  assign CLBLM_L_X70Y136_SLICE_X105Y136_A6 = 1'b1;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_D6 = 1'b1;
  assign CLBLM_L_X70Y111_SLICE_X104Y111_C5 = CLBLM_L_X72Y111_SLICE_X109Y111_AQ;
  assign CLBLM_L_X70Y136_SLICE_X105Y136_B1 = CLBLM_L_X70Y136_SLICE_X105Y136_AQ;
  assign CLBLM_L_X70Y136_SLICE_X105Y136_B2 = CLBLM_L_X70Y136_SLICE_X105Y136_BQ;
  assign CLBLM_L_X70Y136_SLICE_X105Y136_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y111_SLICE_X104Y111_C6 = CLBLM_L_X70Y112_SLICE_X104Y112_AQ;
  assign CLBLM_L_X70Y136_SLICE_X105Y136_B4 = CLBLL_R_X73Y133_SLICE_X111Y133_A5Q;
  assign CLBLM_L_X70Y136_SLICE_X105Y136_B5 = CLBLM_L_X70Y136_SLICE_X104Y136_AQ;
  assign CLBLM_L_X70Y136_SLICE_X105Y136_B6 = 1'b1;
  assign CLBLM_R_X67Y97_SLICE_X100Y97_C2 = 1'b1;
  assign CLBLM_L_X70Y136_SLICE_X105Y136_C1 = CLBLM_L_X70Y136_SLICE_X104Y136_AQ;
  assign CLBLM_L_X70Y136_SLICE_X105Y136_C2 = CLBLL_R_X75Y133_SLICE_X115Y133_BQ;
  assign CLBLM_L_X70Y136_SLICE_X105Y136_C3 = CLBLM_L_X70Y136_SLICE_X105Y136_BQ;
  assign CLBLM_L_X70Y136_SLICE_X105Y136_C4 = CLBLM_L_X70Y136_SLICE_X105Y136_AQ;
  assign CLBLM_L_X70Y136_SLICE_X105Y136_C5 = 1'b1;
  assign CLBLM_L_X70Y136_SLICE_X105Y136_C6 = CLBLM_L_X70Y136_SLICE_X104Y136_BQ;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X70Y136_SLICE_X105Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X70Y111_SLICE_X104Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X70Y136_SLICE_X105Y136_D1 = 1'b1;
  assign CLBLM_L_X70Y136_SLICE_X105Y136_D2 = 1'b1;
  assign CLBLM_L_X70Y136_SLICE_X105Y136_D3 = 1'b1;
  assign CLBLM_L_X70Y136_SLICE_X105Y136_D4 = 1'b1;
  assign CLBLM_L_X70Y136_SLICE_X105Y136_D5 = 1'b1;
  assign CLBLM_L_X70Y136_SLICE_X105Y136_D6 = 1'b1;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_A1 = CLBLM_L_X76Y128_SLICE_X117Y128_A5Q;
  assign CLBLM_L_X70Y136_SLICE_X105Y136_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_A2 = CLBLM_L_X76Y128_SLICE_X116Y128_BQ;
  assign CLBLM_L_X70Y136_SLICE_X104Y136_A1 = CLBLM_L_X70Y136_SLICE_X105Y136_BQ;
  assign CLBLM_L_X70Y136_SLICE_X104Y136_A2 = CLBLM_L_X70Y136_SLICE_X104Y136_BQ;
  assign CLBLM_L_X70Y136_SLICE_X104Y136_A3 = CLBLM_L_X70Y136_SLICE_X104Y136_AQ;
  assign CLBLM_L_X70Y136_SLICE_X104Y136_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y136_SLICE_X104Y136_A5 = CLBLM_L_X70Y136_SLICE_X105Y136_AQ;
  assign CLBLM_L_X70Y136_SLICE_X104Y136_A6 = CLBLL_R_X73Y133_SLICE_X111Y133_A5Q;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_A3 = CLBLM_L_X76Y128_SLICE_X116Y128_AQ;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_A4 = CLBLL_R_X77Y126_SLICE_X118Y126_AQ;
  assign CLBLM_L_X70Y136_SLICE_X104Y136_B1 = CLBLM_L_X70Y136_SLICE_X105Y136_BQ;
  assign CLBLM_L_X70Y136_SLICE_X104Y136_B2 = CLBLM_L_X70Y136_SLICE_X104Y136_BQ;
  assign CLBLM_L_X70Y136_SLICE_X104Y136_B3 = CLBLM_L_X70Y136_SLICE_X104Y136_AQ;
  assign CLBLM_L_X70Y136_SLICE_X104Y136_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y136_SLICE_X104Y136_B5 = CLBLM_L_X70Y136_SLICE_X105Y136_AQ;
  assign CLBLM_L_X70Y136_SLICE_X104Y136_B6 = CLBLL_R_X73Y133_SLICE_X111Y133_A5Q;
  assign CLBLM_L_X72Y106_SLICE_X109Y106_A1 = CLBLL_R_X73Y108_SLICE_X110Y108_A5Q;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_A5 = CLBLL_R_X77Y126_SLICE_X118Y126_BQ;
  assign CLBLM_L_X72Y106_SLICE_X109Y106_A2 = CLBLL_R_X71Y107_SLICE_X106Y107_C5Q;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_A6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y136_SLICE_X104Y136_C1 = 1'b1;
  assign CLBLM_L_X70Y136_SLICE_X104Y136_C2 = 1'b1;
  assign CLBLM_L_X70Y136_SLICE_X104Y136_C3 = 1'b1;
  assign CLBLM_L_X70Y136_SLICE_X104Y136_C4 = 1'b1;
  assign CLBLM_L_X70Y136_SLICE_X104Y136_C5 = 1'b1;
  assign CLBLM_L_X70Y136_SLICE_X104Y136_C6 = 1'b1;
  assign CLBLM_L_X72Y106_SLICE_X109Y106_A3 = CLBLM_L_X62Y90_SLICE_X92Y90_AQ;
  assign CLBLM_L_X72Y106_SLICE_X109Y106_A4 = CLBLL_R_X71Y107_SLICE_X106Y107_CQ;
  assign CLBLM_L_X70Y136_SLICE_X104Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X72Y106_SLICE_X109Y106_A5 = CLBLM_L_X72Y106_SLICE_X108Y106_AQ;
  assign CLBLM_L_X70Y111_SLICE_X104Y111_D4 = CLBLM_L_X72Y111_SLICE_X108Y111_BQ;
  assign CLBLM_L_X70Y136_SLICE_X104Y136_D1 = 1'b1;
  assign CLBLM_L_X70Y136_SLICE_X104Y136_D2 = 1'b1;
  assign CLBLM_L_X70Y111_SLICE_X104Y111_D5 = CLBLM_L_X70Y110_SLICE_X104Y110_AQ;
  assign CLBLM_L_X70Y136_SLICE_X104Y136_D3 = 1'b1;
  assign CLBLM_L_X70Y136_SLICE_X104Y136_D4 = 1'b1;
  assign CLBLM_L_X70Y136_SLICE_X104Y136_D5 = 1'b1;
  assign CLBLM_L_X70Y136_SLICE_X104Y136_D6 = 1'b1;
  assign CLBLM_L_X72Y106_SLICE_X109Y106_A6 = CLBLM_L_X74Y107_SLICE_X112Y107_DQ;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_AX = CLBLM_L_X76Y128_SLICE_X116Y128_CQ;
  assign CLBLM_L_X70Y136_SLICE_X104Y136_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_B1 = CLBLM_L_X76Y128_SLICE_X117Y128_A5Q;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_B2 = CLBLL_R_X77Y126_SLICE_X118Y126_AQ;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_A1 = CLBLM_L_X70Y101_SLICE_X104Y101_DO6;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_A2 = CLBLM_R_X65Y103_SLICE_X99Y103_DO6;
  assign CLBLM_L_X74Y103_SLICE_X113Y103_B2 = CLBLM_L_X74Y103_SLICE_X113Y103_BQ;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_B3 = CLBLM_L_X76Y128_SLICE_X116Y128_AQ;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_A3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_A4 = CLBLM_R_X65Y104_SLICE_X98Y104_C5Q;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_A5 = CLBLM_R_X65Y104_SLICE_X99Y104_DO6;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_A6 = CLBLM_R_X65Y104_SLICE_X98Y104_CQ;
  assign CLBLM_L_X72Y106_SLICE_X109Y106_B1 = CLBLL_R_X71Y107_SLICE_X106Y107_C5Q;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_B1 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_B2 = 1'b1;
  assign CLBLM_L_X72Y106_SLICE_X109Y106_B2 = CLBLL_R_X73Y107_SLICE_X110Y107_BQ;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_B5 = CLBLL_R_X77Y126_SLICE_X118Y126_BQ;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_B3 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_B4 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_B5 = 1'b1;
  assign CLBLM_L_X72Y106_SLICE_X109Y106_B3 = CLBLM_L_X78Y106_SLICE_X120Y106_AQ;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_B6 = CLBLM_L_X76Y128_SLICE_X116Y128_BQ;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_B6 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_C5 = 1'b1;
  assign CLBLM_L_X72Y106_SLICE_X109Y106_B4 = CLBLL_R_X71Y107_SLICE_X106Y107_CQ;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_C6 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_C1 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_C2 = 1'b1;
  assign CLBLM_L_X72Y106_SLICE_X109Y106_B5 = CLBLM_L_X72Y106_SLICE_X108Y106_AQ;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_C3 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_C4 = 1'b1;
  assign CLBLM_L_X76Y122_SLICE_X116Y122_B3 = 1'b1;
  assign CLBLM_L_X72Y106_SLICE_X109Y106_B6 = CLBLL_R_X73Y108_SLICE_X110Y108_A5Q;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_D1 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_D2 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_D3 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_D4 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_D5 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_D6 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_A1 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_A2 = 1'b1;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_C1 = CLBLM_L_X76Y125_SLICE_X116Y125_A5Q;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_A3 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_A4 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_A5 = 1'b1;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_C2 = CLBLM_L_X76Y128_SLICE_X116Y128_AQ;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_A6 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_B1 = 1'b1;
  assign CLBLM_L_X72Y106_SLICE_X109Y106_C1 = CLBLM_L_X72Y106_SLICE_X109Y106_AO6;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_C3 = CLBLM_L_X76Y129_SLICE_X116Y129_B5Q;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_B2 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_B3 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_B4 = 1'b1;
  assign CLBLM_L_X72Y106_SLICE_X109Y106_C2 = CLBLM_L_X72Y106_SLICE_X108Y106_A5Q;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_C4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_B5 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_B6 = 1'b1;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_C5 = CLBLM_L_X76Y130_SLICE_X116Y130_DQ;
  assign CLBLM_L_X72Y106_SLICE_X109Y106_C3 = CLBLM_L_X72Y107_SLICE_X109Y107_BO5;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_C1 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_C2 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_C3 = 1'b1;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_C6 = 1'b1;
  assign CLBLM_L_X72Y106_SLICE_X109Y106_C4 = CLBLM_L_X72Y107_SLICE_X109Y107_CO6;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_C4 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_C5 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_C6 = 1'b1;
  assign CLBLM_L_X72Y106_SLICE_X109Y106_C5 = CLBLM_L_X74Y107_SLICE_X112Y107_BQ;
  assign CLBLM_L_X72Y106_SLICE_X109Y106_C6 = CLBLM_L_X72Y106_SLICE_X109Y106_BO6;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_D1 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_D2 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_D3 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_D4 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_D5 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_D6 = 1'b1;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOB33_X105Y75_IOB_X1Y75_O = CLBLM_R_X103Y75_SLICE_X162Y75_CQ;
  assign RIOB33_X105Y75_IOB_X1Y76_O = CLBLM_R_X103Y75_SLICE_X163Y75_BQ;
  assign CLBLM_L_X76Y122_SLICE_X116Y122_B6 = CLBLL_R_X75Y123_SLICE_X114Y123_AO6;
  assign CLBLM_L_X80Y132_SLICE_X124Y132_AX = CLBLL_R_X77Y128_SLICE_X119Y128_BQ;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_D1 = CLBLL_R_X77Y128_SLICE_X118Y128_AQ;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_D2 = CLBLL_R_X77Y126_SLICE_X118Y126_BQ;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_D3 = CLBLM_L_X76Y128_SLICE_X116Y128_AQ;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_D4 = CLBLM_L_X76Y128_SLICE_X116Y128_BQ;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_D5 = CLBLM_L_X76Y128_SLICE_X117Y128_A5Q;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_D6 = 1'b1;
  assign CLBLM_L_X72Y106_SLICE_X109Y106_D6 = 1'b1;
  assign CLBLM_L_X82Y130_SLICE_X128Y130_D4 = 1'b1;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_T1 = 1'b1;
  assign CLBLM_R_X103Y75_SLICE_X162Y75_B5 = 1'b1;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_D1 = 1'b0;
  assign CLBLM_L_X82Y130_SLICE_X128Y130_D5 = 1'b1;
  assign RIOI3_X105Y55_ILOGIC_X1Y56_D = RIOB33_X105Y55_IOB_X1Y56_I;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_A2 = CLBLM_R_X65Y104_SLICE_X99Y104_DO6;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_A3 = CLBLM_R_X65Y103_SLICE_X99Y103_AQ;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_A4 = CLBLM_R_X65Y104_SLICE_X98Y104_C5Q;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_A5 = CLBLM_R_X65Y102_SLICE_X99Y102_AQ;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_A6 = CLBLM_R_X65Y104_SLICE_X98Y104_CQ;
  assign RIOI3_X105Y55_ILOGIC_X1Y55_D = RIOB33_X105Y55_IOB_X1Y55_I;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_B1 = CLBLM_R_X65Y104_SLICE_X98Y104_B5Q;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_B2 = CLBLM_R_X65Y104_SLICE_X98Y104_BQ;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_B3 = CLBLM_R_X65Y103_SLICE_X98Y103_A5Q;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_B4 = CLBLM_R_X65Y103_SLICE_X98Y103_BQ;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_B5 = CLBLM_R_X65Y103_SLICE_X99Y103_BQ;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_B6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X103Y75_SLICE_X162Y75_B6 = 1'b1;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_C1 = CLBLM_R_X65Y103_SLICE_X99Y103_BQ;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_C2 = CLBLM_R_X65Y104_SLICE_X99Y104_AQ;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_C3 = CLBLM_R_X65Y104_SLICE_X99Y104_A5Q;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_C4 = CLBLM_R_X65Y104_SLICE_X98Y104_B5Q;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_C5 = CLBLM_R_X65Y104_SLICE_X98Y104_BQ;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_C6 = CLBLM_R_X65Y103_SLICE_X98Y103_BQ;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_D1 = 1'b1;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_D2 = CLBLM_R_X65Y104_SLICE_X98Y104_CQ;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_D3 = CLBLM_R_X65Y105_SLICE_X98Y105_B5Q;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_D4 = CLBLM_R_X65Y103_SLICE_X99Y103_CO6;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_D5 = CLBLM_R_X65Y103_SLICE_X99Y103_AQ;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_D6 = CLBLM_R_X65Y104_SLICE_X98Y104_C5Q;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_A1 = CLBLM_R_X65Y104_SLICE_X98Y104_B5Q;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_A2 = CLBLM_R_X65Y103_SLICE_X98Y103_BQ;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_A3 = CLBLM_R_X65Y103_SLICE_X98Y103_AQ;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_A4 = CLBLM_R_X65Y104_SLICE_X98Y104_BQ;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_A6 = CLBLM_R_X65Y103_SLICE_X98Y103_A5Q;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_AX = CLBLM_R_X65Y104_SLICE_X99Y104_B5Q;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_B1 = CLBLM_R_X65Y104_SLICE_X98Y104_B5Q;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_B2 = CLBLM_R_X65Y103_SLICE_X98Y103_BQ;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_B3 = CLBLM_R_X65Y103_SLICE_X98Y103_AQ;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_B4 = CLBLM_R_X65Y104_SLICE_X98Y104_BQ;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_B6 = CLBLM_R_X65Y103_SLICE_X98Y103_A5Q;
  assign RIOB33_X105Y77_IOB_X1Y77_O = CLBLM_R_X103Y76_SLICE_X163Y76_AQ;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_C1 = CLBLM_R_X65Y103_SLICE_X99Y103_AQ;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_C2 = CLBLM_R_X65Y104_SLICE_X98Y104_CQ;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_C3 = CLBLM_L_X64Y103_SLICE_X97Y103_BQ;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_C4 = CLBLM_L_X64Y103_SLICE_X97Y103_AQ;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_C5 = CLBLM_R_X65Y104_SLICE_X98Y104_C5Q;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_C6 = CLBLM_L_X64Y105_SLICE_X97Y105_AQ;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_A1 = CLBLL_R_X71Y109_SLICE_X106Y109_B5Q;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_A3 = CLBLL_R_X71Y117_SLICE_X106Y117_AQ;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_A4 = CLBLM_L_X72Y123_SLICE_X108Y123_A5Q;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_A5 = CLBLM_L_X68Y107_SLICE_X103Y107_AO6;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_A6 = 1'b1;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_D1 = CLBLM_L_X64Y100_SLICE_X97Y100_AQ;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_D2 = CLBLM_R_X65Y104_SLICE_X99Y104_B5Q;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_D3 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_B2 = CLBLL_R_X71Y117_SLICE_X106Y117_BQ;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_B3 = CLBLL_R_X71Y117_SLICE_X106Y117_AQ;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_B4 = CLBLM_R_X67Y111_SLICE_X100Y111_A5Q;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_B5 = CLBLM_L_X68Y105_SLICE_X102Y105_DO6;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_B6 = 1'b1;
  assign CLBLM_L_X82Y130_SLICE_X128Y130_D6 = 1'b1;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_C1 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_C2 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_C3 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_C4 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_C5 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_C6 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_D1 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_T1 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_D1 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_D2 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_D3 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_D4 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_D5 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_D6 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_T1 = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_D1 = CLBLM_L_X72Y119_SLICE_X108Y119_CQ;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_T1 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_A1 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_A2 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_A3 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_A4 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_A5 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_A6 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_B1 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_B2 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_B3 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_B4 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_B5 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_B6 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_C1 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_C2 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_C3 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_C4 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_C5 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_C6 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_D1 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_D2 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_D3 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_D4 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_D5 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_D6 = 1'b1;
  assign LIOB33_X0Y95_IOB_X0Y96_O = CLBLM_R_X63Y97_SLICE_X95Y97_AQ;
  assign LIOB33_X0Y95_IOB_X0Y95_O = CLBLM_L_X70Y101_SLICE_X104Y101_AQ;
  assign LIOB33_SING_X0Y50_IOB_X0Y50_O = CLBLM_L_X60Y97_SLICE_X90Y97_DQ;
  assign CLBLM_L_X68Y96_SLICE_X102Y96_D4 = CLBLM_L_X68Y99_SLICE_X102Y99_BO6;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_A1 = CLBLM_R_X65Y104_SLICE_X99Y104_AQ;
  assign CLBLM_L_X68Y96_SLICE_X102Y96_D5 = CLBLM_L_X62Y95_SLICE_X92Y95_BQ;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_A2 = CLBLM_R_X65Y103_SLICE_X99Y103_BQ;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_A3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_A4 = CLBLM_R_X65Y104_SLICE_X98Y104_AO5;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_A5 = CLBLM_R_X65Y104_SLICE_X99Y104_A5Q;
  assign CLBLM_L_X68Y96_SLICE_X102Y96_D6 = CLBLM_L_X68Y96_SLICE_X102Y96_BO6;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_A6 = 1'b1;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_B1 = 1'b1;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_B2 = CLBLM_R_X65Y104_SLICE_X99Y104_BQ;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_B3 = CLBLM_R_X65Y105_SLICE_X99Y105_C5Q;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_B4 = CLBLM_L_X64Y104_SLICE_X97Y104_AQ;
  assign CLBLM_L_X78Y106_SLICE_X121Y106_B1 = 1'b1;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_B6 = CLBLM_R_X63Y103_SLICE_X95Y103_BO5;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_BX = CLBLM_R_X65Y105_SLICE_X98Y105_B5Q;
  assign CLBLM_L_X78Y106_SLICE_X121Y106_B2 = 1'b1;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_C1 = CLBLM_R_X65Y104_SLICE_X99Y104_A5Q;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_C2 = CLBLM_R_X65Y104_SLICE_X98Y104_C5Q;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_C3 = CLBLM_R_X65Y103_SLICE_X98Y103_CO6;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_C4 = CLBLM_R_X65Y104_SLICE_X98Y104_CQ;
  assign CLBLM_L_X78Y106_SLICE_X121Y106_B3 = 1'b1;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_C5 = CLBLM_R_X65Y104_SLICE_X99Y104_AQ;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_C6 = CLBLM_R_X65Y103_SLICE_X99Y103_BQ;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X78Y106_SLICE_X121Y106_B4 = 1'b1;
  assign RIOI3_X105Y59_ILOGIC_X1Y60_D = RIOB33_X105Y59_IOB_X1Y60_I;
  assign RIOI3_X105Y59_ILOGIC_X1Y59_D = RIOB33_X105Y59_IOB_X1Y59_I;
  assign RIOB33_X105Y79_IOB_X1Y79_O = CLBLL_R_X83Y94_SLICE_X130Y94_A5Q;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_D1 = 1'b1;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_D2 = 1'b1;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_D3 = 1'b1;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_D4 = CLBLM_R_X65Y104_SLICE_X99Y104_A5Q;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_D5 = CLBLM_R_X65Y104_SLICE_X99Y104_AQ;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_D6 = CLBLM_R_X65Y103_SLICE_X99Y103_BQ;
  assign RIOB33_X105Y79_IOB_X1Y80_O = 1'b0;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_A1 = CLBLM_R_X65Y104_SLICE_X98Y104_B5Q;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_A2 = CLBLM_R_X65Y104_SLICE_X98Y104_BQ;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_A3 = CLBLM_R_X65Y103_SLICE_X98Y103_A5Q;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_A4 = CLBLM_R_X65Y103_SLICE_X99Y103_BQ;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_A5 = CLBLM_R_X65Y103_SLICE_X98Y103_BQ;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_A6 = 1'b1;
  assign LIOB33_X0Y143_IOB_X0Y143_O = 1'b1;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_B1 = CLBLM_R_X65Y104_SLICE_X98Y104_B5Q;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_B2 = CLBLM_R_X65Y104_SLICE_X98Y104_BQ;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_B3 = CLBLM_R_X65Y103_SLICE_X98Y103_A5Q;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_B4 = 1'b1;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_B6 = 1'b1;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_C2 = CLBLM_R_X65Y104_SLICE_X98Y104_CQ;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_C3 = CLBLM_R_X65Y104_SLICE_X99Y104_AQ;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_C4 = CLBLM_R_X65Y104_SLICE_X98Y104_C5Q;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_C5 = CLBLM_R_X65Y104_SLICE_X98Y104_DO6;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_C6 = 1'b1;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_D1 = CLBLM_R_X65Y103_SLICE_X98Y103_BQ;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_D2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_D3 = CLBLM_R_X65Y104_SLICE_X98Y104_BQ;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_D4 = CLBLM_R_X65Y103_SLICE_X98Y103_A5Q;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_D5 = CLBLM_R_X65Y104_SLICE_X98Y104_B5Q;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_D6 = CLBLM_R_X65Y103_SLICE_X99Y103_BQ;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_A4 = CLBLM_L_X72Y128_SLICE_X108Y128_A5Q;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_A5 = CLBLM_L_X72Y128_SLICE_X108Y128_AQ;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_A6 = CLBLM_L_X72Y127_SLICE_X108Y127_A5Q;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_T1 = 1'b1;
  assign LIOB33_SING_X0Y99_IOB_X0Y99_O = RIOB33_X105Y61_IOB_X1Y62_I;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_B3 = CLBLM_L_X72Y126_SLICE_X108Y126_CO6;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_B4 = CLBLM_L_X72Y127_SLICE_X109Y127_BQ;
  assign LIOB33_X0Y181_IOB_X0Y182_O = CLBLM_L_X70Y126_SLICE_X104Y126_DO6;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_B5 = CLBLM_L_X72Y127_SLICE_X108Y127_A5Q;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_B6 = 1'b1;
  assign RIOB33_X105Y173_IOB_X1Y174_O = CLBLM_L_X70Y111_SLICE_X105Y111_DO6;
  assign LIOB33_X0Y181_IOB_X0Y181_O = CLBLM_L_X64Y106_SLICE_X97Y106_AO6;
  assign CLBLM_L_X78Y106_SLICE_X120Y106_A3 = 1'b1;
  assign CLBLM_L_X78Y106_SLICE_X120Y106_A4 = 1'b1;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_A4 = 1'b1;
  assign CLBLM_L_X78Y106_SLICE_X120Y106_A5 = 1'b1;
  assign CLBLM_L_X78Y106_SLICE_X120Y106_A6 = 1'b1;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X78Y106_SLICE_X120Y106_AX = CLBLM_L_X72Y106_SLICE_X108Y106_AQ;
  assign CLBLM_L_X78Y106_SLICE_X120Y106_B1 = 1'b1;
  assign CLBLM_L_X78Y106_SLICE_X120Y106_B2 = 1'b1;
  assign CLBLM_L_X78Y106_SLICE_X120Y106_B3 = 1'b1;
  assign CLBLM_L_X78Y106_SLICE_X120Y106_B4 = 1'b1;
  assign LIOB33_SING_X0Y100_IOB_X0Y100_O = RIOB33_X105Y57_IOB_X1Y57_I;
  assign CLBLM_L_X78Y106_SLICE_X120Y106_B5 = 1'b1;
  assign CLBLM_L_X78Y106_SLICE_X120Y106_B6 = 1'b1;
  assign CLBLM_L_X72Y133_SLICE_X108Y133_C5 = CLBLM_L_X72Y132_SLICE_X108Y132_AQ;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_D5 = CLBLM_L_X72Y126_SLICE_X108Y126_CO6;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_D6 = CLBLM_L_X72Y128_SLICE_X108Y128_DQ;
  assign CLBLM_L_X72Y133_SLICE_X108Y133_C6 = CLBLM_L_X72Y133_SLICE_X108Y133_DO6;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_A1 = CLBLM_R_X63Y106_SLICE_X94Y106_AO6;
  assign CLBLM_L_X78Y106_SLICE_X120Y106_C1 = 1'b1;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_A2 = CLBLM_R_X65Y106_SLICE_X99Y106_C5Q;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_A3 = CLBLM_R_X65Y105_SLICE_X99Y105_AQ;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_A5 = CLBLM_R_X65Y105_SLICE_X98Y105_CQ;
  assign CLBLM_L_X78Y106_SLICE_X120Y106_C2 = 1'b1;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_A6 = 1'b1;
  assign RIOB33_X105Y81_IOB_X1Y81_O = CLBLL_R_X71Y110_SLICE_X106Y110_A5Q;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_B1 = CLBLM_R_X65Y100_SLICE_X99Y100_A5Q;
  assign CLBLM_L_X78Y106_SLICE_X120Y106_C3 = 1'b1;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_B2 = CLBLM_R_X65Y100_SLICE_X99Y100_CQ;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_B3 = CLBLM_R_X65Y104_SLICE_X99Y104_BQ;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_B4 = CLBLM_R_X65Y105_SLICE_X99Y105_D5Q;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X78Y106_SLICE_X120Y106_C4 = 1'b1;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_B6 = 1'b1;
  assign LIOB33_X0Y123_IOB_X0Y124_O = CLBLL_L_X34Y123_SLICE_X50Y123_AO6;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_C1 = CLBLM_R_X65Y105_SLICE_X99Y105_C5Q;
  assign CLBLM_L_X78Y106_SLICE_X120Y106_C5 = 1'b1;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_C2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_C3 = CLBLM_R_X65Y105_SLICE_X99Y105_D5Q;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_C4 = CLBLM_L_X72Y118_SLICE_X108Y118_CQ;
  assign CLBLM_L_X74Y122_SLICE_X113Y122_B5 = 1'b1;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_B3 = CLBLM_L_X62Y107_SLICE_X93Y107_A5Q;
  assign CLBLM_L_X78Y106_SLICE_X120Y106_C6 = 1'b1;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_C5 = CLBLM_R_X63Y101_SLICE_X94Y101_BO5;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_C6 = 1'b1;
  assign CLBLM_L_X74Y122_SLICE_X113Y122_B6 = 1'b1;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_B4 = CLBLL_R_X75Y107_SLICE_X114Y107_AQ;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_D1 = CLBLM_L_X64Y105_SLICE_X97Y105_CQ;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_B5 = CLBLM_L_X60Y101_SLICE_X90Y101_BQ;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_D2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_D3 = CLBLM_R_X65Y105_SLICE_X99Y105_DQ;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_D4 = CLBLM_R_X65Y105_SLICE_X99Y105_D5Q;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_D5 = CLBLM_R_X63Y101_SLICE_X94Y101_BO5;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_D6 = 1'b1;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X78Y106_SLICE_X120Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_A1 = CLBLM_R_X65Y105_SLICE_X98Y105_B5Q;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_A2 = CLBLM_R_X65Y104_SLICE_X98Y104_AO6;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_A3 = CLBLM_R_X65Y105_SLICE_X98Y105_AQ;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_A4 = CLBLM_R_X65Y104_SLICE_X99Y104_B5Q;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_A6 = 1'b1;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_B1 = CLBLM_L_X64Y106_SLICE_X97Y106_B5Q;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_B2 = CLBLM_R_X65Y105_SLICE_X98Y105_BQ;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_B4 = CLBLM_L_X64Y106_SLICE_X97Y106_C5Q;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_B5 = CLBLM_R_X65Y105_SLICE_X99Y105_AQ;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_B6 = CLBLM_L_X64Y106_SLICE_X97Y106_AQ;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_BX = CLBLM_R_X65Y105_SLICE_X98Y105_AQ;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_C1 = CLBLM_R_X65Y105_SLICE_X98Y105_BQ;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_C2 = CLBLM_L_X64Y106_SLICE_X97Y106_AO6;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_C3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_C4 = CLBLM_R_X65Y105_SLICE_X99Y105_AQ;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_A2 = CLBLL_R_X71Y124_SLICE_X106Y124_A5Q;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_A3 = CLBLL_R_X71Y125_SLICE_X106Y125_DO6;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_A4 = CLBLL_R_X71Y110_SLICE_X106Y110_A5Q;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_A5 = CLBLL_R_X71Y114_SLICE_X106Y114_AQ;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_A6 = 1'b1;
  assign CLBLM_L_X74Y122_SLICE_X113Y122_C5 = 1'b1;
  assign CLBLM_L_X74Y122_SLICE_X113Y122_C6 = 1'b1;
  assign CLBLM_L_X78Y106_SLICE_X120Y106_D1 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_B1 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_B2 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_B3 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_B4 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_B5 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_B6 = 1'b1;
  assign CLBLM_L_X78Y106_SLICE_X120Y106_D2 = 1'b1;
  assign CLBLM_L_X78Y106_SLICE_X120Y106_D3 = 1'b1;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_D1 = CLBLM_L_X70Y103_SLICE_X104Y103_AQ;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_C1 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_C2 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_C3 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_C4 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_C5 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_C6 = 1'b1;
  assign CLBLM_L_X74Y122_SLICE_X113Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X78Y106_SLICE_X120Y106_D4 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X78Y106_SLICE_X120Y106_D5 = 1'b1;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign LIOB33_SING_X0Y149_IOB_X0Y149_O = CLBLM_R_X67Y105_SLICE_X101Y105_AO6;
  assign CLBLM_L_X78Y106_SLICE_X120Y106_D6 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_D1 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_D2 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_D3 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_D4 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_D5 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_D6 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_T1 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y122_SLICE_X113Y122_D1 = 1'b1;
  assign CLBLM_L_X74Y122_SLICE_X113Y122_D2 = 1'b1;
  assign CLBLM_L_X74Y122_SLICE_X113Y122_D3 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_A1 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_A2 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_A3 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_A4 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_A5 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_A6 = 1'b1;
  assign CLBLM_L_X74Y122_SLICE_X113Y122_D4 = 1'b1;
  assign CLBLM_L_X74Y122_SLICE_X113Y122_D5 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_B1 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_B2 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_B3 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_B4 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_B5 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_B6 = 1'b1;
  assign CLBLM_L_X74Y122_SLICE_X113Y122_D6 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_C1 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_C2 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_C3 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_C4 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_C5 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_C6 = 1'b1;
  assign CLBLM_L_X74Y122_SLICE_X113Y122_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_D1 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_D2 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_D3 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_D4 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_D5 = 1'b1;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_D6 = 1'b1;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y122_SLICE_X112Y122_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y112_SLICE_X105Y112_A6 = 1'b1;
  assign CLBLM_L_X74Y122_SLICE_X112Y122_A2 = CLBLL_R_X75Y128_SLICE_X115Y128_BO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_D1 = 1'b1;
  assign CLBLM_L_X74Y122_SLICE_X112Y122_A3 = CLBLM_L_X74Y122_SLICE_X112Y122_AQ;
  assign CLBLM_L_X74Y122_SLICE_X112Y122_A4 = CLBLL_R_X73Y122_SLICE_X111Y122_AQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_T1 = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_D1 = 1'b0;
  assign CLBLM_L_X74Y122_SLICE_X112Y122_A5 = CLBLM_L_X74Y122_SLICE_X112Y122_A5Q;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_A4 = CLBLM_R_X63Y105_SLICE_X94Y105_CQ;
  assign CLBLM_L_X74Y122_SLICE_X112Y122_A6 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_D1 = 1'b1;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_A5 = CLBLM_R_X63Y105_SLICE_X95Y105_A5Q;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_T1 = 1'b1;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_A6 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_T1 = 1'b1;
  assign CLBLM_L_X70Y112_SLICE_X105Y112_B4 = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_D1 = 1'b0;
  assign LIOB33_SING_X0Y150_IOB_X0Y150_O = CLBLM_L_X74Y129_SLICE_X113Y129_BO6;
  assign CLBLM_L_X70Y112_SLICE_X105Y112_B6 = 1'b1;
  assign CLBLM_L_X74Y122_SLICE_X112Y122_B1 = CLBLM_L_X76Y130_SLICE_X116Y130_DQ;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_T1 = 1'b1;
  assign CLBLM_L_X74Y122_SLICE_X112Y122_B2 = CLBLM_L_X74Y122_SLICE_X112Y122_BQ;
  assign CLBLM_L_X74Y122_SLICE_X112Y122_B3 = CLBLM_L_X76Y125_SLICE_X117Y125_BQ;
  assign CLBLM_L_X74Y122_SLICE_X112Y122_B4 = CLBLM_L_X74Y123_SLICE_X112Y123_BQ;
  assign CLBLM_L_X74Y122_SLICE_X112Y122_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y112_SLICE_X105Y112_C1 = CLBLM_L_X68Y112_SLICE_X103Y112_BQ;
  assign CLBLM_L_X74Y122_SLICE_X112Y122_B6 = CLBLM_L_X72Y122_SLICE_X108Y122_CQ;
  assign CLBLM_L_X70Y112_SLICE_X105Y112_C2 = CLBLL_R_X71Y111_SLICE_X106Y111_A5Q;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_D1 = CLBLL_R_X77Y113_SLICE_X118Y113_AQ;
  assign CLBLM_L_X70Y112_SLICE_X105Y112_C3 = CLBLL_R_X71Y108_SLICE_X107Y108_A5Q;
  assign RIOB33_X105Y83_IOB_X1Y84_O = CLBLM_L_X72Y118_SLICE_X108Y118_D5Q;
  assign RIOB33_X105Y83_IOB_X1Y83_O = CLBLM_R_X63Y105_SLICE_X95Y105_AQ;
  assign CLBLM_L_X70Y112_SLICE_X105Y112_C4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign RIOI3_X105Y105_OLOGIC_X1Y105_D1 = CLBLM_R_X65Y111_SLICE_X98Y111_AQ;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_T1 = 1'b1;
  assign CLBLM_L_X70Y112_SLICE_X105Y112_C5 = CLBLM_L_X70Y112_SLICE_X105Y112_B5Q;
  assign CLBLM_L_X70Y112_SLICE_X105Y112_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_D1 = CLBLM_R_X103Y69_SLICE_X162Y69_AQ;
  assign CLBLM_L_X74Y122_SLICE_X112Y122_C1 = 1'b1;
  assign CLBLM_L_X74Y122_SLICE_X112Y122_C2 = 1'b1;
  assign CLBLM_L_X70Y112_SLICE_X105Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_A1 = CLBLM_R_X65Y105_SLICE_X98Y105_DO6;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_A2 = CLBLM_R_X65Y103_SLICE_X98Y103_A5Q;
  assign CLBLM_L_X74Y122_SLICE_X112Y122_C3 = 1'b1;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_C1 = 1'b1;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_A3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_A4 = CLBLM_R_X65Y105_SLICE_X98Y105_AO6;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_A5 = CLBLM_R_X65Y106_SLICE_X99Y106_DQ;
  assign CLBLM_L_X74Y122_SLICE_X112Y122_C4 = 1'b1;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_A6 = CLBLM_R_X65Y104_SLICE_X99Y104_CO6;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_B1 = CLBLM_L_X64Y106_SLICE_X97Y106_AQ;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_B2 = CLBLM_R_X65Y106_SLICE_X99Y106_BQ;
  assign CLBLM_L_X74Y122_SLICE_X112Y122_C5 = 1'b1;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_B3 = CLBLM_L_X64Y106_SLICE_X97Y106_B5Q;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_B4 = CLBLM_L_X64Y106_SLICE_X97Y106_C5Q;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_B6 = CLBLM_R_X65Y106_SLICE_X98Y106_CQ;
  assign CLBLM_L_X74Y122_SLICE_X112Y122_C6 = 1'b1;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_C4 = 1'b1;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_C1 = CLBLM_R_X65Y106_SLICE_X99Y106_C5Q;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_C2 = CLBLM_R_X65Y106_SLICE_X99Y106_CQ;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_C3 = CLBLM_R_X65Y106_SLICE_X99Y106_BQ;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_C5 = 1'b1;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_C4 = CLBLM_R_X63Y106_SLICE_X94Y106_AO6;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_C5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_C6 = 1'b1;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X76Y129_SLICE_X117Y129_A3 = 1'b1;
  assign CLBLM_L_X70Y112_SLICE_X105Y112_D1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_D1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y122_SLICE_X112Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X76Y129_SLICE_X117Y129_A4 = 1'b1;
  assign CLBLM_L_X70Y112_SLICE_X105Y112_D2 = CLBLM_L_X70Y112_SLICE_X105Y112_CQ;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_D2 = CLBLM_R_X65Y104_SLICE_X99Y104_CO6;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_D3 = CLBLM_R_X65Y105_SLICE_X98Y105_DO6;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_D4 = CLBLM_R_X65Y103_SLICE_X98Y103_A5Q;
  assign CLBLM_L_X76Y129_SLICE_X117Y129_A5 = 1'b1;
  assign CLBLM_L_X70Y112_SLICE_X105Y112_D3 = CLBLM_L_X70Y112_SLICE_X105Y112_DQ;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_D5 = 1'b1;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_D6 = CLBLM_R_X65Y105_SLICE_X98Y105_AO6;
  assign CLBLM_L_X76Y129_SLICE_X117Y129_A6 = 1'b1;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_A1 = 1'b1;
  assign CLBLM_L_X70Y112_SLICE_X105Y112_D4 = 1'b1;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_A2 = CLBLM_R_X65Y106_SLICE_X98Y106_BQ;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_A3 = CLBLM_R_X65Y106_SLICE_X98Y106_AQ;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_A5 = CLBLM_R_X63Y106_SLICE_X94Y106_AO6;
  assign CLBLM_L_X70Y112_SLICE_X105Y112_D5 = CLBLM_L_X70Y112_SLICE_X105Y112_B5Q;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_A6 = CLBLM_L_X62Y106_SLICE_X93Y106_DO6;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_B1 = CLBLM_L_X64Y106_SLICE_X97Y106_AQ;
  assign CLBLM_L_X70Y112_SLICE_X105Y112_D6 = 1'b1;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_B2 = CLBLM_R_X65Y106_SLICE_X98Y106_BQ;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_B4 = CLBLM_L_X64Y106_SLICE_X97Y106_B5Q;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_B5 = CLBLM_R_X65Y106_SLICE_X98Y106_DQ;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_B6 = CLBLM_L_X64Y106_SLICE_X97Y106_C5Q;
  assign RIOI3_X105Y101_OLOGIC_X1Y102_T1 = 1'b1;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_C1 = CLBLM_R_X63Y106_SLICE_X94Y106_AO6;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_C2 = CLBLM_R_X65Y106_SLICE_X98Y106_CQ;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_C3 = CLBLM_R_X65Y106_SLICE_X98Y106_AQ;
  assign CLBLM_L_X74Y122_SLICE_X112Y122_D1 = 1'b1;
  assign CLBLM_L_X76Y129_SLICE_X117Y129_B1 = 1'b1;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_C4 = CLBLM_R_X65Y106_SLICE_X98Y106_BQ;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_C5 = 1'b1;
  assign CLBLM_L_X74Y122_SLICE_X112Y122_D2 = 1'b1;
  assign CLBLM_L_X76Y129_SLICE_X117Y129_B2 = 1'b1;
  assign CLBLM_L_X70Y112_SLICE_X105Y112_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_C6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y122_SLICE_X112Y122_D3 = 1'b1;
  assign CLBLM_L_X76Y129_SLICE_X117Y129_B3 = 1'b1;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_D1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_D2 = CLBLM_L_X64Y106_SLICE_X97Y106_AQ;
  assign CLBLM_L_X74Y122_SLICE_X112Y122_D4 = 1'b1;
  assign CLBLM_L_X76Y129_SLICE_X117Y129_B4 = 1'b1;
  assign CLBLM_L_X78Y127_SLICE_X120Y127_A1 = 1'b1;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_D3 = CLBLM_R_X65Y106_SLICE_X98Y106_DQ;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_D4 = CLBLM_L_X64Y106_SLICE_X97Y106_B5Q;
  assign CLBLM_L_X74Y122_SLICE_X112Y122_D5 = 1'b1;
  assign CLBLM_L_X76Y129_SLICE_X117Y129_B5 = 1'b1;
  assign CLBLM_L_X78Y127_SLICE_X120Y127_A2 = 1'b1;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_D5 = CLBLL_R_X79Y99_SLICE_X122Y99_AO6;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_D6 = CLBLM_L_X64Y106_SLICE_X97Y106_C5Q;
  assign CLBLM_L_X74Y122_SLICE_X112Y122_D6 = 1'b1;
  assign CLBLM_L_X76Y129_SLICE_X117Y129_B6 = 1'b1;
  assign CLBLM_L_X70Y112_SLICE_X104Y112_A1 = CLBLL_R_X71Y111_SLICE_X107Y111_AQ;
  assign CLBLM_L_X78Y127_SLICE_X120Y127_A3 = 1'b1;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X78Y127_SLICE_X120Y127_A4 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_D1 = CLBLL_R_X79Y135_SLICE_X122Y135_AQ;
  assign CLBLM_L_X78Y127_SLICE_X120Y127_A5 = 1'b1;
  assign CLBLM_L_X70Y112_SLICE_X104Y112_A3 = CLBLM_L_X70Y112_SLICE_X104Y112_AQ;
  assign CLBLM_L_X78Y127_SLICE_X120Y127_A6 = 1'b1;
  assign CLBLM_L_X70Y112_SLICE_X104Y112_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y112_SLICE_X104Y112_A5 = CLBLM_L_X72Y111_SLICE_X109Y111_AQ;
  assign CLBLM_L_X74Y122_SLICE_X112Y122_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X76Y129_SLICE_X117Y129_C1 = 1'b1;
  assign CLBLM_L_X70Y112_SLICE_X104Y112_A6 = CLBLM_L_X72Y111_SLICE_X109Y111_A5Q;
  assign CLBLM_L_X76Y129_SLICE_X117Y129_C2 = 1'b1;
  assign CLBLM_L_X76Y129_SLICE_X117Y129_C3 = 1'b1;
  assign RIOI3_X105Y61_ILOGIC_X1Y62_D = RIOB33_X105Y61_IOB_X1Y62_I;
  assign CLBLM_L_X76Y129_SLICE_X117Y129_C4 = 1'b1;
  assign CLBLM_L_X76Y129_SLICE_X117Y129_C5 = 1'b1;
  assign CLBLM_L_X78Y127_SLICE_X120Y127_B1 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_B5 = CLBLM_L_X64Y102_SLICE_X96Y102_DO6;
  assign CLBLM_L_X76Y129_SLICE_X117Y129_C6 = 1'b1;
  assign CLBLM_L_X78Y127_SLICE_X120Y127_B2 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_B6 = CLBLM_R_X65Y104_SLICE_X99Y104_DO6;
  assign CLBLM_L_X78Y127_SLICE_X120Y127_B3 = 1'b1;
  assign CLBLM_L_X78Y127_SLICE_X120Y127_B4 = 1'b1;
  assign CLBLM_L_X78Y127_SLICE_X120Y127_B5 = 1'b1;
  assign CLBLM_L_X78Y127_SLICE_X120Y127_B6 = 1'b1;
  assign CLBLM_L_X70Y112_SLICE_X104Y112_B5 = CLBLM_L_X70Y112_SLICE_X104Y112_A5Q;
  assign CLBLM_L_X70Y112_SLICE_X104Y112_B6 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X163Y67_A1 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X163Y67_A2 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X163Y67_A3 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X163Y67_A4 = 1'b1;
  assign CLBLM_L_X76Y129_SLICE_X117Y129_D1 = 1'b1;
  assign CLBLM_L_X78Y127_SLICE_X120Y127_C1 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X163Y67_A5 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X163Y67_A6 = 1'b1;
  assign CLBLM_L_X76Y129_SLICE_X117Y129_D2 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X163Y67_AX = CLBLM_R_X103Y67_SLICE_X162Y67_AQ;
  assign CLBLM_R_X103Y67_SLICE_X163Y67_B1 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X163Y67_B2 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X163Y67_B3 = 1'b1;
  assign CLBLM_L_X76Y129_SLICE_X117Y129_D3 = 1'b1;
  assign CLBLM_L_X78Y127_SLICE_X120Y127_C3 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X163Y67_B4 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X163Y67_B5 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X163Y67_B6 = 1'b1;
  assign CLBLM_L_X76Y129_SLICE_X117Y129_D4 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X163Y67_BX = CLBLM_R_X103Y67_SLICE_X162Y67_CQ;
  assign CLBLM_R_X103Y67_SLICE_X163Y67_C1 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X163Y67_C2 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X163Y67_C3 = 1'b1;
  assign CLBLM_L_X76Y129_SLICE_X117Y129_D5 = 1'b1;
  assign CLBLM_L_X78Y127_SLICE_X120Y127_C5 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X163Y67_C4 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X163Y67_C5 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X163Y67_C6 = 1'b1;
  assign CLBLM_L_X76Y129_SLICE_X117Y129_D6 = 1'b1;
  assign CLBLM_L_X78Y127_SLICE_X120Y127_C6 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X163Y67_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X103Y67_SLICE_X163Y67_CX = CLBLM_R_X103Y67_SLICE_X163Y67_BQ;
  assign CLBLM_R_X103Y67_SLICE_X163Y67_D1 = 1'b1;
  assign CLBLM_L_X70Y112_SLICE_X104Y112_C5 = CLBLM_L_X70Y113_SLICE_X104Y113_BQ;
  assign CLBLM_R_X103Y67_SLICE_X163Y67_D2 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X163Y67_D3 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X163Y67_D4 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X163Y67_D5 = 1'b1;
  assign CLBLM_L_X70Y112_SLICE_X104Y112_C6 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X163Y67_D6 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X163Y67_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X103Y67_SLICE_X162Y67_A1 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X162Y67_A2 = CLBLM_R_X103Y67_SLICE_X162Y67_BQ;
  assign CLBLM_R_X103Y67_SLICE_X162Y67_A3 = CLBLM_R_X103Y67_SLICE_X162Y67_CQ;
  assign CLBLM_R_X103Y67_SLICE_X162Y67_A4 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X162Y67_A5 = CLBLM_R_X103Y67_SLICE_X162Y67_AQ;
  assign CLBLM_R_X103Y67_SLICE_X162Y67_A6 = CLBLM_R_X103Y67_SLICE_X163Y67_BQ;
  assign CLBLM_R_X103Y67_SLICE_X162Y67_AX = CLBLM_R_X103Y69_SLICE_X162Y69_AQ;
  assign CLBLM_R_X103Y67_SLICE_X162Y67_B1 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X162Y67_B2 = 1'b1;
  assign CLBLM_L_X70Y112_SLICE_X104Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X103Y67_SLICE_X162Y67_B3 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X162Y67_B4 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X162Y67_B5 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X162Y67_B6 = 1'b1;
  assign RIOB33_X105Y85_IOB_X1Y85_O = CLBLL_R_X71Y98_SLICE_X106Y98_AQ;
  assign RIOB33_X105Y85_IOB_X1Y86_O = CLBLM_L_X64Y99_SLICE_X97Y99_A5Q;
  assign CLBLM_R_X103Y67_SLICE_X162Y67_BX = CLBLM_R_X103Y67_SLICE_X163Y67_AQ;
  assign CLBLM_L_X76Y129_SLICE_X116Y129_A1 = CLBLM_L_X76Y128_SLICE_X117Y128_AQ;
  assign CLBLM_R_X103Y67_SLICE_X162Y67_C1 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X162Y67_C2 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X162Y67_C3 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X162Y67_C4 = 1'b1;
  assign CLBLM_L_X76Y129_SLICE_X116Y129_A2 = CLBLM_L_X78Y131_SLICE_X120Y131_AQ;
  assign CLBLM_R_X103Y67_SLICE_X162Y67_C5 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X162Y67_C6 = 1'b1;
  assign CLBLM_L_X76Y129_SLICE_X116Y129_A3 = CLBLL_R_X77Y129_SLICE_X119Y129_BQ;
  assign CLBLM_R_X103Y67_SLICE_X162Y67_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X76Y129_SLICE_X116Y129_A4 = CLBLL_R_X77Y130_SLICE_X118Y130_AQ;
  assign CLBLM_R_X103Y67_SLICE_X162Y67_CX = CLBLM_R_X103Y67_SLICE_X162Y67_BQ;
  assign CLBLM_R_X103Y67_SLICE_X162Y67_D1 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X162Y67_D2 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X162Y67_D3 = 1'b1;
  assign CLBLM_L_X76Y129_SLICE_X116Y129_A5 = CLBLL_R_X75Y129_SLICE_X114Y129_BQ;
  assign CLBLM_R_X103Y67_SLICE_X162Y67_D4 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X162Y67_D5 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X162Y67_D6 = 1'b1;
  assign CLBLM_L_X76Y129_SLICE_X116Y129_A6 = 1'b1;
  assign CLBLM_R_X103Y67_SLICE_X162Y67_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X78Y127_SLICE_X120Y127_D4 = 1'b1;
  assign CLBLM_L_X78Y127_SLICE_X120Y127_D5 = 1'b1;
  assign CLBLM_L_X72Y107_SLICE_X109Y107_A5 = CLBLM_L_X72Y107_SLICE_X108Y107_AQ;
  assign CLBLM_L_X70Y112_SLICE_X104Y112_D4 = CLBLM_L_X70Y110_SLICE_X104Y110_CQ;
  assign CLBLM_L_X78Y127_SLICE_X120Y127_D6 = 1'b1;
  assign CLBLM_L_X76Y129_SLICE_X116Y129_AX = CLBLM_L_X76Y129_SLICE_X116Y129_CQ;
  assign CLBLM_L_X72Y107_SLICE_X109Y107_A6 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X70Y112_SLICE_X104Y112_D5 = CLBLM_L_X70Y112_SLICE_X104Y112_BO5;
  assign CLBLM_R_X103Y75_SLICE_X162Y75_C5 = 1'b1;
  assign CLBLM_L_X76Y129_SLICE_X116Y129_B1 = CLBLL_R_X75Y130_SLICE_X115Y130_BO5;
  assign CLBLM_L_X76Y129_SLICE_X116Y129_B2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X76Y129_SLICE_X116Y129_B3 = CLBLM_L_X76Y130_SLICE_X116Y130_AQ;
  assign CLBLM_L_X76Y129_SLICE_X116Y129_B4 = CLBLM_L_X76Y129_SLICE_X116Y129_DO6;
  assign CLBLM_L_X76Y129_SLICE_X116Y129_B5 = CLBLL_R_X75Y129_SLICE_X114Y129_BQ;
  assign CLBLM_L_X76Y129_SLICE_X116Y129_B6 = CLBLM_L_X76Y129_SLICE_X116Y129_AO5;
  assign CLBLM_L_X76Y129_SLICE_X116Y129_BX = CLBLM_L_X76Y128_SLICE_X116Y128_C5Q;
  assign CLBLM_L_X72Y107_SLICE_X109Y107_BX = CLBLM_L_X72Y107_SLICE_X109Y107_A5Q;
  assign CLBLM_L_X76Y129_SLICE_X116Y129_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y133_SLICE_X105Y133_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_A1 = CLBLM_L_X72Y123_SLICE_X108Y123_CO6;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_A3 = CLBLM_L_X68Y107_SLICE_X103Y107_AO6;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_A4 = CLBLL_R_X71Y121_SLICE_X106Y121_BO6;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_A5 = CLBLM_L_X72Y118_SLICE_X108Y118_AQ;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_A6 = CLBLM_L_X68Y105_SLICE_X102Y105_DO6;
  assign CLBLM_L_X70Y133_SLICE_X105Y133_A3 = CLBLM_L_X70Y133_SLICE_X105Y133_AQ;
  assign CLBLM_L_X72Y107_SLICE_X109Y107_C1 = CLBLL_R_X71Y107_SLICE_X106Y107_CQ;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_AX = CLBLL_R_X71Y121_SLICE_X106Y121_BO5;
  assign CLBLM_L_X76Y129_SLICE_X116Y129_C2 = CLBLM_L_X76Y129_SLICE_X116Y129_CQ;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_B1 = CLBLL_R_X71Y126_SLICE_X107Y126_CO6;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_B2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_B3 = CLBLM_R_X63Y122_SLICE_X95Y122_CQ;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_B4 = CLBLL_R_X83Y94_SLICE_X130Y94_AQ;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_B5 = CLBLL_R_X71Y121_SLICE_X106Y121_A5Q;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_B6 = 1'b1;
  assign CLBLM_L_X72Y107_SLICE_X109Y107_C2 = CLBLM_L_X72Y106_SLICE_X108Y106_A5Q;
  assign CLBLM_L_X72Y107_SLICE_X109Y107_C3 = CLBLM_L_X72Y108_SLICE_X109Y108_DQ;
  assign CLBLM_L_X76Y129_SLICE_X116Y129_C4 = CLBLM_L_X76Y128_SLICE_X116Y128_C5Q;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_C1 = 1'b1;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_C2 = 1'b1;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_C3 = 1'b1;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_C4 = 1'b1;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_C5 = 1'b1;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_C6 = 1'b1;
  assign CLBLM_L_X72Y107_SLICE_X109Y107_C4 = CLBLL_R_X73Y108_SLICE_X110Y108_BQ;
  assign CLBLM_L_X72Y107_SLICE_X109Y107_C5 = CLBLM_L_X62Y90_SLICE_X92Y90_AQ;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X76Y129_SLICE_X116Y129_C6 = CLBLM_L_X76Y125_SLICE_X116Y125_BQ;
  assign CLBLM_L_X72Y107_SLICE_X109Y107_C6 = CLBLL_R_X71Y107_SLICE_X106Y107_C5Q;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_D1 = 1'b1;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_D2 = 1'b1;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_D3 = 1'b1;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_D4 = 1'b1;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_D5 = 1'b1;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_D6 = 1'b1;
  assign CLBLM_L_X76Y129_SLICE_X116Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y107_SLICE_X109Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_A1 = 1'b1;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_A2 = 1'b1;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_A3 = 1'b1;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_A4 = 1'b1;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_A5 = 1'b1;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_A6 = 1'b1;
  assign CLBLM_L_X76Y129_SLICE_X116Y129_D1 = CLBLM_L_X76Y127_SLICE_X116Y127_AQ;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_B1 = 1'b1;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_B2 = 1'b1;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_B3 = 1'b1;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_B4 = 1'b1;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_B5 = 1'b1;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_B6 = 1'b1;
  assign CLBLM_L_X72Y107_SLICE_X109Y107_D1 = CLBLM_L_X72Y106_SLICE_X108Y106_AQ;
  assign CLBLM_L_X72Y107_SLICE_X109Y107_D2 = CLBLM_L_X72Y106_SLICE_X108Y106_A5Q;
  assign CLBLM_L_X76Y129_SLICE_X116Y129_D2 = CLBLM_L_X76Y130_SLICE_X116Y130_BQ;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_C1 = 1'b1;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_C2 = 1'b1;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_C3 = 1'b1;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_C4 = 1'b1;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_C5 = 1'b1;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_C6 = 1'b1;
  assign CLBLM_L_X72Y107_SLICE_X109Y107_D3 = CLBLM_L_X62Y90_SLICE_X92Y90_AQ;
  assign CLBLM_L_X72Y107_SLICE_X109Y107_D4 = 1'b1;
  assign CLBLM_L_X76Y129_SLICE_X116Y129_D4 = CLBLM_L_X76Y130_SLICE_X116Y130_A5Q;
  assign CLBLM_L_X76Y129_SLICE_X116Y129_D5 = CLBLM_L_X76Y129_SLICE_X116Y129_BQ;
  assign CLBLM_L_X76Y129_SLICE_X116Y129_D6 = CLBLL_R_X77Y128_SLICE_X118Y128_CQ;
  assign CLBLM_L_X72Y107_SLICE_X109Y107_D5 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_A2 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_A4 = 1'b1;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_D1 = 1'b1;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_D2 = 1'b1;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_D3 = 1'b1;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_D4 = 1'b1;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_D5 = 1'b1;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_D6 = 1'b1;
  assign CLBLM_L_X72Y107_SLICE_X109Y107_D6 = CLBLM_L_X78Y106_SLICE_X120Y106_AQ;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_B2 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_B4 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_B5 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_B6 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_C1 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_C2 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_C3 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_C4 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_C5 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_C6 = 1'b1;
  assign CLBLM_L_X72Y107_SLICE_X109Y107_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X76Y129_SLICE_X116Y129_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_D1 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_D2 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_D3 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_D4 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_D5 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_D6 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_A1 = CLBLM_L_X78Y121_SLICE_X120Y121_CO6;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_A2 = CLBLM_L_X78Y122_SLICE_X121Y122_AQ;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_A3 = CLBLM_L_X78Y120_SLICE_X120Y120_AQ;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_A4 = CLBLM_L_X76Y122_SLICE_X117Y122_AQ;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_A5 = CLBLL_R_X77Y113_SLICE_X118Y113_AQ;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_A6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_B1 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_B2 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_B3 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_B4 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_B5 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_B6 = 1'b1;
  assign RIOB33_X105Y87_IOB_X1Y88_O = CLBLM_L_X68Y105_SLICE_X102Y105_AQ;
  assign RIOB33_X105Y87_IOB_X1Y87_O = CLBLM_L_X64Y97_SLICE_X97Y97_AQ;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_C1 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_C2 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_C3 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_C4 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_C5 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_C6 = 1'b1;
  assign CLBLM_R_X67Y118_SLICE_X101Y118_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_D1 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_D2 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_D3 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_D4 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_D5 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_D6 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y107_SLICE_X108Y107_B6 = 1'b1;
  assign CLBLM_L_X72Y107_SLICE_X108Y107_BX = CLBLM_L_X72Y107_SLICE_X108Y107_A5Q;
  assign CLBLM_R_X65Y108_SLICE_X99Y108_A1 = CLBLM_R_X65Y109_SLICE_X98Y109_DO6;
  assign CLBLM_R_X65Y108_SLICE_X99Y108_A2 = CLBLM_R_X65Y108_SLICE_X98Y108_BO6;
  assign CLBLM_R_X65Y108_SLICE_X99Y108_A3 = CLBLM_R_X65Y108_SLICE_X98Y108_AO6;
  assign CLBLM_R_X65Y108_SLICE_X99Y108_A4 = CLBLM_R_X65Y108_SLICE_X99Y108_BO6;
  assign CLBLM_R_X65Y108_SLICE_X99Y108_A5 = CLBLM_R_X65Y108_SLICE_X99Y108_CO6;
  assign CLBLM_R_X65Y108_SLICE_X99Y108_A6 = CLBLM_R_X65Y109_SLICE_X99Y109_DO5;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_D1 = 1'b1;
  assign CLBLM_R_X65Y108_SLICE_X99Y108_B1 = CLBLM_L_X68Y108_SLICE_X102Y108_A5Q;
  assign CLBLM_R_X65Y108_SLICE_X99Y108_B2 = CLBLM_R_X65Y109_SLICE_X98Y109_A5Q;
  assign CLBLM_R_X65Y108_SLICE_X99Y108_B3 = CLBLM_L_X68Y108_SLICE_X102Y108_AQ;
  assign CLBLM_R_X65Y108_SLICE_X99Y108_B4 = CLBLM_R_X65Y110_SLICE_X99Y110_BQ;
  assign CLBLM_R_X65Y108_SLICE_X99Y108_B5 = CLBLM_R_X67Y109_SLICE_X101Y109_BQ;
  assign CLBLM_R_X65Y108_SLICE_X99Y108_B6 = CLBLM_R_X65Y110_SLICE_X98Y110_A5Q;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_T1 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_D1 = 1'b0;
  assign CLBLM_R_X65Y108_SLICE_X99Y108_C1 = CLBLM_R_X65Y110_SLICE_X99Y110_CQ;
  assign CLBLM_R_X65Y108_SLICE_X99Y108_C2 = CLBLM_L_X68Y108_SLICE_X102Y108_AQ;
  assign CLBLM_R_X65Y108_SLICE_X99Y108_C3 = CLBLM_R_X65Y109_SLICE_X99Y109_BQ;
  assign CLBLM_R_X65Y108_SLICE_X99Y108_C4 = CLBLM_L_X68Y108_SLICE_X102Y108_A5Q;
  assign CLBLM_R_X65Y108_SLICE_X99Y108_C5 = CLBLM_L_X68Y109_SLICE_X102Y109_A5Q;
  assign CLBLM_R_X65Y108_SLICE_X99Y108_C6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_D1 = 1'b1;
  assign CLBLM_L_X72Y107_SLICE_X108Y107_C5 = CLBLM_L_X72Y107_SLICE_X108Y107_DO6;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_T1 = 1'b1;
  assign CLBLM_L_X72Y107_SLICE_X108Y107_C6 = CLBLM_L_X72Y107_SLICE_X108Y107_BO6;
  assign CLBLM_R_X65Y108_SLICE_X99Y108_D1 = 1'b1;
  assign CLBLM_R_X65Y108_SLICE_X99Y108_D2 = 1'b1;
  assign CLBLM_R_X65Y108_SLICE_X99Y108_D3 = 1'b1;
  assign CLBLM_R_X65Y108_SLICE_X99Y108_D4 = 1'b1;
  assign CLBLM_R_X65Y108_SLICE_X99Y108_D5 = 1'b1;
  assign CLBLM_R_X65Y108_SLICE_X99Y108_D6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_T1 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_D1 = CLBLL_R_X71Y117_SLICE_X106Y117_A5Q;
  assign RIOI3_X105Y65_OLOGIC_X1Y66_D1 = CLBLM_R_X103Y67_SLICE_X162Y67_CQ;
  assign CLBLM_R_X65Y108_SLICE_X98Y108_A1 = CLBLM_R_X65Y110_SLICE_X98Y110_A5Q;
  assign CLBLM_R_X65Y108_SLICE_X98Y108_A2 = CLBLM_L_X68Y108_SLICE_X102Y108_A5Q;
  assign CLBLM_R_X65Y108_SLICE_X98Y108_A3 = CLBLM_R_X65Y111_SLICE_X98Y111_AQ;
  assign CLBLM_R_X65Y108_SLICE_X98Y108_A4 = CLBLM_R_X65Y110_SLICE_X98Y110_BQ;
  assign CLBLM_L_X72Y107_SLICE_X108Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X65Y108_SLICE_X98Y108_A5 = CLBLM_L_X68Y108_SLICE_X102Y108_AQ;
  assign CLBLM_R_X65Y108_SLICE_X98Y108_A6 = CLBLM_R_X65Y109_SLICE_X98Y109_CQ;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_T1 = 1'b1;
  assign CLBLM_R_X65Y108_SLICE_X98Y108_B1 = CLBLM_R_X65Y109_SLICE_X99Y109_CQ;
  assign CLBLM_R_X65Y108_SLICE_X98Y108_B2 = CLBLM_L_X68Y108_SLICE_X102Y108_A5Q;
  assign CLBLM_R_X65Y108_SLICE_X98Y108_B3 = CLBLM_R_X65Y109_SLICE_X98Y109_A5Q;
  assign CLBLM_R_X65Y108_SLICE_X98Y108_B4 = CLBLM_L_X68Y108_SLICE_X102Y108_AQ;
  assign CLBLM_R_X65Y108_SLICE_X98Y108_B5 = CLBLM_L_X62Y92_SLICE_X92Y92_BQ;
  assign CLBLM_R_X65Y108_SLICE_X98Y108_B6 = CLBLM_R_X65Y110_SLICE_X98Y110_AQ;
  assign RIOI3_X105Y65_OLOGIC_X1Y66_T1 = 1'b1;
  assign CLBLM_R_X65Y108_SLICE_X98Y108_C1 = 1'b1;
  assign CLBLM_R_X65Y108_SLICE_X98Y108_C2 = 1'b1;
  assign CLBLM_R_X65Y108_SLICE_X98Y108_C3 = 1'b1;
  assign CLBLM_R_X65Y108_SLICE_X98Y108_C4 = 1'b1;
  assign CLBLM_R_X65Y108_SLICE_X98Y108_C5 = 1'b1;
  assign CLBLM_R_X65Y108_SLICE_X98Y108_C6 = 1'b1;
  assign RIOI3_X105Y65_OLOGIC_X1Y65_D1 = CLBLM_R_X103Y67_SLICE_X162Y67_BQ;
  assign CLBLM_L_X74Y103_SLICE_X112Y103_D4 = CLBLM_L_X72Y104_SLICE_X109Y104_BQ;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_D1 = CLBLM_L_X62Y106_SLICE_X93Y106_AQ;
  assign RIOI3_X105Y65_OLOGIC_X1Y65_T1 = 1'b1;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1 = CLBLM_L_X74Y109_SLICE_X113Y109_AQ;
  assign CLBLM_R_X65Y108_SLICE_X98Y108_D1 = 1'b1;
  assign CLBLM_R_X65Y108_SLICE_X98Y108_D2 = 1'b1;
  assign CLBLM_R_X65Y108_SLICE_X98Y108_D3 = 1'b1;
  assign CLBLM_R_X65Y108_SLICE_X98Y108_D4 = 1'b1;
  assign CLBLM_R_X65Y108_SLICE_X98Y108_D5 = 1'b1;
  assign CLBLM_R_X65Y108_SLICE_X98Y108_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_T1 = 1'b1;
  assign CLBLM_L_X72Y107_SLICE_X108Y107_D4 = CLBLL_R_X71Y107_SLICE_X107Y107_BQ;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_D1 = CLBLM_L_X76Y128_SLICE_X116Y128_CQ;
  assign CLBLM_L_X72Y107_SLICE_X108Y107_D5 = CLBLM_L_X78Y106_SLICE_X120Y106_AQ;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_T1 = 1'b1;
  assign LIOB33_X0Y163_IOB_X0Y164_O = CLBLL_R_X73Y123_SLICE_X110Y123_AQ;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_D1 = CLBLL_R_X73Y103_SLICE_X110Y103_B5Q;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1 = 1'b1;
  assign LIOB33_X0Y163_IOB_X0Y163_O = CLBLM_R_X63Y106_SLICE_X95Y106_AQ;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_A1 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_A2 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_A3 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_A4 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_A5 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_A6 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_B1 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_B2 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_B3 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_B4 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_B5 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_B6 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_C1 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_C2 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_C3 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_C4 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_C5 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_C6 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_D1 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_D2 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_D3 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_D4 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_D5 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_D6 = 1'b1;
  assign CLBLM_R_X103Y69_SLICE_X163Y69_A1 = 1'b1;
  assign CLBLM_R_X103Y69_SLICE_X163Y69_A2 = 1'b1;
  assign CLBLM_R_X103Y69_SLICE_X163Y69_A3 = 1'b1;
  assign CLBLM_R_X103Y69_SLICE_X163Y69_A4 = 1'b1;
  assign CLBLM_R_X103Y69_SLICE_X163Y69_A5 = 1'b1;
  assign CLBLM_R_X103Y69_SLICE_X163Y69_A6 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_A2 = CLBLM_L_X78Y123_SLICE_X121Y123_BQ;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_A3 = CLBLM_L_X78Y121_SLICE_X120Y121_AQ;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_A4 = CLBLM_L_X78Y123_SLICE_X120Y123_BO6;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_A5 = CLBLL_R_X77Y113_SLICE_X118Y113_AQ;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_A6 = CLBLM_L_X76Y122_SLICE_X117Y122_AQ;
  assign CLBLM_R_X103Y69_SLICE_X163Y69_AX = CLBLM_R_X103Y67_SLICE_X163Y67_CQ;
  assign CLBLM_R_X103Y69_SLICE_X163Y69_B1 = 1'b1;
  assign CLBLM_R_X103Y69_SLICE_X163Y69_B2 = 1'b1;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_A6 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_B1 = CLBLM_L_X78Y123_SLICE_X120Y123_BO6;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_B2 = CLBLM_L_X78Y121_SLICE_X120Y121_BQ;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_B3 = CLBLM_L_X78Y121_SLICE_X120Y121_AQ;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_B4 = CLBLM_L_X76Y122_SLICE_X117Y122_AQ;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_B5 = CLBLL_R_X77Y113_SLICE_X118Y113_AQ;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_B6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X103Y69_SLICE_X163Y69_B6 = 1'b1;
  assign CLBLM_R_X103Y69_SLICE_X163Y69_C1 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_B2 = 1'b1;
  assign CLBLM_R_X103Y69_SLICE_X163Y69_C3 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_C1 = CLBLL_R_X77Y113_SLICE_X118Y113_AQ;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_C2 = CLBLM_L_X78Y121_SLICE_X120Y121_AQ;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_C3 = CLBLM_L_X78Y121_SLICE_X120Y121_BQ;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_C4 = CLBLM_L_X76Y122_SLICE_X117Y122_AQ;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_C5 = CLBLM_L_X78Y123_SLICE_X120Y123_BO6;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_C6 = 1'b1;
  assign CLBLM_R_X103Y69_SLICE_X163Y69_D1 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X103Y69_SLICE_X163Y69_D2 = 1'b1;
  assign CLBLM_R_X103Y69_SLICE_X163Y69_D3 = 1'b1;
  assign CLBLM_R_X103Y69_SLICE_X163Y69_D4 = 1'b1;
  assign CLBLM_R_X103Y69_SLICE_X163Y69_D5 = 1'b1;
  assign CLBLM_R_X103Y69_SLICE_X163Y69_D6 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_D1 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_D2 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_D3 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_D4 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_D5 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_D6 = 1'b1;
  assign CLBLM_R_X103Y69_SLICE_X162Y69_A1 = 1'b1;
  assign CLBLM_R_X103Y69_SLICE_X162Y69_A2 = CLBLM_R_X103Y67_SLICE_X162Y67_CQ;
  assign CLBLM_R_X103Y69_SLICE_X162Y69_A3 = CLBLL_R_X83Y94_SLICE_X130Y94_AQ;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X103Y69_SLICE_X162Y69_A4 = CLBLM_R_X103Y69_SLICE_X162Y69_BO6;
  assign CLBLM_R_X103Y69_SLICE_X162Y69_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X103Y69_SLICE_X162Y69_A6 = CLBLM_R_X103Y69_SLICE_X162Y69_A5Q;
  assign CLBLM_R_X103Y69_SLICE_X162Y69_AX = CLBLM_R_X103Y69_SLICE_X163Y69_AQ;
  assign CLBLM_R_X103Y69_SLICE_X162Y69_B1 = CLBLM_R_X103Y67_SLICE_X163Y67_AQ;
  assign CLBLM_R_X103Y69_SLICE_X162Y69_B2 = CLBLM_R_X103Y67_SLICE_X162Y67_AO6;
  assign CLBLM_R_X103Y69_SLICE_X162Y69_B3 = CLBLM_R_X103Y69_SLICE_X162Y69_AQ;
  assign CLBLM_R_X103Y69_SLICE_X162Y69_B4 = CLBLM_R_X103Y69_SLICE_X163Y69_AQ;
  assign CLBLM_R_X103Y69_SLICE_X162Y69_B5 = CLBLM_R_X103Y67_SLICE_X163Y67_CQ;
  assign CLBLM_R_X103Y69_SLICE_X162Y69_B6 = CLBLM_R_X103Y69_SLICE_X162Y69_A5Q;
  assign CLBLM_R_X103Y69_SLICE_X162Y69_C1 = 1'b1;
  assign CLBLM_R_X103Y69_SLICE_X162Y69_C2 = 1'b1;
  assign CLBLM_R_X103Y69_SLICE_X162Y69_C3 = 1'b1;
  assign CLBLM_R_X103Y69_SLICE_X162Y69_C4 = 1'b1;
  assign CLBLM_L_X76Y134_SLICE_X117Y134_D2 = 1'b1;
  assign CLBLM_R_X103Y69_SLICE_X162Y69_C5 = 1'b1;
  assign CLBLM_R_X103Y69_SLICE_X162Y69_C6 = 1'b1;
  assign CLBLM_R_X103Y69_SLICE_X163Y69_C6 = 1'b1;
  assign CLBLM_R_X103Y69_SLICE_X162Y69_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X103Y69_SLICE_X162Y69_D1 = 1'b1;
  assign CLBLM_R_X103Y69_SLICE_X162Y69_D2 = 1'b1;
  assign CLBLM_R_X103Y69_SLICE_X162Y69_D3 = 1'b1;
  assign CLBLM_R_X103Y69_SLICE_X162Y69_D4 = 1'b1;
  assign CLBLM_R_X103Y69_SLICE_X162Y69_D5 = 1'b1;
  assign CLBLM_R_X103Y69_SLICE_X162Y69_D6 = 1'b1;
  assign CLBLM_R_X103Y69_SLICE_X163Y69_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X67Y115_SLICE_X100Y115_D3 = 1'b1;
  assign CLBLM_R_X103Y69_SLICE_X162Y69_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_A2 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X67Y118_SLICE_X100Y118_B1 = 1'b1;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_A3 = CLBLM_R_X63Y103_SLICE_X95Y103_AQ;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_A4 = CLBLM_L_X64Y105_SLICE_X96Y105_CQ;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_A5 = CLBLM_R_X63Y102_SLICE_X95Y102_AO5;
  assign CLBLM_R_X65Y109_SLICE_X99Y109_A1 = CLBLM_R_X65Y109_SLICE_X99Y109_AQ;
  assign CLBLM_R_X65Y109_SLICE_X99Y109_A2 = CLBLM_R_X67Y111_SLICE_X101Y111_CO6;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_A6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y109_SLICE_X99Y109_A3 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X65Y109_SLICE_X99Y109_A4 = CLBLM_R_X67Y111_SLICE_X100Y111_A5Q;
  assign CLBLM_R_X65Y109_SLICE_X99Y109_A5 = CLBLM_R_X67Y111_SLICE_X101Y111_A5Q;
  assign CLBLM_R_X65Y109_SLICE_X99Y109_A6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y109_SLICE_X99Y109_AX = CLBLM_R_X65Y109_SLICE_X98Y109_A5Q;
  assign CLBLM_R_X65Y109_SLICE_X99Y109_B1 = CLBLM_R_X67Y111_SLICE_X101Y111_DO6;
  assign CLBLM_R_X65Y109_SLICE_X99Y109_B2 = CLBLM_R_X65Y109_SLICE_X99Y109_BQ;
  assign CLBLM_R_X65Y109_SLICE_X99Y109_B3 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X65Y109_SLICE_X99Y109_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y109_SLICE_X99Y109_B5 = CLBLM_R_X65Y111_SLICE_X99Y111_AO6;
  assign CLBLM_R_X65Y109_SLICE_X99Y109_B6 = CLBLM_R_X65Y109_SLICE_X98Y109_CQ;
  assign CLBLM_R_X65Y109_SLICE_X99Y109_C1 = CLBLM_R_X65Y111_SLICE_X99Y111_AO6;
  assign CLBLM_R_X65Y109_SLICE_X99Y109_C2 = CLBLM_R_X65Y109_SLICE_X99Y109_CQ;
  assign CLBLM_R_X65Y109_SLICE_X99Y109_C3 = CLBLM_R_X67Y111_SLICE_X101Y111_DO5;
  assign CLBLM_R_X65Y109_SLICE_X99Y109_C4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y109_SLICE_X99Y109_C5 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X65Y109_SLICE_X99Y109_C6 = CLBLM_R_X65Y109_SLICE_X99Y109_BQ;
  assign CLBLM_R_X65Y109_SLICE_X99Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X65Y109_SLICE_X99Y109_D1 = CLBLM_L_X68Y108_SLICE_X102Y108_AQ;
  assign CLBLM_R_X65Y109_SLICE_X99Y109_D2 = CLBLM_L_X68Y109_SLICE_X102Y109_A5Q;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_B3 = 1'b1;
  assign CLBLM_R_X65Y109_SLICE_X99Y109_D3 = CLBLM_L_X68Y108_SLICE_X102Y108_A5Q;
  assign CLBLM_R_X65Y109_SLICE_X99Y109_D4 = CLBLM_R_X65Y109_SLICE_X99Y109_AQ;
  assign CLBLM_R_X65Y109_SLICE_X99Y109_D5 = CLBLM_R_X65Y110_SLICE_X99Y110_AQ;
  assign CLBLM_R_X65Y109_SLICE_X99Y109_D6 = 1'b1;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_B4 = CLBLM_L_X64Y105_SLICE_X96Y105_C5Q;
  assign CLBLM_R_X65Y109_SLICE_X99Y109_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X103Y69_SLICE_X163Y69_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_B5 = CLBLM_L_X64Y105_SLICE_X96Y105_CQ;
  assign CLBLM_R_X65Y109_SLICE_X98Y109_A1 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X65Y109_SLICE_X98Y109_A2 = CLBLM_R_X65Y111_SLICE_X99Y111_AO6;
  assign CLBLM_R_X65Y109_SLICE_X98Y109_A3 = CLBLM_R_X65Y109_SLICE_X98Y109_AQ;
  assign CLBLM_R_X65Y109_SLICE_X98Y109_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y109_SLICE_X98Y109_A5 = CLBLM_R_X65Y110_SLICE_X98Y110_AQ;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_B6 = 1'b1;
  assign CLBLM_R_X65Y109_SLICE_X98Y109_A6 = CLBLM_R_X67Y111_SLICE_X101Y111_CO6;
  assign CLBLM_R_X65Y109_SLICE_X98Y109_AX = CLBLM_R_X65Y110_SLICE_X99Y110_CQ;
  assign CLBLM_R_X65Y109_SLICE_X98Y109_B1 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X65Y109_SLICE_X98Y109_B2 = CLBLM_R_X65Y109_SLICE_X98Y109_BQ;
  assign CLBLM_R_X65Y109_SLICE_X98Y109_B3 = CLBLM_R_X67Y111_SLICE_X101Y111_B5Q;
  assign CLBLM_R_X65Y109_SLICE_X98Y109_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y109_SLICE_X98Y109_B5 = CLBLM_R_X65Y111_SLICE_X99Y111_AO6;
  assign CLBLM_R_X65Y109_SLICE_X98Y109_B6 = CLBLM_R_X65Y109_SLICE_X99Y109_CQ;
  assign CLBLM_R_X65Y109_SLICE_X98Y109_C1 = CLBLM_R_X65Y111_SLICE_X99Y111_AO6;
  assign CLBLM_R_X65Y109_SLICE_X98Y109_C2 = CLBLM_R_X65Y109_SLICE_X98Y109_CQ;
  assign CLBLM_R_X65Y109_SLICE_X98Y109_C3 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X65Y109_SLICE_X98Y109_C4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y109_SLICE_X98Y109_C5 = CLBLM_R_X67Y111_SLICE_X101Y111_CO5;
  assign CLBLM_R_X65Y109_SLICE_X98Y109_C6 = CLBLM_R_X65Y109_SLICE_X98Y109_AQ;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_C1 = CLBLM_L_X62Y103_SLICE_X92Y103_B5Q;
  assign CLBLM_R_X65Y109_SLICE_X98Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_C2 = CLBLM_L_X64Y102_SLICE_X96Y102_CQ;
  assign CLBLM_R_X65Y109_SLICE_X98Y109_D1 = CLBLM_L_X68Y108_SLICE_X102Y108_AQ;
  assign CLBLM_R_X65Y109_SLICE_X98Y109_D2 = CLBLM_R_X65Y109_SLICE_X99Y109_A5Q;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_C3 = CLBLM_L_X64Y101_SLICE_X96Y101_B5Q;
  assign CLBLM_R_X65Y109_SLICE_X98Y109_D3 = CLBLM_R_X65Y109_SLICE_X98Y109_AQ;
  assign CLBLM_R_X65Y109_SLICE_X98Y109_D4 = CLBLM_R_X65Y110_SLICE_X99Y110_AQ;
  assign CLBLM_R_X65Y109_SLICE_X98Y109_D5 = CLBLM_R_X65Y109_SLICE_X98Y109_BQ;
  assign CLBLM_R_X65Y109_SLICE_X98Y109_D6 = CLBLM_L_X68Y108_SLICE_X102Y108_A5Q;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_C4 = CLBLM_L_X64Y101_SLICE_X96Y101_A5Q;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_B1 = 1'b1;
  assign CLBLM_R_X65Y109_SLICE_X98Y109_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_C5 = 1'b1;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_C6 = CLBLM_L_X64Y101_SLICE_X96Y101_BQ;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_A3 = CLBLM_L_X72Y128_SLICE_X108Y128_AQ;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_A4 = CLBLM_L_X72Y127_SLICE_X108Y127_BO6;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_A5 = CLBLM_L_X72Y126_SLICE_X108Y126_CO6;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_D1 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_B2 = CLBLM_L_X72Y128_SLICE_X108Y128_A5Q;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_A1 = CLBLM_L_X76Y122_SLICE_X117Y122_AQ;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_A2 = CLBLM_L_X78Y121_SLICE_X120Y121_BQ;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_A3 = CLBLM_L_X78Y122_SLICE_X121Y122_AQ;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_B3 = CLBLM_L_X72Y127_SLICE_X108Y127_AQ;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_A4 = CLBLM_L_X78Y121_SLICE_X120Y121_CO6;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_A5 = CLBLL_R_X77Y113_SLICE_X118Y113_AQ;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_A6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_D2 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_B2 = CLBLM_L_X78Y122_SLICE_X121Y122_BQ;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_B3 = CLBLM_L_X78Y122_SLICE_X121Y122_AQ;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_B5 = CLBLM_L_X72Y126_SLICE_X108Y126_CO6;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_B4 = CLBLM_L_X78Y123_SLICE_X121Y123_CO6;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_B5 = CLBLM_L_X78Y121_SLICE_X120Y121_CO6;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_B6 = CLBLM_L_X78Y120_SLICE_X120Y120_AQ;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_D4 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_B6 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_C1 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_C2 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_C3 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_C4 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_C5 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_C6 = 1'b1;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_D6 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_D1 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_D2 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_D3 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_D4 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_D5 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_D6 = 1'b1;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y98_SLICE_X109Y98_A1 = 1'b1;
  assign CLBLM_L_X72Y98_SLICE_X109Y98_A2 = 1'b1;
  assign CLBLM_L_X72Y98_SLICE_X109Y98_A3 = 1'b1;
  assign CLBLM_L_X72Y98_SLICE_X109Y98_A4 = 1'b1;
  assign CLBLM_L_X72Y98_SLICE_X109Y98_A5 = 1'b1;
  assign CLBLM_L_X72Y98_SLICE_X109Y98_A6 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_A1 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_A2 = CLBLM_L_X76Y122_SLICE_X117Y122_AQ;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_A3 = CLBLM_L_X78Y120_SLICE_X120Y120_AQ;
  assign CLBLM_L_X72Y98_SLICE_X109Y98_B1 = 1'b1;
  assign CLBLM_L_X72Y98_SLICE_X109Y98_B2 = 1'b1;
  assign CLBLM_L_X72Y98_SLICE_X109Y98_B3 = 1'b1;
  assign CLBLM_L_X72Y98_SLICE_X109Y98_B4 = 1'b1;
  assign CLBLM_L_X72Y98_SLICE_X109Y98_B5 = 1'b1;
  assign CLBLM_L_X72Y98_SLICE_X109Y98_B6 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_B2 = CLBLL_R_X75Y121_SLICE_X114Y121_AQ;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_B1 = CLBLM_L_X78Y123_SLICE_X121Y123_CO6;
  assign CLBLM_L_X72Y98_SLICE_X109Y98_C1 = 1'b1;
  assign CLBLM_L_X72Y98_SLICE_X109Y98_C2 = 1'b1;
  assign CLBLM_L_X72Y98_SLICE_X109Y98_C3 = 1'b1;
  assign CLBLM_L_X72Y98_SLICE_X109Y98_C4 = 1'b1;
  assign CLBLM_L_X72Y98_SLICE_X109Y98_C5 = 1'b1;
  assign CLBLM_L_X72Y98_SLICE_X109Y98_C6 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_C1 = CLBLM_L_X78Y122_SLICE_X120Y122_AO6;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_C2 = CLBLM_L_X78Y120_SLICE_X120Y120_AQ;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_A1 = CLBLL_R_X75Y128_SLICE_X114Y128_DO6;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_C3 = CLBLM_L_X78Y121_SLICE_X120Y121_BQ;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_C4 = CLBLM_L_X78Y123_SLICE_X120Y123_CO6;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_C5 = CLBLL_R_X77Y122_SLICE_X119Y122_AO5;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_C6 = CLBLM_L_X78Y122_SLICE_X121Y122_BQ;
  assign CLBLM_L_X72Y98_SLICE_X109Y98_D1 = 1'b1;
  assign CLBLM_L_X72Y98_SLICE_X109Y98_D2 = 1'b1;
  assign CLBLM_L_X72Y98_SLICE_X109Y98_D3 = 1'b1;
  assign CLBLM_L_X72Y98_SLICE_X109Y98_D4 = 1'b1;
  assign CLBLM_L_X72Y98_SLICE_X109Y98_D5 = 1'b1;
  assign CLBLM_L_X72Y98_SLICE_X109Y98_D6 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_D1 = CLBLL_R_X77Y122_SLICE_X119Y122_BQ;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_D2 = CLBLM_L_X78Y123_SLICE_X120Y123_CO6;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_D3 = CLBLM_L_X78Y121_SLICE_X120Y121_BQ;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_D4 = CLBLM_L_X78Y122_SLICE_X120Y122_AO5;
  assign CLBLM_L_X72Y98_SLICE_X108Y98_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y98_SLICE_X108Y98_A2 = 1'b1;
  assign CLBLM_L_X72Y98_SLICE_X108Y98_A3 = CLBLM_L_X72Y98_SLICE_X108Y98_AQ;
  assign CLBLM_L_X72Y98_SLICE_X108Y98_A4 = CLBLL_R_X71Y98_SLICE_X106Y98_AQ;
  assign CLBLM_L_X72Y98_SLICE_X108Y98_A5 = CLBLM_L_X72Y118_SLICE_X108Y118_D5Q;
  assign CLBLM_L_X72Y98_SLICE_X108Y98_A6 = CLBLM_L_X72Y98_SLICE_X108Y98_A5Q;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_A2 = CLBLM_L_X74Y128_SLICE_X112Y128_BQ;
  assign CLBLM_L_X72Y98_SLICE_X108Y98_AX = CLBLM_L_X72Y118_SLICE_X108Y118_D5Q;
  assign CLBLM_L_X72Y98_SLICE_X108Y98_B1 = CLBLM_L_X72Y98_SLICE_X108Y98_B5Q;
  assign CLBLM_L_X72Y98_SLICE_X108Y98_B2 = CLBLM_L_X72Y98_SLICE_X108Y98_BQ;
  assign CLBLM_L_X72Y98_SLICE_X108Y98_B3 = CLBLM_L_X68Y98_SLICE_X103Y98_AQ;
  assign CLBLM_L_X72Y98_SLICE_X108Y98_B4 = CLBLM_L_X72Y119_SLICE_X108Y119_C5Q;
  assign CLBLM_L_X72Y98_SLICE_X108Y98_B5 = 1'b1;
  assign CLBLM_L_X72Y98_SLICE_X108Y98_B6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_AX = CLBLM_L_X62Y103_SLICE_X92Y103_B5Q;
  assign CLBLM_L_X72Y98_SLICE_X108Y98_BX = CLBLM_L_X72Y119_SLICE_X108Y119_C5Q;
  assign CLBLM_L_X72Y98_SLICE_X108Y98_C1 = 1'b1;
  assign CLBLM_L_X72Y98_SLICE_X108Y98_C2 = 1'b1;
  assign CLBLM_L_X72Y98_SLICE_X108Y98_C3 = 1'b1;
  assign CLBLM_L_X72Y98_SLICE_X108Y98_C4 = 1'b1;
  assign CLBLM_L_X72Y98_SLICE_X108Y98_C5 = 1'b1;
  assign CLBLM_L_X72Y98_SLICE_X108Y98_C6 = 1'b1;
  assign CLBLM_L_X72Y98_SLICE_X108Y98_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_A3 = CLBLM_L_X74Y128_SLICE_X112Y128_AQ;
  assign CLBLM_L_X72Y98_SLICE_X108Y98_D1 = 1'b1;
  assign CLBLM_L_X72Y98_SLICE_X108Y98_D2 = 1'b1;
  assign CLBLM_L_X72Y98_SLICE_X108Y98_D3 = 1'b1;
  assign CLBLM_L_X72Y98_SLICE_X108Y98_D4 = 1'b1;
  assign CLBLM_L_X72Y98_SLICE_X108Y98_D5 = 1'b1;
  assign CLBLM_L_X72Y98_SLICE_X108Y98_D6 = 1'b1;
  assign CLBLM_L_X72Y98_SLICE_X108Y98_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_A4 = CLBLM_L_X74Y127_SLICE_X113Y127_A5Q;
  assign CLBLM_R_X65Y110_SLICE_X99Y110_A1 = CLBLM_R_X67Y111_SLICE_X101Y111_A5Q;
  assign CLBLM_R_X65Y110_SLICE_X99Y110_A2 = CLBLM_R_X67Y111_SLICE_X100Y111_A5Q;
  assign CLBLM_R_X65Y110_SLICE_X99Y110_A3 = 1'b1;
  assign CLBLM_R_X65Y110_SLICE_X99Y110_A4 = 1'b1;
  assign CLBLM_R_X65Y110_SLICE_X99Y110_A5 = 1'b1;
  assign CLBLM_R_X65Y110_SLICE_X99Y110_A6 = 1'b1;
  assign CLBLM_R_X65Y110_SLICE_X99Y110_AX = CLBLM_L_X62Y92_SLICE_X92Y92_BQ;
  assign CLBLM_R_X65Y110_SLICE_X99Y110_B1 = CLBLM_R_X67Y111_SLICE_X101Y111_CO5;
  assign CLBLM_R_X65Y110_SLICE_X99Y110_B2 = CLBLM_R_X65Y110_SLICE_X99Y110_BQ;
  assign CLBLM_R_X65Y110_SLICE_X99Y110_B3 = CLBLM_R_X65Y109_SLICE_X99Y109_AQ;
  assign CLBLM_R_X65Y110_SLICE_X99Y110_B4 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X65Y110_SLICE_X99Y110_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y110_SLICE_X99Y110_B6 = CLBLM_R_X65Y110_SLICE_X99Y110_AO5;
  assign CLBLM_R_X65Y110_SLICE_X99Y110_BX = CLBLM_L_X76Y111_SLICE_X116Y111_AQ;
  assign CLBLM_R_X65Y110_SLICE_X99Y110_C1 = CLBLM_R_X67Y110_SLICE_X100Y110_DO6;
  assign CLBLM_R_X65Y110_SLICE_X99Y110_C2 = CLBLM_L_X76Y111_SLICE_X116Y111_AQ;
  assign CLBLM_R_X65Y110_SLICE_X99Y110_C3 = CLBLM_R_X65Y109_SLICE_X99Y109_DO6;
  assign CLBLM_R_X65Y110_SLICE_X99Y110_C4 = CLBLM_R_X65Y110_SLICE_X98Y110_CQ;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y110_SLICE_X99Y110_C5 = CLBLM_R_X65Y110_SLICE_X99Y110_DO6;
  assign CLBLM_R_X65Y110_SLICE_X99Y110_C6 = CLBLM_R_X67Y109_SLICE_X100Y109_DO6;
  assign CLBLM_R_X65Y110_SLICE_X99Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X65Y110_SLICE_X99Y110_CX = CLBLM_R_X65Y110_SLICE_X98Y110_A5Q;
  assign CLBLM_R_X65Y110_SLICE_X99Y110_D1 = 1'b1;
  assign CLBLM_R_X65Y110_SLICE_X99Y110_D2 = CLBLM_L_X68Y108_SLICE_X102Y108_AQ;
  assign CLBLM_R_X65Y110_SLICE_X99Y110_D3 = 1'b1;
  assign CLBLM_R_X65Y110_SLICE_X99Y110_D4 = CLBLM_L_X68Y108_SLICE_X102Y108_A5Q;
  assign CLBLM_R_X65Y110_SLICE_X99Y110_D5 = CLBLM_R_X65Y110_SLICE_X98Y110_DQ;
  assign CLBLM_R_X65Y110_SLICE_X99Y110_D6 = CLBLM_R_X65Y110_SLICE_X99Y110_B5Q;
  assign CLBLM_R_X65Y110_SLICE_X99Y110_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X65Y110_SLICE_X98Y110_A1 = CLBLM_R_X67Y110_SLICE_X100Y110_BQ;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_A6 = CLBLM_L_X74Y128_SLICE_X113Y128_BO6;
  assign CLBLL_R_X71Y124_SLICE_X106Y124_A1 = CLBLM_L_X70Y125_SLICE_X105Y125_CO6;
  assign CLBLL_R_X71Y124_SLICE_X106Y124_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y124_SLICE_X106Y124_A3 = CLBLM_L_X70Y124_SLICE_X104Y124_BQ;
  assign CLBLL_R_X71Y124_SLICE_X106Y124_A4 = CLBLL_R_X73Y125_SLICE_X111Y125_A5Q;
  assign CLBLL_R_X71Y124_SLICE_X106Y124_A5 = CLBLL_R_X71Y125_SLICE_X106Y125_DO6;
  assign CLBLL_R_X71Y124_SLICE_X106Y124_A6 = 1'b1;
  assign CLBLM_R_X65Y110_SLICE_X98Y110_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y110_SLICE_X98Y110_A3 = CLBLM_R_X65Y110_SLICE_X98Y110_AQ;
  assign CLBLM_R_X65Y110_SLICE_X98Y110_A4 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLL_R_X71Y124_SLICE_X106Y124_B1 = CLBLL_R_X73Y125_SLICE_X110Y125_DO6;
  assign CLBLL_R_X71Y124_SLICE_X106Y124_B2 = CLBLL_R_X71Y124_SLICE_X106Y124_BQ;
  assign CLBLL_R_X71Y124_SLICE_X106Y124_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y124_SLICE_X106Y124_B4 = CLBLL_R_X71Y129_SLICE_X107Y129_BO6;
  assign CLBLL_R_X71Y124_SLICE_X106Y124_B5 = CLBLL_R_X71Y117_SLICE_X106Y117_BQ;
  assign CLBLL_R_X71Y124_SLICE_X106Y124_B6 = 1'b1;
  assign CLBLM_R_X65Y110_SLICE_X98Y110_B6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y110_SLICE_X98Y110_B1 = CLBLM_R_X65Y111_SLICE_X99Y111_AO5;
  assign CLBLL_R_X71Y124_SLICE_X106Y124_C1 = CLBLL_R_X71Y126_SLICE_X107Y126_AQ;
  assign CLBLL_R_X71Y124_SLICE_X106Y124_C2 = CLBLL_R_X71Y126_SLICE_X107Y126_BQ;
  assign CLBLL_R_X71Y124_SLICE_X106Y124_C3 = CLBLM_L_X70Y123_SLICE_X104Y123_AQ;
  assign CLBLL_R_X71Y124_SLICE_X106Y124_C4 = CLBLM_L_X70Y124_SLICE_X105Y124_BO6;
  assign CLBLL_R_X71Y124_SLICE_X106Y124_C5 = CLBLM_L_X70Y126_SLICE_X104Y126_CQ;
  assign CLBLL_R_X71Y124_SLICE_X106Y124_C6 = CLBLM_L_X70Y125_SLICE_X105Y125_AQ;
  assign CLBLM_R_X65Y110_SLICE_X98Y110_C1 = CLBLM_R_X65Y110_SLICE_X98Y110_BQ;
  assign CLBLM_R_X65Y110_SLICE_X98Y110_C2 = CLBLM_R_X65Y110_SLICE_X98Y110_CQ;
  assign CLBLL_R_X71Y124_SLICE_X106Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X65Y110_SLICE_X98Y110_C3 = CLBLM_R_X67Y111_SLICE_X101Y111_CO5;
  assign CLBLM_R_X65Y110_SLICE_X98Y110_C4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y110_SLICE_X98Y110_C5 = CLBLM_R_X65Y111_SLICE_X99Y111_AO5;
  assign CLBLM_R_X65Y110_SLICE_X98Y110_C6 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X65Y110_SLICE_X98Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X71Y124_SLICE_X106Y124_D1 = 1'b1;
  assign CLBLL_R_X71Y124_SLICE_X106Y124_D2 = 1'b1;
  assign CLBLL_R_X71Y124_SLICE_X106Y124_D3 = 1'b1;
  assign CLBLL_R_X71Y124_SLICE_X106Y124_D4 = 1'b1;
  assign CLBLL_R_X71Y124_SLICE_X106Y124_D5 = 1'b1;
  assign CLBLL_R_X71Y124_SLICE_X106Y124_D6 = 1'b1;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_C5 = CLBLL_R_X75Y113_SLICE_X114Y113_AQ;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_C6 = 1'b1;
  assign CLBLL_R_X71Y124_SLICE_X106Y124_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X65Y110_SLICE_X98Y110_D1 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X65Y110_SLICE_X98Y110_D2 = CLBLM_R_X65Y110_SLICE_X98Y110_CQ;
  assign CLBLM_R_X65Y110_SLICE_X98Y110_D3 = CLBLM_R_X65Y110_SLICE_X98Y110_DQ;
  assign CLBLM_R_X65Y110_SLICE_X98Y110_D4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y110_SLICE_X98Y110_D5 = CLBLM_R_X65Y111_SLICE_X99Y111_AO5;
  assign CLBLM_R_X65Y110_SLICE_X98Y110_D6 = CLBLM_R_X67Y111_SLICE_X101Y111_DO6;
  assign CLBLM_R_X65Y110_SLICE_X98Y110_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_D1 = CLBLM_L_X72Y123_SLICE_X108Y123_BO6;
  assign CLBLL_R_X71Y124_SLICE_X107Y124_A1 = 1'b1;
  assign CLBLL_R_X71Y124_SLICE_X107Y124_A2 = 1'b1;
  assign CLBLL_R_X71Y124_SLICE_X107Y124_A3 = 1'b1;
  assign CLBLL_R_X71Y124_SLICE_X107Y124_A4 = 1'b1;
  assign CLBLL_R_X71Y124_SLICE_X107Y124_A5 = 1'b1;
  assign CLBLL_R_X71Y124_SLICE_X107Y124_A6 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_T1 = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_D1 = CLBLM_L_X76Y128_SLICE_X116Y128_C5Q;
  assign CLBLL_R_X71Y124_SLICE_X107Y124_B1 = 1'b1;
  assign CLBLL_R_X71Y124_SLICE_X107Y124_B2 = 1'b1;
  assign CLBLL_R_X71Y124_SLICE_X107Y124_B3 = 1'b1;
  assign CLBLL_R_X71Y124_SLICE_X107Y124_B4 = 1'b1;
  assign CLBLL_R_X71Y124_SLICE_X107Y124_B5 = 1'b1;
  assign CLBLL_R_X71Y124_SLICE_X107Y124_B6 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_D1 = CLBLL_R_X71Y130_SLICE_X106Y130_DO6;
  assign CLBLL_R_X71Y124_SLICE_X107Y124_C1 = 1'b1;
  assign CLBLL_R_X71Y124_SLICE_X107Y124_C2 = 1'b1;
  assign CLBLL_R_X71Y124_SLICE_X107Y124_C3 = 1'b1;
  assign CLBLL_R_X71Y124_SLICE_X107Y124_C4 = 1'b1;
  assign CLBLL_R_X71Y124_SLICE_X107Y124_C5 = 1'b1;
  assign CLBLL_R_X71Y124_SLICE_X107Y124_C6 = 1'b1;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_D1 = CLBLM_L_X74Y123_SLICE_X113Y123_CO5;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_D2 = CLBLL_R_X75Y123_SLICE_X114Y123_BQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_T1 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_T1 = 1'b1;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_D3 = CLBLM_L_X74Y123_SLICE_X113Y123_DQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_D1 = 1'b0;
  assign CLBLL_R_X71Y124_SLICE_X107Y124_D1 = 1'b1;
  assign CLBLL_R_X71Y124_SLICE_X107Y124_D2 = 1'b1;
  assign CLBLL_R_X71Y124_SLICE_X107Y124_D3 = 1'b1;
  assign CLBLL_R_X71Y124_SLICE_X107Y124_D4 = 1'b1;
  assign CLBLL_R_X71Y124_SLICE_X107Y124_D5 = 1'b1;
  assign CLBLL_R_X71Y124_SLICE_X107Y124_D6 = 1'b1;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_D4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_D5 = 1'b1;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_A2 = CLBLM_L_X78Y123_SLICE_X121Y123_A5Q;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_D6 = CLBLL_R_X75Y121_SLICE_X114Y121_AO5;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_A3 = CLBLM_L_X78Y123_SLICE_X121Y123_AQ;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_A4 = CLBLM_L_X78Y123_SLICE_X120Y123_AO6;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_A5 = CLBLM_L_X78Y127_SLICE_X121Y127_DO6;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_A6 = 1'b1;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_B1 = CLBLM_L_X76Y122_SLICE_X117Y122_AQ;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_B2 = CLBLM_L_X78Y123_SLICE_X121Y123_BQ;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_B3 = CLBLL_R_X77Y113_SLICE_X118Y113_AQ;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_B4 = CLBLM_L_X72Y111_SLICE_X108Y111_C5Q;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_B6 = CLBLL_R_X77Y123_SLICE_X119Y123_BO5;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_C1 = CLBLL_R_X77Y113_SLICE_X118Y113_AQ;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_C2 = 1'b1;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_C3 = CLBLM_L_X72Y111_SLICE_X108Y111_C5Q;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_C4 = 1'b1;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_C5 = CLBLM_L_X76Y122_SLICE_X117Y122_AQ;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_C6 = 1'b1;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOI3_X105Y67_OLOGIC_X1Y67_D1 = CLBLM_R_X103Y67_SLICE_X163Y67_BQ;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_D1 = 1'b1;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_D2 = 1'b1;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_D3 = 1'b1;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_D4 = 1'b1;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_D5 = 1'b1;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_D6 = 1'b1;
  assign CLBLM_L_X70Y113_SLICE_X105Y113_A4 = 1'b1;
  assign RIOI3_X105Y67_OLOGIC_X1Y67_T1 = 1'b1;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_D1 = CLBLL_R_X79Y104_SLICE_X122Y104_A5Q;
  assign CLBLM_L_X70Y113_SLICE_X105Y113_A5 = 1'b1;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_A1 = CLBLM_L_X78Y124_SLICE_X120Y124_CQ;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_A1 = CLBLM_L_X74Y123_SLICE_X112Y123_DO6;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_A2 = CLBLL_R_X75Y123_SLICE_X114Y123_AO6;
  assign CLBLM_L_X70Y113_SLICE_X105Y113_A6 = 1'b1;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_A3 = CLBLL_R_X77Y124_SLICE_X118Y124_BQ;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_A4 = CLBLM_L_X78Y124_SLICE_X120Y124_AQ;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_A5 = CLBLM_L_X78Y124_SLICE_X120Y124_BQ;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_A6 = CLBLL_R_X77Y123_SLICE_X118Y123_AQ;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_A3 = CLBLM_L_X74Y123_SLICE_X112Y123_AQ;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_B1 = CLBLM_L_X78Y123_SLICE_X120Y123_DO6;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_B2 = CLBLL_R_X75Y123_SLICE_X114Y123_AO6;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_B3 = CLBLL_R_X77Y121_SLICE_X118Y121_AO6;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_B4 = CLBLM_L_X78Y123_SLICE_X121Y123_BQ;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_A4 = CLBLL_R_X73Y125_SLICE_X111Y125_AQ;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_B5 = CLBLL_R_X77Y113_SLICE_X118Y113_AQ;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_B6 = CLBLM_L_X72Y111_SLICE_X108Y111_C5Q;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_D1 = CLBLM_L_X76Y111_SLICE_X116Y111_AQ;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_A5 = CLBLM_L_X74Y123_SLICE_X113Y123_AQ;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_C1 = CLBLM_L_X78Y121_SLICE_X120Y121_CO5;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_C2 = CLBLM_L_X78Y123_SLICE_X121Y123_CO5;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_C3 = CLBLL_R_X75Y123_SLICE_X114Y123_AO6;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_C4 = CLBLL_R_X77Y121_SLICE_X118Y121_AO6;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_A6 = CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_C5 = CLBLM_L_X78Y123_SLICE_X120Y123_DO6;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_C6 = CLBLM_L_X78Y123_SLICE_X121Y123_BQ;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_T1 = 1'b1;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_D1 = CLBLM_L_X78Y124_SLICE_X120Y124_BQ;
  assign CLBLM_L_X70Y113_SLICE_X105Y113_B3 = 1'b1;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_D2 = CLBLM_L_X78Y124_SLICE_X120Y124_CQ;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_D3 = 1'b1;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_D4 = CLBLM_L_X78Y124_SLICE_X120Y124_AQ;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_D5 = CLBLL_R_X77Y124_SLICE_X118Y124_BQ;
  assign CLBLM_L_X70Y113_SLICE_X105Y113_B4 = 1'b1;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_B3 = CLBLM_L_X74Y128_SLICE_X113Y128_BO5;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_D6 = CLBLL_R_X77Y123_SLICE_X118Y123_AQ;
  assign CLBLM_L_X70Y113_SLICE_X105Y113_B5 = 1'b1;
  assign CLBLM_L_X70Y113_SLICE_X105Y113_B6 = 1'b1;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_B1 = CLBLM_L_X74Y123_SLICE_X112Y123_B5Q;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_B2 = CLBLM_L_X74Y123_SLICE_X112Y123_CO6;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_B3 = CLBLM_L_X74Y123_SLICE_X112Y123_AQ;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_B4 = 1'b1;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_B5 = CLBLM_L_X74Y123_SLICE_X113Y123_AQ;
  assign CLBLM_L_X70Y113_SLICE_X105Y113_C1 = 1'b1;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_B6 = 1'b1;
  assign CLBLM_L_X70Y113_SLICE_X105Y113_C2 = 1'b1;
  assign CLBLM_L_X70Y113_SLICE_X105Y113_C4 = 1'b1;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y113_SLICE_X105Y113_C5 = 1'b1;
  assign CLBLM_L_X70Y113_SLICE_X105Y113_C6 = 1'b1;
  assign CLBLM_R_X65Y111_SLICE_X99Y111_A1 = CLBLM_R_X67Y111_SLICE_X101Y111_A5Q;
  assign CLBLM_R_X65Y111_SLICE_X99Y111_A2 = 1'b1;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_C1 = CLBLM_L_X76Y125_SLICE_X117Y125_AQ;
  assign CLBLM_R_X65Y111_SLICE_X99Y111_A3 = 1'b1;
  assign CLBLM_R_X65Y111_SLICE_X99Y111_A4 = CLBLM_R_X67Y111_SLICE_X100Y111_A5Q;
  assign CLBLM_R_X65Y111_SLICE_X99Y111_A6 = 1'b1;
  assign CLBLM_R_X65Y111_SLICE_X99Y111_A5 = 1'b1;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_C2 = CLBLL_R_X75Y124_SLICE_X114Y124_BQ;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_B6 = CLBLM_L_X74Y128_SLICE_X113Y128_CQ;
  assign CLBLM_R_X65Y111_SLICE_X99Y111_B1 = 1'b1;
  assign CLBLM_R_X65Y111_SLICE_X99Y111_B2 = 1'b1;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_C3 = CLBLL_R_X75Y123_SLICE_X115Y123_DO6;
  assign CLBLM_R_X65Y111_SLICE_X99Y111_B3 = 1'b1;
  assign CLBLM_R_X65Y111_SLICE_X99Y111_B4 = 1'b1;
  assign CLBLM_R_X65Y111_SLICE_X99Y111_B5 = 1'b1;
  assign CLBLM_R_X65Y111_SLICE_X99Y111_B6 = 1'b1;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_C4 = CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  assign CLBLM_R_X65Y111_SLICE_X99Y111_C1 = 1'b1;
  assign CLBLM_R_X65Y111_SLICE_X99Y111_C2 = 1'b1;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_C5 = CLBLL_R_X75Y124_SLICE_X114Y124_AQ;
  assign CLBLM_R_X65Y111_SLICE_X99Y111_C3 = 1'b1;
  assign CLBLM_R_X65Y111_SLICE_X99Y111_C4 = 1'b1;
  assign CLBLM_R_X65Y111_SLICE_X99Y111_C5 = 1'b1;
  assign CLBLM_R_X65Y111_SLICE_X99Y111_C6 = 1'b1;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_C6 = CLBLL_R_X73Y125_SLICE_X111Y125_AQ;
  assign CLBLM_R_X65Y111_SLICE_X99Y111_D1 = 1'b1;
  assign CLBLM_R_X65Y111_SLICE_X99Y111_D2 = 1'b1;
  assign CLBLM_R_X65Y111_SLICE_X99Y111_D3 = 1'b1;
  assign CLBLM_R_X65Y111_SLICE_X99Y111_D4 = 1'b1;
  assign CLBLM_R_X65Y111_SLICE_X99Y111_D5 = 1'b1;
  assign CLBLM_R_X65Y111_SLICE_X99Y111_D6 = 1'b1;
  assign CLBLM_L_X70Y113_SLICE_X105Y113_D1 = 1'b1;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_A2 = CLBLL_R_X71Y125_SLICE_X106Y125_BQ;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_A3 = CLBLL_R_X71Y125_SLICE_X106Y125_AQ;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_A4 = 1'b1;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_A5 = CLBLL_R_X71Y125_SLICE_X107Y125_AQ;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_A6 = CLBLM_L_X70Y124_SLICE_X105Y124_CO6;
  assign CLBLM_L_X70Y113_SLICE_X105Y113_D2 = 1'b1;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X70Y113_SLICE_X105Y113_D3 = 1'b1;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_B1 = CLBLM_L_X70Y125_SLICE_X105Y125_AO5;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_B2 = CLBLL_R_X71Y125_SLICE_X106Y125_BQ;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_B3 = CLBLM_L_X70Y125_SLICE_X105Y125_BO6;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_B4 = CLBLM_L_X70Y126_SLICE_X104Y126_BQ;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_B6 = CLBLL_R_X71Y130_SLICE_X106Y130_CQ;
  assign CLBLM_L_X70Y113_SLICE_X105Y113_D4 = 1'b1;
  assign CLBLM_R_X65Y111_SLICE_X98Y111_A6 = CLBLM_R_X65Y110_SLICE_X99Y110_B5Q;
  assign CLBLM_L_X70Y113_SLICE_X105Y113_D5 = 1'b1;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_C1 = CLBLL_R_X71Y132_SLICE_X107Y132_BQ;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_C2 = CLBLL_R_X71Y125_SLICE_X106Y125_CQ;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_C3 = CLBLL_R_X71Y125_SLICE_X106Y125_BQ;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_C4 = CLBLM_L_X70Y125_SLICE_X105Y125_BO6;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_C5 = CLBLM_L_X70Y125_SLICE_X105Y125_AO5;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_C6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y113_SLICE_X105Y113_D6 = 1'b1;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X65Y111_SLICE_X98Y111_C1 = 1'b1;
  assign CLBLM_R_X65Y111_SLICE_X98Y111_C2 = 1'b1;
  assign CLBLM_R_X65Y111_SLICE_X98Y111_C3 = 1'b1;
  assign CLBLM_R_X65Y111_SLICE_X98Y111_C4 = 1'b1;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_D1 = CLBLM_L_X70Y124_SLICE_X104Y124_BQ;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_D2 = CLBLL_R_X71Y126_SLICE_X107Y126_AQ;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_D3 = CLBLL_R_X71Y125_SLICE_X107Y125_DO6;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_D4 = CLBLM_L_X70Y126_SLICE_X104Y126_CQ;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_D5 = CLBLL_R_X71Y126_SLICE_X106Y126_DO6;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_D6 = CLBLM_L_X70Y125_SLICE_X105Y125_AQ;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_D1 = CLBLM_L_X76Y125_SLICE_X117Y125_AQ;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_D2 = CLBLL_R_X75Y123_SLICE_X115Y123_DO6;
  assign CLBLM_L_X76Y130_SLICE_X117Y130_B2 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_A2 = CLBLM_R_X65Y104_SLICE_X99Y104_DO6;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_D3 = CLBLL_R_X75Y124_SLICE_X114Y124_AQ;
  assign CLBLM_L_X76Y130_SLICE_X117Y130_B3 = 1'b1;
  assign CLBLM_R_X65Y111_SLICE_X98Y111_D1 = 1'b1;
  assign CLBLM_R_X65Y111_SLICE_X98Y111_D2 = 1'b1;
  assign CLBLM_R_X65Y111_SLICE_X98Y111_D3 = 1'b1;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_D4 = CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  assign CLBLM_L_X76Y130_SLICE_X117Y130_B4 = 1'b1;
  assign CLBLM_R_X65Y111_SLICE_X98Y111_D6 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_A4 = CLBLM_R_X65Y104_SLICE_X98Y104_CQ;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_D5 = 1'b1;
  assign CLBLM_L_X76Y130_SLICE_X117Y130_B5 = 1'b1;
  assign CLBLM_R_X65Y111_SLICE_X98Y111_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign RIOI3_X105Y105_OLOGIC_X1Y105_T1 = 1'b1;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_D6 = CLBLL_R_X75Y124_SLICE_X114Y124_BQ;
  assign CLBLM_L_X76Y130_SLICE_X117Y130_B6 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X120Y128_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_A1 = CLBLL_R_X71Y125_SLICE_X107Y125_AQ;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_A2 = CLBLM_L_X70Y123_SLICE_X104Y123_AQ;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_A3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_A4 = CLBLL_R_X71Y126_SLICE_X107Y126_BQ;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_A5 = CLBLM_L_X70Y125_SLICE_X105Y125_BO5;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_A6 = CLBLL_R_X71Y125_SLICE_X106Y125_CQ;
  assign CLBLM_L_X78Y128_SLICE_X120Y128_A5 = CLBLL_R_X77Y128_SLICE_X118Y128_BQ;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_D1 = 1'b1;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_B1 = CLBLM_L_X70Y125_SLICE_X105Y125_AQ;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_B2 = CLBLM_L_X70Y123_SLICE_X104Y123_AQ;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_B3 = CLBLL_R_X71Y126_SLICE_X107Y126_AQ;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_B4 = CLBLM_L_X70Y124_SLICE_X105Y124_BO6;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_B5 = CLBLL_R_X71Y125_SLICE_X106Y125_AQ;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_B6 = CLBLL_R_X71Y126_SLICE_X107Y126_BQ;
  assign CLBLM_L_X70Y113_SLICE_X104Y113_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_C1 = CLBLM_L_X70Y124_SLICE_X105Y124_BO6;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_C2 = CLBLM_L_X70Y123_SLICE_X104Y123_AQ;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_C3 = CLBLM_L_X70Y125_SLICE_X105Y125_AQ;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_C4 = CLBLL_R_X71Y126_SLICE_X107Y126_AQ;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_C5 = CLBLL_R_X71Y125_SLICE_X107Y125_AQ;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_C6 = CLBLL_R_X71Y126_SLICE_X107Y126_BQ;
  assign CLBLM_L_X70Y113_SLICE_X104Y113_A6 = 1'b1;
  assign CLBLM_L_X76Y130_SLICE_X117Y130_C1 = 1'b1;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X76Y130_SLICE_X117Y130_C2 = 1'b1;
  assign CLBLM_L_X76Y130_SLICE_X117Y130_C3 = 1'b1;
  assign CLBLM_L_X76Y130_SLICE_X117Y130_C4 = 1'b1;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_D1 = CLBLM_L_X72Y123_SLICE_X108Y123_AQ;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_D2 = CLBLM_L_X72Y125_SLICE_X108Y125_AQ;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_D3 = CLBLL_R_X71Y126_SLICE_X107Y126_BO5;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_D4 = CLBLL_R_X71Y126_SLICE_X107Y126_AQ;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_D5 = CLBLM_L_X70Y124_SLICE_X105Y124_DO6;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_D6 = CLBLM_L_X70Y125_SLICE_X105Y125_AQ;
  assign CLBLM_L_X76Y130_SLICE_X117Y130_C5 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_A1 = 1'b1;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X76Y130_SLICE_X117Y130_C6 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_A2 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_A3 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_A4 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_A5 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_A6 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_B1 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_B2 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_B3 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_B4 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_B5 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_B6 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X120Y128_B3 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X120Y128_B4 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X120Y128_B5 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_C1 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_C2 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_C3 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_C4 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_C5 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_C6 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X120Y128_B6 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_T1 = 1'b1;
  assign CLBLM_L_X70Y113_SLICE_X104Y113_B6 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_D1 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_D2 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_D3 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_D4 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_D5 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_D6 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_A2 = CLBLL_R_X77Y124_SLICE_X118Y124_CO6;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_A3 = CLBLM_L_X78Y124_SLICE_X120Y124_AQ;
  assign CLBLM_L_X76Y130_SLICE_X117Y130_D1 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_A4 = CLBLM_L_X76Y124_SLICE_X117Y124_BQ;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_A5 = CLBLL_R_X77Y124_SLICE_X118Y124_BQ;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_A6 = CLBLL_R_X77Y123_SLICE_X119Y123_CQ;
  assign CLBLM_L_X76Y130_SLICE_X117Y130_D2 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_B1 = CLBLL_R_X77Y124_SLICE_X118Y124_CO6;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_B2 = CLBLM_L_X78Y124_SLICE_X120Y124_BQ;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_B3 = CLBLM_L_X78Y124_SLICE_X120Y124_AQ;
  assign CLBLM_L_X76Y130_SLICE_X117Y130_D3 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_B4 = CLBLL_R_X77Y123_SLICE_X119Y123_CQ;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_B6 = CLBLM_L_X76Y124_SLICE_X117Y124_BQ;
  assign CLBLM_L_X76Y130_SLICE_X117Y130_D4 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_C1 = CLBLL_R_X77Y123_SLICE_X119Y123_AQ;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_C2 = CLBLM_L_X78Y124_SLICE_X120Y124_CQ;
  assign CLBLM_L_X76Y130_SLICE_X117Y130_D5 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_C3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_C4 = CLBLL_R_X77Y123_SLICE_X119Y123_CQ;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_C5 = CLBLM_L_X76Y123_SLICE_X117Y123_AO5;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_C6 = CLBLM_L_X76Y124_SLICE_X117Y124_BQ;
  assign CLBLM_L_X76Y130_SLICE_X117Y130_D6 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X120Y128_C6 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X70Y113_SLICE_X104Y113_C5 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_D1 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_D2 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_D3 = 1'b1;
  assign CLBLM_L_X70Y113_SLICE_X104Y113_C6 = CLBLM_L_X72Y111_SLICE_X108Y111_BQ;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_D4 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_D5 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_D6 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X78Y128_SLICE_X120Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X70Y113_SLICE_X104Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X76Y130_SLICE_X116Y130_A1 = CLBLL_R_X75Y130_SLICE_X114Y130_AQ;
  assign CLBLM_L_X76Y130_SLICE_X116Y130_A2 = CLBLM_L_X76Y130_SLICE_X116Y130_BQ;
  assign CLBLM_L_X76Y130_SLICE_X116Y130_A3 = CLBLM_L_X76Y130_SLICE_X116Y130_AQ;
  assign CLBLM_L_X76Y130_SLICE_X116Y130_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X76Y130_SLICE_X116Y130_A5 = CLBLM_L_X76Y129_SLICE_X116Y129_BQ;
  assign CLBLM_L_X76Y130_SLICE_X116Y130_A6 = CLBLL_R_X75Y130_SLICE_X115Y130_BO5;
  assign CLBLM_L_X78Y128_SLICE_X120Y128_D4 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X120Y128_D5 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X120Y128_D6 = 1'b1;
  assign CLBLM_L_X70Y113_SLICE_X104Y113_D4 = 1'b1;
  assign CLBLM_L_X76Y130_SLICE_X116Y130_AX = CLBLM_L_X76Y130_SLICE_X116Y130_CO5;
  assign CLBLM_L_X70Y113_SLICE_X104Y113_D5 = 1'b1;
  assign CLBLM_L_X76Y130_SLICE_X116Y130_B1 = CLBLL_R_X75Y130_SLICE_X114Y130_AQ;
  assign CLBLM_L_X76Y130_SLICE_X116Y130_B2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X76Y130_SLICE_X116Y130_B3 = CLBLL_R_X77Y128_SLICE_X118Y128_CQ;
  assign CLBLM_L_X76Y130_SLICE_X116Y130_B4 = CLBLL_R_X77Y129_SLICE_X118Y129_CQ;
  assign CLBLM_L_X76Y130_SLICE_X116Y130_B5 = CLBLM_L_X76Y127_SLICE_X116Y127_AQ;
  assign CLBLM_L_X76Y130_SLICE_X116Y130_B6 = CLBLM_L_X76Y130_SLICE_X116Y130_BQ;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_A2 = CLBLL_R_X71Y126_SLICE_X106Y126_BQ;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_A3 = CLBLL_R_X71Y126_SLICE_X106Y126_AQ;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_A4 = CLBLL_R_X71Y126_SLICE_X107Y126_BQ;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_A5 = CLBLM_L_X70Y125_SLICE_X105Y125_BO5;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_A6 = CLBLM_L_X70Y123_SLICE_X104Y123_AQ;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_B1 = CLBLM_L_X72Y128_SLICE_X108Y128_AQ;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_B2 = CLBLL_R_X71Y126_SLICE_X106Y126_BQ;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_B3 = CLBLM_L_X70Y125_SLICE_X105Y125_BO6;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_B4 = CLBLM_L_X70Y125_SLICE_X105Y125_AO5;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_B5 = CLBLM_L_X70Y126_SLICE_X105Y126_BQ;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_B6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_D3 = 1'b1;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_C1 = CLBLM_L_X70Y124_SLICE_X105Y124_BO6;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_C2 = CLBLM_L_X70Y123_SLICE_X104Y123_AQ;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_C3 = CLBLM_L_X70Y125_SLICE_X105Y125_AQ;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_C4 = CLBLL_R_X71Y126_SLICE_X107Y126_AQ;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_C5 = CLBLL_R_X71Y126_SLICE_X107Y126_BQ;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_C6 = CLBLM_L_X70Y126_SLICE_X105Y126_AQ;
  assign CLBLL_R_X79Y127_SLICE_X122Y127_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X65Y111_SLICE_X98Y111_B1 = CLBLM_R_X65Y110_SLICE_X99Y110_AQ;
  assign CLBLM_L_X76Y130_SLICE_X116Y130_C1 = CLBLL_R_X75Y130_SLICE_X115Y130_BO5;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_D1 = CLBLL_R_X71Y126_SLICE_X107Y126_AQ;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_D2 = CLBLM_L_X70Y125_SLICE_X105Y125_AQ;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_D3 = CLBLL_R_X71Y126_SLICE_X106Y126_AQ;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_D4 = CLBLM_L_X70Y124_SLICE_X105Y124_DO6;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_D5 = 1'b1;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_D6 = CLBLM_L_X70Y126_SLICE_X105Y126_AQ;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_D4 = 1'b1;
  assign CLBLM_L_X76Y130_SLICE_X116Y130_C2 = CLBLL_R_X75Y130_SLICE_X114Y130_AQ;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X76Y130_SLICE_X116Y130_C3 = CLBLM_L_X76Y130_SLICE_X116Y130_BQ;
  assign CLBLM_L_X76Y130_SLICE_X116Y130_C4 = CLBLM_L_X76Y130_SLICE_X116Y130_A5Q;
  assign CLBLL_R_X79Y127_SLICE_X122Y127_A5 = CLBLL_R_X77Y125_SLICE_X118Y125_AQ;
  assign CLBLM_L_X76Y130_SLICE_X116Y130_C5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y111_SLICE_X98Y111_B2 = CLBLM_L_X76Y111_SLICE_X116Y111_AQ;
  assign CLBLM_L_X76Y130_SLICE_X116Y130_C6 = 1'b1;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_D5 = 1'b1;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_A1 = CLBLM_L_X70Y125_SLICE_X105Y125_AQ;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_A2 = CLBLM_L_X72Y129_SLICE_X108Y129_BQ;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_A3 = CLBLL_R_X71Y132_SLICE_X107Y132_CQ;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_A4 = CLBLL_R_X71Y126_SLICE_X107Y126_AQ;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_A6 = 1'b1;
  assign CLBLM_L_X76Y130_SLICE_X116Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_T1 = 1'b1;
  assign CLBLM_R_X65Y111_SLICE_X98Y111_B3 = CLBLM_R_X65Y111_SLICE_X98Y111_AQ;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_B1 = CLBLM_L_X72Y127_SLICE_X108Y127_CQ;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_B2 = CLBLL_R_X71Y127_SLICE_X107Y127_BQ;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_B3 = CLBLL_R_X71Y126_SLICE_X107Y126_AQ;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_B4 = CLBLM_L_X70Y125_SLICE_X105Y125_AQ;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_B6 = 1'b1;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_D6 = 1'b1;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_C1 = CLBLL_R_X73Y124_SLICE_X111Y124_BQ;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_C2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_C3 = CLBLL_R_X71Y127_SLICE_X107Y127_DQ;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_C4 = CLBLM_L_X72Y125_SLICE_X109Y125_AQ;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_C5 = CLBLM_L_X72Y128_SLICE_X108Y128_DQ;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_C6 = CLBLL_R_X71Y130_SLICE_X106Y130_DO5;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X65Y111_SLICE_X98Y111_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_D1 = CLBLL_R_X73Y124_SLICE_X111Y124_BQ;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_D2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_D3 = CLBLM_L_X72Y128_SLICE_X108Y128_DQ;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_D4 = CLBLM_L_X72Y125_SLICE_X109Y125_AQ;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_D5 = CLBLL_R_X71Y127_SLICE_X107Y127_DQ;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_D6 = 1'b1;
  assign CLBLM_L_X76Y130_SLICE_X116Y130_D1 = CLBLM_L_X76Y128_SLICE_X116Y128_C5Q;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X76Y130_SLICE_X116Y130_D2 = CLBLM_L_X76Y129_SLICE_X116Y129_CQ;
  assign CLBLM_L_X76Y130_SLICE_X116Y130_D3 = CLBLM_L_X76Y130_SLICE_X116Y130_DQ;
  assign CLBLM_L_X76Y130_SLICE_X116Y130_D4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y108_SLICE_X109Y108_D3 = CLBLM_L_X72Y108_SLICE_X109Y108_DQ;
  assign CLBLM_R_X65Y111_SLICE_X98Y111_B5 = CLBLM_L_X62Y92_SLICE_X92Y92_BQ;
  assign CLBLM_L_X76Y130_SLICE_X116Y130_D5 = CLBLM_L_X76Y129_SLICE_X116Y129_B5Q;
  assign CLBLM_L_X72Y108_SLICE_X109Y108_D4 = CLBLM_L_X72Y108_SLICE_X109Y108_CO6;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_D1 = CLBLM_L_X76Y125_SLICE_X116Y125_AQ;
  assign CLBLM_L_X76Y130_SLICE_X116Y130_D6 = CLBLM_L_X76Y129_SLICE_X116Y129_AQ;
  assign CLBLM_L_X72Y108_SLICE_X109Y108_D5 = CLBLM_L_X72Y109_SLICE_X108Y109_BO6;
  assign CLBLM_L_X72Y108_SLICE_X109Y108_D6 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X76Y111_SLICE_X116Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X79Y127_SLICE_X122Y127_AX = CLBLL_R_X83Y130_SLICE_X130Y130_DQ;
  assign CLBLM_R_X65Y111_SLICE_X98Y111_B6 = CLBLM_R_X65Y110_SLICE_X99Y110_B5Q;
  assign CLBLM_L_X76Y130_SLICE_X116Y130_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y108_SLICE_X109Y108_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_D1 = CLBLL_R_X73Y134_SLICE_X110Y134_AO5;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_T1 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_T1 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_D1 = CLBLM_L_X72Y118_SLICE_X109Y118_A5Q;
  assign CLBLM_R_X67Y110_SLICE_X101Y110_C3 = CLBLM_R_X67Y111_SLICE_X101Y111_DO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_D1 = CLBLL_R_X71Y124_SLICE_X106Y124_BO6;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_T1 = 1'b1;
  assign CLBLM_L_X70Y134_SLICE_X105Y134_D4 = 1'b1;
  assign CLBLM_L_X70Y134_SLICE_X105Y134_D5 = CLBLM_L_X72Y133_SLICE_X109Y133_CO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_T1 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_D1 = CLBLM_L_X68Y109_SLICE_X102Y109_AQ;
  assign CLBLM_L_X70Y134_SLICE_X105Y134_D6 = 1'b1;
  assign CLBLM_R_X67Y110_SLICE_X101Y110_C4 = CLBLM_R_X65Y110_SLICE_X99Y110_AO5;
  assign CLBLM_L_X76Y119_SLICE_X116Y119_C5 = 1'b1;
  assign RIOI3_X105Y71_OLOGIC_X1Y72_D1 = CLBLM_R_X103Y76_SLICE_X162Y76_AQ;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_T1 = 1'b1;
  assign RIOI3_X105Y71_OLOGIC_X1Y72_T1 = 1'b1;
  assign CLBLM_R_X67Y110_SLICE_X101Y110_C5 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X67Y115_SLICE_X101Y115_D4 = 1'b1;
  assign RIOI3_X105Y71_OLOGIC_X1Y71_D1 = CLBLM_R_X103Y75_SLICE_X162Y75_BQ;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_D1 = CLBLM_L_X70Y101_SLICE_X105Y101_AQ;
  assign RIOI3_X105Y71_OLOGIC_X1Y71_T1 = 1'b1;
  assign CLBLL_R_X79Y127_SLICE_X122Y127_B4 = CLBLL_R_X79Y127_SLICE_X122Y127_CQ;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_T1 = 1'b1;
  assign CLBLM_R_X67Y110_SLICE_X101Y110_C6 = CLBLM_R_X65Y110_SLICE_X99Y110_BQ;
  assign RIOB33_X105Y81_IOB_X1Y82_O = CLBLL_R_X77Y104_SLICE_X119Y104_A5Q;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_D1 = CLBLM_L_X62Y106_SLICE_X92Y106_BQ;
  assign CLBLM_L_X78Y104_SLICE_X120Y104_B2 = 1'b1;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_D6 = CLBLM_L_X72Y124_SLICE_X108Y124_BO6;
  assign CLBLL_R_X79Y127_SLICE_X122Y127_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_T1 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_A1 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_A2 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_A3 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_A4 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_A5 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_A6 = 1'b1;
  assign CLBLM_L_X72Y108_SLICE_X108Y108_C5 = CLBLL_R_X71Y109_SLICE_X106Y109_CO6;
  assign CLBLM_L_X72Y108_SLICE_X108Y108_C6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_B1 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_B2 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_B3 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_B4 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_B5 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_B6 = 1'b1;
  assign CLBLL_R_X79Y127_SLICE_X122Y127_B6 = 1'b1;
  assign CLBLM_L_X78Y104_SLICE_X120Y104_B3 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_C1 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_C2 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_C3 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_C4 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_C5 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_C6 = 1'b1;
  assign CLBLM_L_X70Y134_SLICE_X104Y134_B3 = CLBLM_L_X72Y134_SLICE_X109Y134_AO6;
  assign CLBLM_L_X72Y108_SLICE_X108Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A1 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A4 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A5 = CLBLL_R_X73Y123_SLICE_X110Y123_AQ;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_D1 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_D2 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_D3 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_D4 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_D5 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_D6 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A6 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B1 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B4 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B5 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B6 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C1 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C4 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C5 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C6 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_AX = CLBLM_L_X74Y126_SLICE_X113Y126_AQ;
  assign CLBLM_L_X78Y130_SLICE_X121Y130_B1 = 1'b1;
  assign CLBLM_L_X78Y104_SLICE_X120Y104_B5 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D1 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D4 = 1'b1;
  assign CLBLM_L_X68Y98_SLICE_X103Y98_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D5 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D6 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_A2 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_A5 = CLBLM_L_X72Y126_SLICE_X109Y126_AQ;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_A6 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_A3 = CLBLL_R_X71Y127_SLICE_X107Y127_AQ;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_A4 = CLBLL_R_X71Y126_SLICE_X106Y126_CO6;
  assign CLBLM_L_X70Y134_SLICE_X104Y134_C2 = CLBLM_L_X70Y133_SLICE_X104Y133_A5Q;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_B1 = CLBLL_R_X73Y126_SLICE_X110Y126_A5Q;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_B2 = CLBLL_R_X71Y127_SLICE_X107Y127_BQ;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_B3 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_B4 = CLBLM_L_X72Y127_SLICE_X109Y127_AO6;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_B5 = CLBLL_R_X71Y126_SLICE_X106Y126_CO6;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_B6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y134_SLICE_X104Y134_C3 = CLBLM_L_X70Y133_SLICE_X105Y133_AQ;
  assign CLBLM_L_X70Y134_SLICE_X104Y134_C5 = CLBLM_L_X70Y135_SLICE_X104Y135_BQ;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_C1 = CLBLL_R_X71Y127_SLICE_X107Y127_BQ;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_C2 = CLBLL_R_X71Y127_SLICE_X107Y127_CQ;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_C3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_C4 = CLBLM_L_X72Y126_SLICE_X109Y126_AQ;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_C5 = CLBLL_R_X71Y127_SLICE_X107Y127_AQ;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_C6 = CLBLL_R_X71Y126_SLICE_X106Y126_CO6;
  assign CLBLM_L_X70Y134_SLICE_X104Y134_C6 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X65Y111_SLICE_X98Y111_C5 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A1 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A4 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_D1 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_D2 = CLBLL_R_X71Y127_SLICE_X107Y127_CQ;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_D3 = CLBLL_R_X75Y127_SLICE_X114Y127_DQ;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_D4 = CLBLL_R_X71Y127_SLICE_X107Y127_AO5;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A5 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_D6 = CLBLL_R_X71Y127_SLICE_X107Y127_DQ;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_D5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A6 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B1 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B4 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B5 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B6 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C1 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C4 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C5 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C6 = 1'b1;
  assign CLBLM_L_X74Y103_SLICE_X113Y103_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y111_SLICE_X98Y111_C6 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D1 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D4 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D5 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D6 = 1'b1;
  assign CLBLM_L_X68Y98_SLICE_X102Y98_B1 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X74Y103_SLICE_X113Y103_C1 = CLBLM_L_X74Y102_SLICE_X112Y102_AQ;
  assign CLBLM_L_X70Y134_SLICE_X104Y134_D3 = CLBLM_L_X70Y134_SLICE_X104Y134_BQ;
  assign CLBLM_L_X74Y103_SLICE_X113Y103_C2 = CLBLM_L_X72Y104_SLICE_X109Y104_B5Q;
  assign CLBLM_L_X70Y134_SLICE_X104Y134_D4 = CLBLM_L_X70Y135_SLICE_X104Y135_AQ;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_A6 = 1'b1;
  assign CLBLM_L_X70Y134_SLICE_X104Y134_D5 = 1'b1;
  assign CLBLM_L_X70Y134_SLICE_X104Y134_D6 = CLBLM_L_X70Y133_SLICE_X104Y133_AQ;
  assign CLBLM_L_X74Y103_SLICE_X113Y103_C5 = CLBLL_R_X75Y103_SLICE_X115Y103_AQ;
  assign CLBLM_L_X78Y130_SLICE_X121Y130_B2 = 1'b1;
  assign CLBLM_L_X68Y98_SLICE_X102Y98_C3 = CLBLM_L_X68Y98_SLICE_X102Y98_BQ;
  assign CLBLM_L_X68Y98_SLICE_X102Y98_C4 = CLBLM_R_X67Y98_SLICE_X101Y98_BO6;
  assign CLBLM_R_X67Y110_SLICE_X101Y110_D1 = CLBLM_R_X67Y111_SLICE_X100Y111_CO5;
  assign CLBLM_L_X68Y98_SLICE_X102Y98_C6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X78Y104_SLICE_X120Y104_C1 = 1'b1;
  assign CLBLM_L_X74Y103_SLICE_X113Y103_D3 = CLBLL_R_X73Y103_SLICE_X111Y103_A5Q;
  assign CLBLM_L_X68Y98_SLICE_X102Y98_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X67Y110_SLICE_X101Y110_D2 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X74Y103_SLICE_X113Y103_D5 = CLBLL_R_X73Y101_SLICE_X110Y101_AQ;
  assign CLBLM_L_X74Y103_SLICE_X113Y103_D6 = CLBLM_L_X72Y104_SLICE_X109Y104_BQ;
  assign CLBLM_R_X67Y110_SLICE_X101Y110_D3 = CLBLM_R_X67Y110_SLICE_X101Y110_DQ;
  assign CLBLM_L_X74Y103_SLICE_X113Y103_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign RIOB33_X105Y103_IOB_X1Y104_O = CLBLM_L_X72Y106_SLICE_X108Y106_AQ;
  assign RIOB33_X105Y103_IOB_X1Y103_O = CLBLL_R_X77Y128_SLICE_X119Y128_DQ;
  assign CLBLM_R_X67Y110_SLICE_X101Y110_D4 = CLBLM_R_X67Y110_SLICE_X100Y110_CQ;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_A1 = CLBLM_L_X70Y129_SLICE_X105Y129_DQ;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_A3 = CLBLL_R_X71Y128_SLICE_X106Y128_AQ;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_A4 = CLBLM_L_X70Y126_SLICE_X105Y126_CO6;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_A5 = CLBLM_L_X70Y128_SLICE_X104Y128_BQ;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_A6 = CLBLM_L_X70Y129_SLICE_X104Y129_AQ;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_B1 = CLBLM_L_X70Y129_SLICE_X105Y129_DQ;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_B2 = CLBLL_R_X71Y128_SLICE_X106Y128_BQ;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_B3 = CLBLL_R_X71Y128_SLICE_X106Y128_AQ;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_B4 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_B6 = CLBLL_R_X71Y128_SLICE_X106Y128_CO6;
  assign CLBLM_R_X67Y110_SLICE_X101Y110_D5 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_C1 = CLBLM_L_X70Y128_SLICE_X104Y128_BQ;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_C2 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_C3 = CLBLM_L_X70Y129_SLICE_X104Y129_AQ;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_C4 = CLBLM_L_X70Y126_SLICE_X105Y126_CO6;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_C5 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_C6 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_D1 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_D2 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_D3 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_D4 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_D5 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_D6 = 1'b1;
  assign CLBLM_R_X67Y110_SLICE_X101Y110_D6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y103_SLICE_X112Y103_B2 = CLBLM_L_X74Y103_SLICE_X112Y103_BQ;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y103_SLICE_X112Y103_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y103_SLICE_X112Y103_B4 = CLBLL_R_X73Y103_SLICE_X111Y103_AQ;
  assign CLBLM_L_X74Y103_SLICE_X112Y103_B6 = CLBLM_L_X72Y103_SLICE_X108Y103_A5Q;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_D1 = CLBLM_R_X67Y118_SLICE_X101Y118_AQ;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_A1 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_A2 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_A3 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_A4 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_A5 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_A6 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_B1 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_B2 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_B3 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_B4 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_B5 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_B6 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_A2 = CLBLM_L_X72Y129_SLICE_X108Y129_AQ;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_A3 = CLBLL_R_X71Y125_SLICE_X107Y125_BO6;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_C1 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_C2 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_C3 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_C4 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_C5 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_C6 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_A4 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_A5 = CLBLL_R_X71Y130_SLICE_X106Y130_BQ;
  assign CLBLM_L_X74Y103_SLICE_X112Y103_C1 = CLBLM_L_X72Y104_SLICE_X109Y104_BQ;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_A6 = 1'b1;
  assign CLBLM_L_X74Y103_SLICE_X112Y103_C2 = CLBLL_R_X73Y103_SLICE_X110Y103_A5Q;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_D1 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_D2 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_D3 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_D4 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_D5 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_D6 = 1'b1;
  assign CLBLM_L_X74Y103_SLICE_X112Y103_C3 = CLBLM_L_X74Y103_SLICE_X112Y103_AQ;
  assign CLBLM_L_X74Y103_SLICE_X112Y103_C4 = CLBLL_R_X73Y102_SLICE_X110Y102_A5Q;
  assign CLBLM_L_X74Y103_SLICE_X112Y103_C5 = CLBLM_L_X74Y103_SLICE_X112Y103_BQ;
  assign CLBLM_L_X74Y103_SLICE_X112Y103_C6 = CLBLM_L_X72Y104_SLICE_X109Y104_B5Q;
  assign CLBLM_L_X78Y127_SLICE_X121Y127_A1 = CLBLL_R_X79Y128_SLICE_X122Y128_CQ;
  assign CLBLM_L_X78Y127_SLICE_X121Y127_A2 = CLBLL_R_X79Y128_SLICE_X122Y128_BQ;
  assign CLBLM_L_X78Y127_SLICE_X121Y127_A3 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_B1 = CLBLL_R_X71Y130_SLICE_X107Y130_AO6;
  assign CLBLM_L_X78Y127_SLICE_X121Y127_A4 = CLBLL_R_X79Y128_SLICE_X122Y128_AQ;
  assign CLBLM_L_X78Y127_SLICE_X121Y127_A5 = CLBLL_R_X79Y127_SLICE_X122Y127_BQ;
  assign CLBLM_L_X78Y127_SLICE_X121Y127_A6 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_B2 = CLBLM_L_X72Y129_SLICE_X108Y129_BQ;
  assign CLBLM_L_X78Y127_SLICE_X121Y127_B1 = 1'b1;
  assign CLBLM_L_X78Y127_SLICE_X121Y127_B2 = CLBLL_R_X79Y127_SLICE_X122Y127_CQ;
  assign CLBLM_L_X78Y127_SLICE_X121Y127_B3 = CLBLL_R_X79Y128_SLICE_X122Y128_DQ;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X78Y127_SLICE_X121Y127_B4 = CLBLL_R_X77Y127_SLICE_X119Y127_AQ;
  assign CLBLM_L_X78Y127_SLICE_X121Y127_B5 = CLBLL_R_X79Y127_SLICE_X122Y127_AQ;
  assign CLBLM_L_X74Y103_SLICE_X112Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X78Y127_SLICE_X121Y127_B6 = CLBLM_L_X78Y127_SLICE_X121Y127_AO5;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_B4 = 1'b1;
  assign CLBLM_L_X78Y127_SLICE_X121Y127_C1 = CLBLM_L_X78Y127_SLICE_X121Y127_AO6;
  assign CLBLM_L_X78Y127_SLICE_X121Y127_C2 = CLBLL_R_X79Y127_SLICE_X122Y127_CQ;
  assign CLBLM_L_X78Y127_SLICE_X121Y127_C3 = CLBLL_R_X79Y128_SLICE_X122Y128_DQ;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_B5 = CLBLL_R_X71Y125_SLICE_X107Y125_BO6;
  assign CLBLM_L_X78Y127_SLICE_X121Y127_C4 = 1'b1;
  assign CLBLM_L_X78Y127_SLICE_X121Y127_C5 = 1'b1;
  assign CLBLM_L_X78Y127_SLICE_X121Y127_C6 = CLBLL_R_X79Y127_SLICE_X122Y127_AQ;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_B6 = CLBLL_R_X71Y129_SLICE_X106Y129_AQ;
  assign CLBLM_L_X78Y127_SLICE_X121Y127_D1 = CLBLL_R_X79Y127_SLICE_X122Y127_AQ;
  assign CLBLM_L_X78Y127_SLICE_X121Y127_D2 = CLBLL_R_X79Y127_SLICE_X122Y127_BQ;
  assign CLBLM_L_X78Y127_SLICE_X121Y127_D3 = 1'b1;
  assign CLBLM_L_X78Y127_SLICE_X121Y127_D4 = CLBLL_R_X79Y127_SLICE_X122Y127_DO6;
  assign CLBLM_L_X78Y127_SLICE_X121Y127_D5 = 1'b1;
  assign CLBLM_L_X78Y127_SLICE_X121Y127_D6 = CLBLL_R_X79Y128_SLICE_X122Y128_BQ;
  assign CLBLM_R_X103Y75_SLICE_X163Y75_A1 = 1'b1;
  assign CLBLM_R_X103Y75_SLICE_X163Y75_A2 = 1'b1;
  assign CLBLM_R_X103Y75_SLICE_X163Y75_A3 = 1'b1;
  assign CLBLM_R_X103Y75_SLICE_X163Y75_A4 = 1'b1;
  assign CLBLM_R_X103Y75_SLICE_X163Y75_A5 = 1'b1;
  assign CLBLM_L_X72Y103_SLICE_X109Y103_A1 = CLBLM_L_X72Y104_SLICE_X109Y104_B5Q;
  assign CLBLM_L_X72Y103_SLICE_X109Y103_A2 = CLBLL_R_X73Y104_SLICE_X110Y104_A5Q;
  assign CLBLM_L_X72Y103_SLICE_X109Y103_A3 = CLBLM_L_X60Y101_SLICE_X90Y101_AQ;
  assign CLBLM_L_X72Y103_SLICE_X109Y103_A4 = CLBLM_L_X72Y104_SLICE_X109Y104_BQ;
  assign CLBLM_L_X72Y103_SLICE_X109Y103_A5 = CLBLM_L_X70Y105_SLICE_X104Y105_BO6;
  assign CLBLM_L_X72Y103_SLICE_X109Y103_A6 = 1'b1;
  assign CLBLM_L_X74Y103_SLICE_X112Y103_D1 = CLBLM_L_X74Y103_SLICE_X113Y103_AQ;
  assign CLBLM_L_X72Y103_SLICE_X109Y103_AX = CLBLL_R_X73Y103_SLICE_X110Y103_A5Q;
  assign CLBLM_L_X74Y103_SLICE_X112Y103_D2 = CLBLM_L_X72Y103_SLICE_X109Y103_AQ;
  assign CLBLM_L_X72Y103_SLICE_X109Y103_B1 = CLBLL_R_X73Y104_SLICE_X110Y104_CQ;
  assign CLBLM_L_X72Y103_SLICE_X109Y103_B2 = CLBLM_L_X72Y103_SLICE_X109Y103_BQ;
  assign CLBLM_L_X72Y103_SLICE_X109Y103_B3 = CLBLM_L_X72Y103_SLICE_X108Y103_CO5;
  assign CLBLM_L_X72Y103_SLICE_X109Y103_B4 = CLBLM_L_X72Y103_SLICE_X108Y103_BO5;
  assign CLBLM_L_X72Y103_SLICE_X109Y103_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y103_SLICE_X109Y103_B6 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_C1 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_C2 = 1'b1;
  assign CLBLM_L_X74Y103_SLICE_X112Y103_D3 = CLBLL_R_X75Y103_SLICE_X115Y103_AQ;
  assign CLBLM_L_X72Y103_SLICE_X109Y103_C1 = CLBLM_L_X70Y105_SLICE_X104Y105_BO6;
  assign CLBLM_L_X72Y103_SLICE_X109Y103_C2 = CLBLL_R_X73Y104_SLICE_X110Y104_A5Q;
  assign CLBLM_L_X72Y103_SLICE_X109Y103_C3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y103_SLICE_X109Y103_C4 = CLBLM_L_X60Y101_SLICE_X90Y101_AQ;
  assign CLBLM_L_X72Y103_SLICE_X109Y103_C5 = CLBLM_L_X72Y104_SLICE_X109Y104_B5Q;
  assign CLBLM_L_X72Y103_SLICE_X109Y103_C6 = CLBLM_L_X72Y104_SLICE_X109Y104_BQ;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_C3 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_C4 = 1'b1;
  assign CLBLM_L_X72Y103_SLICE_X109Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y103_SLICE_X112Y103_D5 = CLBLM_L_X72Y104_SLICE_X109Y104_B5Q;
  assign CLBLM_L_X74Y103_SLICE_X112Y103_D6 = CLBLM_L_X74Y104_SLICE_X112Y104_AQ;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_C5 = 1'b1;
  assign CLBLM_L_X78Y127_SLICE_X120Y127_C2 = 1'b1;
  assign CLBLM_L_X78Y127_SLICE_X120Y127_C4 = 1'b1;
  assign CLBLM_L_X72Y103_SLICE_X109Y103_D1 = CLBLM_L_X72Y103_SLICE_X109Y103_BQ;
  assign CLBLM_L_X72Y103_SLICE_X109Y103_D2 = CLBLL_R_X73Y104_SLICE_X110Y104_CQ;
  assign CLBLM_L_X72Y103_SLICE_X109Y103_D3 = CLBLM_L_X72Y104_SLICE_X109Y104_B5Q;
  assign CLBLM_L_X72Y103_SLICE_X109Y103_D4 = CLBLL_R_X73Y103_SLICE_X110Y103_A5Q;
  assign CLBLM_L_X72Y103_SLICE_X109Y103_D5 = CLBLM_L_X72Y103_SLICE_X109Y103_AQ;
  assign CLBLM_L_X72Y103_SLICE_X109Y103_D6 = CLBLM_L_X72Y104_SLICE_X109Y104_BQ;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_C6 = 1'b1;
  assign CLBLM_L_X72Y103_SLICE_X109Y103_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X78Y127_SLICE_X120Y127_D1 = 1'b1;
  assign CLBLM_L_X78Y127_SLICE_X120Y127_D2 = 1'b1;
  assign CLBLM_L_X78Y127_SLICE_X120Y127_D3 = 1'b1;
  assign CLBLM_L_X72Y103_SLICE_X108Y103_A1 = 1'b1;
  assign CLBLM_L_X72Y103_SLICE_X108Y103_A2 = CLBLM_L_X72Y103_SLICE_X108Y103_A5Q;
  assign CLBLM_L_X72Y103_SLICE_X108Y103_A3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y103_SLICE_X108Y103_A4 = CLBLM_L_X72Y103_SLICE_X108Y103_AQ;
  assign CLBLM_L_X72Y103_SLICE_X108Y103_A5 = CLBLM_L_X72Y104_SLICE_X109Y104_AQ;
  assign CLBLM_L_X72Y103_SLICE_X108Y103_A6 = 1'b1;
  assign CLBLM_L_X74Y103_SLICE_X112Y103_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X103Y75_SLICE_X162Y75_B1 = 1'b1;
  assign CLBLM_L_X72Y103_SLICE_X108Y103_B1 = 1'b1;
  assign CLBLM_L_X72Y103_SLICE_X108Y103_B2 = CLBLM_L_X72Y103_SLICE_X108Y103_A5Q;
  assign CLBLM_L_X72Y103_SLICE_X108Y103_B3 = 1'b1;
  assign CLBLM_L_X72Y103_SLICE_X108Y103_B4 = CLBLM_L_X72Y103_SLICE_X108Y103_AQ;
  assign CLBLM_L_X72Y103_SLICE_X108Y103_B5 = CLBLM_L_X72Y104_SLICE_X109Y104_AQ;
  assign CLBLM_L_X72Y103_SLICE_X108Y103_B6 = 1'b1;
  assign CLBLM_R_X103Y75_SLICE_X162Y75_BX = CLBLM_R_X103Y75_SLICE_X162Y75_AQ;
  assign CLBLM_R_X103Y75_SLICE_X162Y75_C1 = 1'b1;
  assign CLBLM_R_X103Y75_SLICE_X162Y75_C2 = 1'b1;
  assign CLBLM_R_X103Y75_SLICE_X162Y75_C3 = 1'b1;
  assign CLBLM_L_X72Y103_SLICE_X108Y103_C1 = 1'b1;
  assign CLBLM_L_X72Y103_SLICE_X108Y103_C2 = CLBLM_L_X72Y104_SLICE_X109Y104_A5Q;
  assign CLBLM_L_X72Y103_SLICE_X108Y103_C3 = CLBLL_R_X73Y104_SLICE_X110Y104_BQ;
  assign CLBLM_L_X72Y103_SLICE_X108Y103_C4 = 1'b1;
  assign CLBLM_L_X72Y103_SLICE_X108Y103_C5 = 1'b1;
  assign CLBLM_L_X72Y103_SLICE_X108Y103_C6 = 1'b1;
  assign CLBLM_R_X103Y75_SLICE_X162Y75_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X103Y75_SLICE_X162Y75_CX = CLBLM_R_X103Y75_SLICE_X162Y75_BQ;
  assign CLBLM_R_X103Y75_SLICE_X162Y75_D1 = 1'b1;
  assign CLBLM_L_X72Y103_SLICE_X108Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X103Y75_SLICE_X162Y75_D2 = 1'b1;
  assign CLBLM_R_X103Y75_SLICE_X162Y75_D3 = 1'b1;
  assign CLBLM_R_X103Y75_SLICE_X162Y75_D4 = 1'b1;
  assign CLBLM_R_X103Y75_SLICE_X162Y75_D5 = 1'b1;
  assign CLBLM_L_X72Y103_SLICE_X108Y103_D1 = CLBLM_L_X72Y104_SLICE_X109Y104_AQ;
  assign CLBLM_L_X72Y103_SLICE_X108Y103_D2 = CLBLM_L_X72Y103_SLICE_X108Y103_AQ;
  assign CLBLM_L_X72Y103_SLICE_X108Y103_D3 = 1'b1;
  assign CLBLM_L_X72Y103_SLICE_X108Y103_D4 = 1'b1;
  assign CLBLM_L_X72Y103_SLICE_X108Y103_D5 = 1'b1;
  assign CLBLM_L_X72Y103_SLICE_X108Y103_D6 = 1'b1;
  assign CLBLM_R_X103Y75_SLICE_X162Y75_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign RIOB33_X105Y105_IOB_X1Y105_O = CLBLM_R_X65Y111_SLICE_X98Y111_AQ;
  assign CLBLM_L_X72Y103_SLICE_X108Y103_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_D2 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_D3 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_D4 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_D5 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_D6 = 1'b1;
  assign RIOI3_X105Y83_OLOGIC_X1Y83_T1 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_A1 = CLBLM_L_X72Y129_SLICE_X108Y129_AQ;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_A2 = CLBLL_R_X71Y125_SLICE_X107Y125_BO6;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_A3 = CLBLL_R_X71Y129_SLICE_X106Y129_AQ;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_A4 = CLBLL_R_X71Y129_SLICE_X107Y129_BQ;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_A6 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_D1 = CLBLM_L_X64Y105_SLICE_X97Y105_DO6;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_B1 = CLBLM_L_X72Y130_SLICE_X109Y130_CQ;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_B2 = CLBLL_R_X71Y130_SLICE_X106Y130_BQ;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_B3 = CLBLL_R_X71Y129_SLICE_X106Y129_AQ;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_B5 = CLBLL_R_X71Y125_SLICE_X107Y125_BO6;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_B6 = CLBLL_R_X71Y129_SLICE_X106Y129_BQ;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_T1 = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_D1 = 1'b0;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_C2 = CLBLL_R_X71Y129_SLICE_X106Y129_CQ;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_C3 = CLBLL_R_X71Y129_SLICE_X106Y129_BQ;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_C4 = CLBLM_L_X72Y130_SLICE_X109Y130_CQ;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_C5 = CLBLL_R_X71Y129_SLICE_X106Y129_DO6;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_C6 = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_D1 = CLBLM_L_X72Y128_SLICE_X109Y128_AO6;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_T1 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_D1 = CLBLL_R_X71Y125_SLICE_X107Y125_BO6;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_D2 = CLBLL_R_X71Y129_SLICE_X106Y129_AQ;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_D3 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_D4 = CLBLL_R_X71Y130_SLICE_X106Y130_BQ;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_D5 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_D6 = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_T1 = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_D1 = CLBLL_R_X73Y104_SLICE_X110Y104_AQ;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign RIOI3_X105Y73_OLOGIC_X1Y74_D1 = CLBLM_R_X103Y75_SLICE_X162Y75_AQ;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_T1 = 1'b1;
  assign CLBLM_R_X67Y110_SLICE_X100Y110_A6 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign RIOI3_X105Y73_OLOGIC_X1Y74_T1 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_A1 = CLBLL_R_X71Y130_SLICE_X107Y130_DO6;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_A2 = CLBLM_L_X72Y130_SLICE_X109Y130_BQ;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_A3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_A4 = CLBLL_R_X71Y128_SLICE_X106Y128_BQ;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_A5 = CLBLL_R_X71Y133_SLICE_X106Y133_DQ;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_A6 = CLBLL_R_X71Y129_SLICE_X106Y129_CQ;
  assign RIOI3_X105Y73_OLOGIC_X1Y73_D1 = CLBLM_R_X103Y75_SLICE_X163Y75_AQ;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_AX = CLBLM_L_X70Y130_SLICE_X105Y130_AQ;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_B1 = CLBLM_L_X72Y132_SLICE_X109Y132_AQ;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_B2 = CLBLM_L_X70Y132_SLICE_X105Y132_BQ;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_B3 = CLBLL_R_X71Y129_SLICE_X107Y129_AQ;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_B4 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_B5 = CLBLL_R_X71Y130_SLICE_X107Y130_AQ;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_B6 = CLBLL_R_X71Y129_SLICE_X107Y129_CO6;
  assign RIOI3_X105Y73_OLOGIC_X1Y73_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_BX = CLBLM_L_X72Y129_SLICE_X108Y129_AQ;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_C1 = CLBLL_R_X71Y130_SLICE_X107Y130_BQ;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_C2 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_C3 = CLBLL_R_X71Y129_SLICE_X107Y129_BQ;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_C4 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_C5 = CLBLM_L_X70Y128_SLICE_X105Y128_AQ;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_C6 = CLBLM_L_X70Y132_SLICE_X105Y132_AQ;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_CE = CLBLM_L_X76Y109_SLICE_X116Y109_AO6;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_D1 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_D2 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_D3 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_D4 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_D5 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X121Y128_A1 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X121Y128_A2 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X121Y128_A3 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X121Y128_A4 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X121Y128_A5 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X121Y128_A6 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X121Y128_B1 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X121Y128_B2 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X121Y128_B3 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X121Y128_B4 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X121Y128_B5 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X121Y128_B6 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X121Y128_C1 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X121Y128_C2 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X121Y128_C3 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X121Y128_C4 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X121Y128_C5 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X121Y128_C6 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X121Y128_D1 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X121Y128_D2 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X121Y128_D3 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X121Y128_D4 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X121Y128_D5 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X121Y128_D6 = 1'b1;
  assign CLBLM_R_X103Y76_SLICE_X163Y76_A1 = 1'b1;
  assign CLBLM_R_X103Y76_SLICE_X163Y76_A2 = 1'b1;
  assign CLBLM_R_X103Y76_SLICE_X163Y76_A3 = 1'b1;
  assign CLBLM_R_X103Y76_SLICE_X163Y76_A4 = 1'b1;
  assign CLBLM_R_X103Y76_SLICE_X163Y76_A5 = 1'b1;
  assign CLBLM_R_X103Y76_SLICE_X163Y76_A6 = 1'b1;
  assign CLBLM_L_X72Y104_SLICE_X109Y104_A1 = CLBLM_L_X72Y103_SLICE_X108Y103_A5Q;
  assign CLBLM_L_X72Y104_SLICE_X109Y104_A2 = CLBLM_L_X72Y104_SLICE_X109Y104_A5Q;
  assign CLBLM_L_X72Y104_SLICE_X109Y104_A3 = CLBLM_L_X72Y104_SLICE_X109Y104_AQ;
  assign CLBLM_L_X72Y104_SLICE_X109Y104_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y104_SLICE_X109Y104_A5 = 1'b1;
  assign CLBLM_L_X72Y104_SLICE_X109Y104_A6 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X120Y128_A1 = CLBLL_R_X77Y128_SLICE_X119Y128_BQ;
  assign CLBLM_L_X78Y128_SLICE_X120Y128_A2 = CLBLL_R_X77Y128_SLICE_X118Y128_CQ;
  assign CLBLM_L_X78Y128_SLICE_X120Y128_A3 = CLBLM_L_X78Y128_SLICE_X120Y128_AQ;
  assign CLBLM_L_X72Y104_SLICE_X109Y104_B1 = CLBLM_L_X70Y105_SLICE_X104Y105_BO6;
  assign CLBLM_L_X72Y104_SLICE_X109Y104_B2 = CLBLM_L_X72Y104_SLICE_X109Y104_BQ;
  assign CLBLM_L_X72Y104_SLICE_X109Y104_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y114_SLICE_X105Y114_A6 = 1'b1;
  assign CLBLM_L_X72Y104_SLICE_X109Y104_B4 = CLBLM_L_X72Y104_SLICE_X109Y104_B5Q;
  assign CLBLM_L_X72Y104_SLICE_X109Y104_B5 = CLBLM_L_X72Y104_SLICE_X109Y104_C5Q;
  assign CLBLM_L_X72Y104_SLICE_X109Y104_B6 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X120Y128_B1 = 1'b1;
  assign CLBLM_L_X72Y104_SLICE_X109Y104_C1 = CLBLM_L_X72Y104_SLICE_X109Y104_C5Q;
  assign CLBLM_L_X72Y104_SLICE_X109Y104_C2 = CLBLM_L_X72Y104_SLICE_X109Y104_CQ;
  assign CLBLM_L_X72Y104_SLICE_X109Y104_C3 = CLBLL_R_X73Y104_SLICE_X110Y104_A5Q;
  assign CLBLM_L_X72Y104_SLICE_X109Y104_C4 = CLBLL_R_X73Y104_SLICE_X111Y104_DO6;
  assign CLBLM_L_X72Y104_SLICE_X109Y104_C5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y104_SLICE_X109Y104_C6 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X120Y128_C1 = 1'b1;
  assign CLBLM_L_X72Y104_SLICE_X109Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X78Y128_SLICE_X120Y128_C2 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X120Y128_C3 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X120Y128_C4 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X120Y128_C5 = 1'b1;
  assign CLBLM_L_X72Y104_SLICE_X109Y104_D1 = CLBLM_L_X72Y104_SLICE_X109Y104_C5Q;
  assign CLBLM_L_X72Y104_SLICE_X109Y104_D2 = CLBLM_L_X72Y104_SLICE_X109Y104_CQ;
  assign CLBLM_L_X72Y104_SLICE_X109Y104_D3 = CLBLM_L_X72Y104_SLICE_X109Y104_BQ;
  assign CLBLM_L_X70Y114_SLICE_X105Y114_B1 = 1'b1;
  assign CLBLM_L_X72Y104_SLICE_X109Y104_D4 = CLBLM_L_X70Y105_SLICE_X105Y105_BQ;
  assign CLBLM_L_X72Y104_SLICE_X109Y104_D5 = CLBLM_L_X72Y104_SLICE_X109Y104_B5Q;
  assign CLBLM_L_X72Y104_SLICE_X109Y104_D6 = CLBLM_L_X70Y105_SLICE_X104Y105_BO6;
  assign CLBLM_L_X72Y104_SLICE_X109Y104_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X78Y128_SLICE_X120Y128_D1 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X120Y128_D2 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X120Y128_D3 = 1'b1;
  assign CLBLM_L_X72Y104_SLICE_X108Y104_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y104_SLICE_X108Y104_A2 = CLBLL_R_X73Y103_SLICE_X111Y103_BO6;
  assign CLBLM_L_X72Y104_SLICE_X108Y104_A3 = CLBLM_L_X72Y104_SLICE_X108Y104_AQ;
  assign CLBLM_L_X72Y104_SLICE_X108Y104_A4 = CLBLM_L_X72Y105_SLICE_X108Y105_BQ;
  assign CLBLM_L_X72Y104_SLICE_X108Y104_A5 = CLBLM_L_X72Y103_SLICE_X109Y103_AO6;
  assign CLBLM_L_X70Y114_SLICE_X105Y114_B4 = 1'b1;
  assign CLBLM_L_X72Y104_SLICE_X108Y104_A6 = 1'b1;
  assign CLBLM_L_X78Y128_SLICE_X120Y128_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X103Y76_SLICE_X162Y76_B1 = 1'b1;
  assign CLBLM_L_X72Y104_SLICE_X108Y104_B1 = CLBLM_L_X72Y105_SLICE_X108Y105_A5Q;
  assign CLBLM_L_X72Y104_SLICE_X108Y104_B2 = CLBLM_L_X72Y104_SLICE_X108Y104_BQ;
  assign CLBLM_L_X72Y104_SLICE_X108Y104_B3 = CLBLM_L_X72Y104_SLICE_X109Y104_A5Q;
  assign CLBLM_L_X72Y104_SLICE_X108Y104_B4 = CLBLL_R_X73Y104_SLICE_X110Y104_BQ;
  assign CLBLM_L_X70Y114_SLICE_X105Y114_B6 = 1'b1;
  assign CLBLM_L_X72Y104_SLICE_X108Y104_B5 = CLBLM_L_X72Y103_SLICE_X108Y103_A5Q;
  assign CLBLM_L_X72Y104_SLICE_X108Y104_B6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X103Y76_SLICE_X162Y76_BX = CLBLM_R_X103Y76_SLICE_X163Y76_AQ;
  assign CLBLM_R_X103Y76_SLICE_X162Y76_C1 = 1'b1;
  assign CLBLM_R_X103Y76_SLICE_X162Y76_C2 = 1'b1;
  assign CLBLM_L_X72Y104_SLICE_X108Y104_C1 = CLBLM_L_X72Y104_SLICE_X108Y104_BQ;
  assign CLBLM_L_X72Y104_SLICE_X108Y104_C2 = CLBLM_L_X72Y104_SLICE_X108Y104_CQ;
  assign CLBLM_L_X72Y104_SLICE_X108Y104_C3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y104_SLICE_X108Y104_C4 = 1'b1;
  assign CLBLM_L_X72Y104_SLICE_X108Y104_C5 = CLBLM_L_X72Y105_SLICE_X108Y105_A5Q;
  assign CLBLM_L_X72Y104_SLICE_X108Y104_C6 = CLBLL_R_X73Y104_SLICE_X110Y104_BO5;
  assign CLBLM_R_X103Y76_SLICE_X162Y76_D1 = 1'b1;
  assign CLBLM_R_X103Y76_SLICE_X162Y76_D2 = 1'b1;
  assign CLBLM_R_X103Y76_SLICE_X162Y76_D3 = 1'b1;
  assign CLBLM_L_X72Y104_SLICE_X108Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X103Y76_SLICE_X162Y76_D4 = 1'b1;
  assign CLBLM_R_X103Y76_SLICE_X162Y76_D5 = 1'b1;
  assign CLBLM_R_X103Y76_SLICE_X162Y76_D6 = 1'b1;
  assign CLBLM_L_X72Y104_SLICE_X108Y104_D1 = CLBLL_R_X73Y104_SLICE_X111Y104_BQ;
  assign CLBLM_L_X72Y104_SLICE_X108Y104_D2 = CLBLM_L_X70Y105_SLICE_X104Y105_BO6;
  assign CLBLM_L_X72Y104_SLICE_X108Y104_D3 = CLBLM_L_X72Y104_SLICE_X108Y104_DQ;
  assign CLBLM_L_X70Y114_SLICE_X105Y114_C1 = 1'b1;
  assign CLBLM_L_X72Y104_SLICE_X108Y104_D4 = CLBLL_R_X73Y103_SLICE_X111Y103_BO6;
  assign CLBLM_L_X72Y104_SLICE_X108Y104_D5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y104_SLICE_X108Y104_D6 = 1'b1;
  assign CLBLM_R_X103Y76_SLICE_X162Y76_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X70Y114_SLICE_X105Y114_C2 = 1'b1;
  assign CLBLM_L_X72Y104_SLICE_X108Y104_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X70Y114_SLICE_X105Y114_C3 = 1'b1;
  assign CLBLM_L_X70Y114_SLICE_X105Y114_C4 = 1'b1;
  assign CLBLM_L_X70Y114_SLICE_X105Y114_C5 = 1'b1;
  assign CLBLM_L_X70Y114_SLICE_X105Y114_C6 = 1'b1;
  assign CLBLL_R_X71Y130_SLICE_X106Y130_A1 = CLBLM_L_X72Y132_SLICE_X109Y132_AO6;
  assign CLBLL_R_X71Y130_SLICE_X106Y130_A2 = CLBLL_R_X71Y129_SLICE_X107Y129_AQ;
  assign CLBLL_R_X71Y130_SLICE_X106Y130_A3 = CLBLL_R_X71Y130_SLICE_X106Y130_AQ;
  assign CLBLL_R_X71Y130_SLICE_X106Y130_A4 = CLBLM_L_X70Y130_SLICE_X105Y130_AQ;
  assign CLBLL_R_X71Y130_SLICE_X106Y130_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y130_SLICE_X106Y130_A6 = 1'b1;
  assign CLBLL_R_X71Y130_SLICE_X106Y130_B1 = CLBLL_R_X71Y130_SLICE_X106Y130_CQ;
  assign CLBLL_R_X71Y130_SLICE_X106Y130_B2 = CLBLL_R_X71Y130_SLICE_X106Y130_BQ;
  assign CLBLL_R_X71Y130_SLICE_X106Y130_B3 = CLBLM_L_X72Y129_SLICE_X108Y129_AQ;
  assign CLBLL_R_X71Y130_SLICE_X106Y130_B4 = CLBLL_R_X71Y125_SLICE_X107Y125_BO6;
  assign CLBLL_R_X71Y130_SLICE_X106Y130_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y130_SLICE_X106Y130_B6 = CLBLL_R_X71Y129_SLICE_X106Y129_AQ;
  assign CLBLL_R_X71Y130_SLICE_X106Y130_C1 = CLBLL_R_X71Y131_SLICE_X107Y131_AQ;
  assign CLBLL_R_X71Y130_SLICE_X106Y130_C2 = CLBLM_L_X72Y130_SLICE_X108Y130_AO6;
  assign CLBLL_R_X71Y130_SLICE_X106Y130_C3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y130_SLICE_X106Y130_C4 = CLBLL_R_X71Y129_SLICE_X106Y129_AO6;
  assign CLBLL_R_X71Y130_SLICE_X106Y130_C5 = CLBLL_R_X71Y130_SLICE_X106Y130_CQ;
  assign CLBLL_R_X71Y130_SLICE_X106Y130_C6 = CLBLL_R_X71Y125_SLICE_X107Y125_BO6;
  assign CLBLL_R_X71Y130_SLICE_X106Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X70Y114_SLICE_X105Y114_D1 = 1'b1;
  assign CLBLL_R_X71Y130_SLICE_X106Y130_D1 = CLBLM_L_X70Y129_SLICE_X104Y129_CQ;
  assign CLBLL_R_X71Y130_SLICE_X106Y130_D2 = CLBLL_R_X71Y126_SLICE_X107Y126_DO6;
  assign CLBLL_R_X71Y130_SLICE_X106Y130_D3 = CLBLM_L_X72Y130_SLICE_X108Y130_CQ;
  assign CLBLL_R_X71Y130_SLICE_X106Y130_D4 = CLBLL_R_X71Y132_SLICE_X106Y132_BQ;
  assign CLBLL_R_X71Y130_SLICE_X106Y130_D5 = CLBLM_L_X70Y133_SLICE_X105Y133_DQ;
  assign CLBLL_R_X71Y130_SLICE_X106Y130_D6 = 1'b1;
  assign CLBLM_L_X70Y114_SLICE_X105Y114_D2 = 1'b1;
  assign CLBLL_R_X71Y130_SLICE_X106Y130_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X70Y114_SLICE_X105Y114_D3 = 1'b1;
  assign CLBLM_L_X70Y114_SLICE_X105Y114_D4 = 1'b1;
  assign CLBLM_L_X70Y114_SLICE_X105Y114_D5 = 1'b1;
  assign CLBLM_L_X70Y114_SLICE_X105Y114_D6 = 1'b1;
  assign CLBLL_R_X71Y130_SLICE_X107Y130_A1 = CLBLL_R_X71Y129_SLICE_X106Y129_AQ;
  assign CLBLL_R_X71Y130_SLICE_X107Y130_A2 = CLBLM_L_X72Y131_SLICE_X109Y131_BQ;
  assign CLBLL_R_X71Y130_SLICE_X107Y130_A3 = CLBLL_R_X71Y130_SLICE_X106Y130_BQ;
  assign CLBLL_R_X71Y130_SLICE_X107Y130_A4 = CLBLL_R_X71Y130_SLICE_X107Y130_BO6;
  assign CLBLL_R_X71Y130_SLICE_X107Y130_A5 = CLBLL_R_X71Y131_SLICE_X107Y131_AQ;
  assign CLBLL_R_X71Y130_SLICE_X107Y130_A6 = CLBLL_R_X71Y130_SLICE_X107Y130_CO6;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_D4 = 1'b1;
  assign CLBLL_R_X71Y130_SLICE_X107Y130_AX = CLBLM_L_X72Y131_SLICE_X108Y131_AQ;
  assign CLBLL_R_X71Y130_SLICE_X107Y130_B1 = CLBLL_R_X71Y129_SLICE_X106Y129_AQ;
  assign CLBLL_R_X71Y130_SLICE_X107Y130_B2 = CLBLM_L_X72Y131_SLICE_X108Y131_BQ;
  assign CLBLL_R_X71Y130_SLICE_X107Y130_B3 = CLBLM_L_X72Y129_SLICE_X108Y129_AQ;
  assign CLBLL_R_X71Y130_SLICE_X107Y130_B4 = CLBLL_R_X71Y130_SLICE_X106Y130_BQ;
  assign CLBLL_R_X71Y130_SLICE_X107Y130_B5 = 1'b1;
  assign CLBLL_R_X71Y130_SLICE_X107Y130_B6 = CLBLL_R_X71Y131_SLICE_X107Y131_CQ;
  assign CLBLL_R_X71Y130_SLICE_X107Y130_BX = CLBLL_R_X71Y132_SLICE_X106Y132_AQ;
  assign CLBLL_R_X71Y130_SLICE_X107Y130_C1 = CLBLM_L_X72Y129_SLICE_X108Y129_AQ;
  assign CLBLL_R_X71Y130_SLICE_X107Y130_C2 = CLBLL_R_X71Y129_SLICE_X106Y129_AQ;
  assign CLBLL_R_X71Y130_SLICE_X107Y130_C3 = 1'b1;
  assign CLBLL_R_X71Y130_SLICE_X107Y130_C4 = CLBLM_L_X72Y131_SLICE_X108Y131_CQ;
  assign CLBLL_R_X71Y130_SLICE_X107Y130_C5 = CLBLL_R_X71Y131_SLICE_X107Y131_BQ;
  assign CLBLL_R_X71Y130_SLICE_X107Y130_C6 = CLBLL_R_X71Y130_SLICE_X106Y130_BQ;
  assign CLBLL_R_X71Y130_SLICE_X107Y130_CE = CLBLM_L_X76Y109_SLICE_X116Y109_AO6;
  assign CLBLL_R_X71Y130_SLICE_X107Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_D5 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_A4 = CLBLL_R_X77Y130_SLICE_X118Y130_AQ;
  assign CLBLL_R_X71Y130_SLICE_X107Y130_D1 = CLBLL_R_X71Y133_SLICE_X107Y133_BQ;
  assign CLBLL_R_X71Y130_SLICE_X107Y130_D2 = CLBLM_L_X70Y130_SLICE_X104Y130_DQ;
  assign CLBLL_R_X71Y130_SLICE_X107Y130_D3 = CLBLL_R_X71Y131_SLICE_X106Y131_CQ;
  assign CLBLL_R_X71Y130_SLICE_X107Y130_D4 = 1'b1;
  assign CLBLL_R_X71Y130_SLICE_X107Y130_D5 = 1'b1;
  assign CLBLL_R_X71Y130_SLICE_X107Y130_D6 = CLBLL_R_X71Y134_SLICE_X107Y134_BQ;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_A5 = CLBLL_R_X77Y128_SLICE_X118Y128_BQ;
  assign CLBLL_R_X71Y130_SLICE_X107Y130_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_A6 = CLBLL_R_X77Y128_SLICE_X119Y128_A5Q;
  assign CLBLM_L_X70Y114_SLICE_X104Y114_A6 = CLBLM_L_X70Y114_SLICE_X104Y114_A5Q;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_D6 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_A1 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_A2 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_A3 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_A4 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_A5 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_A6 = 1'b1;
  assign CLBLM_L_X70Y114_SLICE_X104Y114_AX = CLBLL_R_X71Y117_SLICE_X106Y117_B5Q;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_B1 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_B2 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_B2 = CLBLL_R_X77Y128_SLICE_X119Y128_CQ;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_B3 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_B4 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_B5 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_B6 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_B3 = CLBLL_R_X77Y128_SLICE_X118Y128_BQ;
  assign CLBLM_L_X70Y114_SLICE_X104Y114_B1 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_C1 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_C2 = 1'b1;
  assign CLBLM_L_X76Y111_SLICE_X116Y111_D4 = 1'b1;
  assign CLBLM_L_X70Y114_SLICE_X104Y114_B2 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_B4 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_C3 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_C4 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_B5 = CLBLM_L_X78Y128_SLICE_X120Y128_AQ;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_C5 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_C6 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_B6 = 1'b1;
  assign CLBLM_L_X70Y114_SLICE_X104Y114_B4 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_D1 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_D2 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_D3 = 1'b1;
  assign CLBLM_L_X70Y114_SLICE_X104Y114_B5 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_D4 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_D5 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_D6 = 1'b1;
  assign CLBLM_L_X70Y114_SLICE_X104Y114_B6 = 1'b1;
  assign CLBLM_L_X72Y105_SLICE_X109Y105_A1 = CLBLM_L_X72Y104_SLICE_X109Y104_A5Q;
  assign CLBLM_L_X72Y105_SLICE_X109Y105_A2 = CLBLM_L_X72Y103_SLICE_X108Y103_A5Q;
  assign CLBLM_L_X72Y105_SLICE_X109Y105_A3 = CLBLM_L_X72Y105_SLICE_X109Y105_AQ;
  assign CLBLM_L_X72Y105_SLICE_X109Y105_A4 = CLBLL_R_X73Y104_SLICE_X110Y104_BQ;
  assign CLBLM_L_X72Y105_SLICE_X109Y105_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y105_SLICE_X109Y105_A6 = CLBLM_L_X72Y105_SLICE_X108Y105_CQ;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_A1 = CLBLL_R_X77Y130_SLICE_X119Y130_AQ;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_A2 = CLBLM_L_X78Y131_SLICE_X120Y131_AQ;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_A3 = CLBLL_R_X77Y128_SLICE_X118Y128_AQ;
  assign CLBLM_L_X72Y105_SLICE_X109Y105_B1 = CLBLM_L_X72Y105_SLICE_X109Y105_B5Q;
  assign CLBLM_L_X72Y105_SLICE_X109Y105_B2 = CLBLM_L_X72Y105_SLICE_X109Y105_BQ;
  assign CLBLM_L_X72Y105_SLICE_X109Y105_B3 = CLBLM_L_X72Y105_SLICE_X109Y105_AQ;
  assign CLBLM_L_X72Y105_SLICE_X109Y105_B4 = CLBLM_L_X72Y103_SLICE_X109Y103_CO6;
  assign CLBLM_L_X72Y105_SLICE_X109Y105_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y105_SLICE_X109Y105_B6 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_B1 = 1'b1;
  assign CLBLM_L_X72Y105_SLICE_X109Y105_C1 = 1'b1;
  assign CLBLM_L_X72Y105_SLICE_X109Y105_C2 = 1'b1;
  assign CLBLM_L_X72Y105_SLICE_X109Y105_C3 = 1'b1;
  assign CLBLM_L_X72Y105_SLICE_X109Y105_C4 = 1'b1;
  assign CLBLM_L_X72Y105_SLICE_X109Y105_C5 = 1'b1;
  assign CLBLM_L_X72Y105_SLICE_X109Y105_C6 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_C1 = 1'b1;
  assign CLBLM_L_X72Y105_SLICE_X109Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_C2 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_C3 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_C4 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_C5 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_C6 = 1'b1;
  assign CLBLM_L_X72Y105_SLICE_X109Y105_D1 = 1'b1;
  assign CLBLM_L_X72Y105_SLICE_X109Y105_D2 = 1'b1;
  assign CLBLM_L_X72Y105_SLICE_X109Y105_D3 = 1'b1;
  assign CLBLM_L_X72Y105_SLICE_X109Y105_D4 = 1'b1;
  assign CLBLM_L_X72Y105_SLICE_X109Y105_D5 = 1'b1;
  assign CLBLM_L_X72Y105_SLICE_X109Y105_D6 = 1'b1;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_DX = CLBLM_L_X72Y121_SLICE_X108Y121_CQ;
  assign CLBLM_L_X72Y105_SLICE_X109Y105_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X70Y114_SLICE_X104Y114_C5 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_D1 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_D2 = 1'b1;
  assign CLBLM_L_X72Y105_SLICE_X108Y105_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y105_SLICE_X108Y105_A2 = CLBLM_L_X72Y105_SLICE_X109Y105_B5Q;
  assign CLBLM_L_X70Y114_SLICE_X104Y114_C6 = 1'b1;
  assign CLBLM_L_X72Y105_SLICE_X108Y105_A3 = CLBLM_L_X72Y103_SLICE_X109Y103_AO6;
  assign CLBLM_L_X72Y105_SLICE_X108Y105_A4 = CLBLM_L_X72Y128_SLICE_X109Y128_AQ;
  assign CLBLM_L_X72Y105_SLICE_X108Y105_A5 = CLBLM_L_X72Y105_SLICE_X108Y105_A5Q;
  assign CLBLM_L_X72Y105_SLICE_X108Y105_A6 = 1'b1;
  assign CLBLM_L_X72Y105_SLICE_X108Y105_B1 = CLBLM_L_X72Y103_SLICE_X108Y103_A5Q;
  assign CLBLM_L_X72Y105_SLICE_X108Y105_B2 = CLBLM_L_X72Y105_SLICE_X108Y105_BQ;
  assign CLBLM_L_X72Y105_SLICE_X108Y105_B3 = CLBLM_L_X72Y105_SLICE_X108Y105_DQ;
  assign CLBLM_L_X72Y105_SLICE_X108Y105_B4 = CLBLL_R_X73Y104_SLICE_X110Y104_BQ;
  assign CLBLM_L_X72Y105_SLICE_X108Y105_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y105_SLICE_X108Y105_B6 = CLBLM_L_X72Y104_SLICE_X109Y104_A5Q;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y105_SLICE_X108Y105_C1 = CLBLM_L_X72Y104_SLICE_X108Y104_AQ;
  assign CLBLM_L_X72Y105_SLICE_X108Y105_C2 = CLBLM_L_X72Y105_SLICE_X108Y105_CQ;
  assign CLBLM_L_X72Y105_SLICE_X108Y105_C3 = CLBLM_L_X72Y105_SLICE_X108Y105_BQ;
  assign CLBLM_L_X72Y105_SLICE_X108Y105_C4 = 1'b1;
  assign CLBLM_L_X72Y105_SLICE_X108Y105_C5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y105_SLICE_X108Y105_C6 = CLBLM_L_X72Y103_SLICE_X109Y103_CO6;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_D3 = 1'b1;
  assign CLBLM_L_X72Y105_SLICE_X108Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_D4 = 1'b1;
  assign CLBLM_L_X72Y105_SLICE_X108Y105_D1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y105_SLICE_X108Y105_D2 = CLBLL_R_X73Y104_SLICE_X110Y104_BQ;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_D5 = 1'b1;
  assign CLBLM_L_X72Y105_SLICE_X108Y105_D3 = CLBLM_L_X72Y105_SLICE_X108Y105_DQ;
  assign CLBLM_L_X72Y105_SLICE_X108Y105_D4 = CLBLM_L_X72Y104_SLICE_X109Y104_A5Q;
  assign CLBLM_L_X72Y105_SLICE_X108Y105_D5 = CLBLL_R_X79Y99_SLICE_X122Y99_AO6;
  assign CLBLL_R_X77Y104_SLICE_X118Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_D6 = 1'b1;
  assign CLBLM_L_X72Y105_SLICE_X108Y105_D6 = CLBLM_L_X72Y103_SLICE_X108Y103_A5Q;
  assign CLBLM_L_X72Y105_SLICE_X108Y105_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_D3 = 1'b1;
  assign CLBLM_L_X70Y110_SLICE_X105Y110_B5 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_D4 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_D5 = 1'b1;
  assign CLBLM_L_X70Y114_SLICE_X104Y114_D3 = 1'b1;
  assign CLBLM_R_X67Y115_SLICE_X100Y115_D2 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_D6 = 1'b1;
  assign CLBLM_L_X70Y114_SLICE_X104Y114_D4 = 1'b1;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1 = RIOB33_X105Y57_IOB_X1Y57_I;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_A1 = CLBLL_R_X71Y131_SLICE_X107Y131_A5Q;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_A2 = CLBLL_R_X71Y132_SLICE_X107Y132_BQ;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_A3 = CLBLL_R_X71Y131_SLICE_X106Y131_AQ;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_A4 = CLBLL_R_X71Y125_SLICE_X107Y125_CO6;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_A6 = CLBLL_R_X71Y132_SLICE_X106Y132_AQ;
  assign CLBLM_L_X70Y114_SLICE_X104Y114_D5 = 1'b1;
  assign CLBLM_L_X70Y110_SLICE_X105Y110_B6 = 1'b1;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1 = 1'b1;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_B1 = CLBLL_R_X71Y131_SLICE_X107Y131_A5Q;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_B2 = CLBLL_R_X71Y131_SLICE_X106Y131_BQ;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_B3 = CLBLL_R_X71Y131_SLICE_X106Y131_AQ;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_B4 = CLBLL_R_X71Y125_SLICE_X107Y125_CO6;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_B6 = CLBLL_R_X71Y132_SLICE_X106Y132_DQ;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_C2 = CLBLL_R_X71Y131_SLICE_X106Y131_CQ;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_C3 = CLBLL_R_X71Y132_SLICE_X106Y132_DQ;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_C4 = CLBLL_R_X71Y131_SLICE_X106Y131_BQ;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_C5 = CLBLL_R_X71Y131_SLICE_X106Y131_DO6;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_C6 = 1'b1;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_D1 = 1'b1;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_D2 = 1'b1;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_D3 = CLBLL_R_X71Y131_SLICE_X106Y131_AQ;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_D4 = 1'b1;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_D5 = CLBLL_R_X71Y131_SLICE_X107Y131_A5Q;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_D6 = CLBLL_R_X71Y125_SLICE_X107Y125_CO6;
  assign LIOB33_X0Y55_IOB_X0Y56_O = CLBLM_L_X62Y92_SLICE_X92Y92_BQ;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_A1 = CLBLM_L_X72Y131_SLICE_X108Y131_A5Q;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_A2 = CLBLL_R_X71Y131_SLICE_X107Y131_BQ;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_A3 = CLBLL_R_X71Y131_SLICE_X107Y131_AQ;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_A4 = CLBLM_L_X72Y131_SLICE_X109Y131_AO6;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_A6 = CLBLM_L_X72Y134_SLICE_X109Y134_AO5;
  assign CLBLM_L_X72Y109_SLICE_X109Y109_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_AX = CLBLL_R_X71Y131_SLICE_X107Y131_DO5;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_B4 = CLBLM_L_X64Y102_SLICE_X96Y102_A5Q;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_B1 = CLBLM_L_X72Y133_SLICE_X109Y133_DO6;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_B2 = CLBLL_R_X71Y131_SLICE_X107Y131_BQ;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_B3 = CLBLL_R_X71Y131_SLICE_X107Y131_CQ;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_B4 = CLBLM_L_X72Y130_SLICE_X108Y130_AO6;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_B6 = CLBLM_L_X72Y134_SLICE_X109Y134_AO5;
  assign CLBLM_L_X60Y94_SLICE_X91Y94_C1 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_B6 = CLBLM_L_X64Y104_SLICE_X96Y104_DQ;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_C2 = CLBLM_L_X72Y134_SLICE_X109Y134_AO5;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_C3 = CLBLM_L_X72Y131_SLICE_X108Y131_CQ;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_C4 = CLBLM_L_X72Y131_SLICE_X108Y131_DO5;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_C5 = CLBLM_L_X72Y133_SLICE_X109Y133_DO6;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_C6 = CLBLL_R_X71Y131_SLICE_X107Y131_CQ;
  assign CLBLM_L_X72Y109_SLICE_X109Y109_C4 = CLBLM_L_X72Y109_SLICE_X109Y109_BQ;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X72Y109_SLICE_X109Y109_C6 = 1'b1;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_D1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X60Y94_SLICE_X91Y94_C5 = 1'b1;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_D2 = CLBLL_R_X71Y132_SLICE_X106Y132_AQ;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_D3 = CLBLL_R_X71Y130_SLICE_X107Y130_BQ;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_D4 = CLBLL_R_X71Y131_SLICE_X107Y131_A5Q;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_D5 = CLBLL_R_X71Y125_SLICE_X107Y125_CO6;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_D6 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_A1 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_A2 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_A3 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_A4 = 1'b1;
  assign CLBLL_R_X79Y127_SLICE_X122Y127_A2 = 1'b1;
  assign CLBLL_R_X79Y127_SLICE_X122Y127_A3 = CLBLL_R_X79Y127_SLICE_X122Y127_AQ;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_A5 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_A6 = CLBLM_R_X53Y122_SLICE_X80Y122_AQ;
  assign CLBLL_R_X79Y127_SLICE_X122Y127_A6 = CLBLL_R_X79Y127_SLICE_X122Y127_A5Q;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X79Y127_SLICE_X122Y127_A1 = CLBLL_R_X77Y125_SLICE_X118Y125_BO5;
  assign CLBLL_R_X79Y127_SLICE_X122Y127_B1 = CLBLL_R_X77Y125_SLICE_X118Y125_BO5;
  assign CLBLL_R_X79Y127_SLICE_X122Y127_B2 = CLBLL_R_X79Y127_SLICE_X122Y127_BQ;
  assign CLBLL_R_X79Y127_SLICE_X122Y127_B3 = CLBLL_R_X83Y130_SLICE_X130Y130_DQ;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_B1 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_B2 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_B3 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_B4 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_B5 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_B6 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_C1 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_C2 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_C3 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_C4 = 1'b1;
  assign CLBLL_R_X79Y127_SLICE_X122Y127_C5 = CLBLL_R_X77Y125_SLICE_X118Y125_BO5;
  assign CLBLL_R_X79Y127_SLICE_X122Y127_C6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_C5 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_C6 = 1'b1;
  assign CLBLL_R_X79Y127_SLICE_X122Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X79Y127_SLICE_X122Y127_C1 = 1'b1;
  assign CLBLL_R_X79Y127_SLICE_X122Y127_C2 = CLBLL_R_X79Y127_SLICE_X122Y127_CQ;
  assign CLBLL_R_X79Y127_SLICE_X122Y127_C3 = CLBLL_R_X79Y128_SLICE_X122Y128_BQ;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_D1 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_D2 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_D3 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_D4 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_D5 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_D6 = 1'b1;
  assign CLBLL_R_X79Y127_SLICE_X122Y127_D1 = CLBLL_R_X79Y128_SLICE_X122Y128_AQ;
  assign CLBLL_R_X79Y127_SLICE_X122Y127_D2 = CLBLL_R_X79Y127_SLICE_X122Y127_CQ;
  assign CLBLL_R_X79Y127_SLICE_X122Y127_D3 = 1'b1;
  assign CLBLL_R_X79Y127_SLICE_X122Y127_D4 = CLBLL_R_X79Y128_SLICE_X122Y128_CQ;
  assign CLBLL_R_X79Y127_SLICE_X122Y127_D5 = CLBLL_R_X79Y128_SLICE_X122Y128_DQ;
  assign CLBLL_R_X79Y127_SLICE_X122Y127_D6 = 1'b1;
  assign CLBLL_R_X79Y127_SLICE_X122Y127_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X78Y130_SLICE_X121Y130_B6 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_B3 = CLBLM_L_X70Y105_SLICE_X105Y105_AQ;
  assign CLBLM_L_X78Y130_SLICE_X121Y130_C1 = 1'b1;
  assign CLBLM_L_X78Y130_SLICE_X121Y130_C2 = 1'b1;
  assign CLBLM_L_X78Y130_SLICE_X121Y130_C3 = 1'b1;
  assign CLBLM_L_X78Y130_SLICE_X121Y130_C4 = 1'b1;
  assign CLBLM_L_X78Y130_SLICE_X121Y130_C5 = 1'b1;
  assign CLBLM_L_X78Y130_SLICE_X121Y130_C6 = 1'b1;
  assign CLBLM_L_X60Y94_SLICE_X91Y94_D4 = 1'b1;
  assign CLBLM_L_X72Y109_SLICE_X109Y109_D6 = CLBLM_L_X72Y111_SLICE_X109Y111_BQ;
  assign CLBLM_L_X78Y130_SLICE_X121Y130_D1 = 1'b1;
  assign CLBLM_L_X78Y130_SLICE_X121Y130_D2 = 1'b1;
  assign CLBLM_L_X78Y130_SLICE_X121Y130_D3 = 1'b1;
  assign CLBLM_L_X60Y94_SLICE_X91Y94_D5 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_A1 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_A2 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_A3 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_A4 = 1'b1;
  assign CLBLM_L_X60Y94_SLICE_X91Y94_D6 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_A5 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_A6 = 1'b1;
  assign CLBLL_R_X79Y127_SLICE_X123Y127_A4 = 1'b1;
  assign CLBLL_R_X79Y127_SLICE_X123Y127_A5 = 1'b1;
  assign CLBLL_R_X79Y127_SLICE_X123Y127_A6 = 1'b1;
  assign CLBLL_R_X79Y127_SLICE_X123Y127_A1 = 1'b1;
  assign CLBLL_R_X79Y127_SLICE_X123Y127_A2 = 1'b1;
  assign CLBLL_R_X79Y127_SLICE_X123Y127_B1 = 1'b1;
  assign CLBLL_R_X79Y127_SLICE_X123Y127_B2 = 1'b1;
  assign CLBLL_R_X79Y127_SLICE_X123Y127_B3 = 1'b1;
  assign CLBLL_R_X79Y127_SLICE_X123Y127_B4 = 1'b1;
  assign CLBLL_R_X79Y127_SLICE_X123Y127_B5 = 1'b1;
  assign CLBLL_R_X79Y127_SLICE_X123Y127_B6 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_B2 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_B3 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_B5 = 1'b1;
  assign CLBLL_R_X79Y127_SLICE_X123Y127_C1 = 1'b1;
  assign CLBLL_R_X79Y127_SLICE_X123Y127_C2 = 1'b1;
  assign CLBLL_R_X79Y127_SLICE_X123Y127_C3 = 1'b1;
  assign CLBLL_R_X79Y127_SLICE_X123Y127_C4 = 1'b1;
  assign CLBLL_R_X79Y127_SLICE_X123Y127_C5 = 1'b1;
  assign CLBLL_R_X79Y127_SLICE_X123Y127_C6 = 1'b1;
  assign CLBLL_R_X79Y127_SLICE_X123Y127_A3 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_C3 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_C4 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_C5 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_C6 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X118Y104_D4 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_D1 = 1'b1;
  assign CLBLL_R_X79Y127_SLICE_X123Y127_D1 = 1'b1;
  assign CLBLL_R_X79Y127_SLICE_X123Y127_D2 = 1'b1;
  assign CLBLL_R_X79Y127_SLICE_X123Y127_D3 = 1'b1;
  assign CLBLL_R_X79Y127_SLICE_X123Y127_D4 = 1'b1;
  assign CLBLL_R_X79Y127_SLICE_X123Y127_D5 = 1'b1;
  assign CLBLL_R_X79Y127_SLICE_X123Y127_D6 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_D2 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_D3 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_D5 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_D6 = 1'b1;
  assign CLBLM_L_X72Y106_SLICE_X109Y106_D1 = 1'b1;
  assign CLBLM_L_X72Y106_SLICE_X109Y106_D2 = 1'b1;
  assign CLBLM_L_X72Y106_SLICE_X109Y106_D3 = 1'b1;
  assign CLBLM_L_X72Y106_SLICE_X109Y106_D4 = 1'b1;
  assign CLBLM_L_X72Y106_SLICE_X109Y106_D5 = 1'b1;
  assign CLBLM_L_X72Y106_SLICE_X108Y106_A1 = CLBLM_L_X72Y106_SLICE_X108Y106_BO6;
  assign CLBLM_L_X72Y106_SLICE_X108Y106_A2 = CLBLM_L_X62Y90_SLICE_X92Y90_AQ;
  assign CLBLM_L_X72Y106_SLICE_X108Y106_A3 = CLBLM_L_X72Y106_SLICE_X108Y106_AQ;
  assign CLBLM_L_X72Y106_SLICE_X108Y106_A4 = CLBLM_L_X78Y106_SLICE_X120Y106_AQ;
  assign CLBLM_L_X72Y106_SLICE_X108Y106_A5 = CLBLM_L_X62Y92_SLICE_X92Y92_AQ;
  assign CLBLM_L_X72Y106_SLICE_X108Y106_A6 = CLBLM_L_X72Y106_SLICE_X108Y106_A5Q;
  assign CLBLM_L_X78Y130_SLICE_X120Y130_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y106_SLICE_X108Y106_AX = CLBLM_L_X78Y106_SLICE_X120Y106_AQ;
  assign CLBLM_R_X67Y115_SLICE_X100Y115_D4 = 1'b1;
  assign CLBLM_L_X72Y106_SLICE_X108Y106_B1 = CLBLM_L_X72Y107_SLICE_X109Y107_A5Q;
  assign CLBLM_L_X72Y106_SLICE_X108Y106_B2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y106_SLICE_X108Y106_B3 = CLBLM_L_X72Y106_SLICE_X108Y106_AQ;
  assign CLBLM_L_X72Y106_SLICE_X108Y106_B4 = CLBLM_L_X78Y106_SLICE_X120Y106_AQ;
  assign CLBLM_L_X72Y106_SLICE_X108Y106_B5 = CLBLM_L_X62Y92_SLICE_X92Y92_AQ;
  assign CLBLM_L_X72Y106_SLICE_X108Y106_B6 = CLBLM_L_X72Y106_SLICE_X108Y106_A5Q;
  assign CLBLM_L_X72Y106_SLICE_X108Y106_C1 = CLBLL_R_X73Y106_SLICE_X110Y106_BO6;
  assign CLBLM_L_X72Y106_SLICE_X108Y106_C2 = CLBLM_L_X72Y106_SLICE_X109Y106_CO6;
  assign CLBLM_L_X72Y106_SLICE_X108Y106_C3 = CLBLM_L_X70Y106_SLICE_X105Y106_CO6;
  assign CLBLM_L_X72Y106_SLICE_X108Y106_C4 = CLBLM_L_X72Y107_SLICE_X108Y107_CO6;
  assign CLBLM_L_X72Y106_SLICE_X108Y106_C5 = CLBLL_R_X73Y107_SLICE_X110Y107_DO6;
  assign CLBLM_L_X72Y106_SLICE_X108Y106_C6 = CLBLM_L_X72Y106_SLICE_X108Y106_DO6;
  assign CLBLL_R_X77Y104_SLICE_X118Y104_D6 = 1'b1;
  assign CLBLM_L_X72Y106_SLICE_X108Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X72Y106_SLICE_X108Y106_D1 = CLBLM_L_X72Y108_SLICE_X108Y108_AQ;
  assign CLBLM_L_X72Y106_SLICE_X108Y106_D2 = CLBLL_R_X71Y107_SLICE_X106Y107_C5Q;
  assign CLBLM_L_X72Y106_SLICE_X108Y106_D3 = CLBLL_R_X71Y107_SLICE_X107Y107_DO6;
  assign CLBLM_L_X72Y106_SLICE_X108Y106_D4 = CLBLL_R_X73Y108_SLICE_X110Y108_A5Q;
  assign CLBLM_L_X72Y106_SLICE_X108Y106_D5 = CLBLM_L_X72Y107_SLICE_X109Y107_A5Q;
  assign CLBLM_L_X72Y106_SLICE_X108Y106_D6 = CLBLL_R_X71Y107_SLICE_X106Y107_CQ;
  assign CLBLM_L_X72Y106_SLICE_X108Y106_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y109_SLICE_X108Y109_B6 = CLBLL_R_X71Y109_SLICE_X106Y109_B5Q;
  assign CLBLM_L_X60Y94_SLICE_X90Y94_B4 = 1'b1;
  assign CLBLM_L_X60Y94_SLICE_X90Y94_B5 = 1'b1;
  assign CLBLL_R_X71Y132_SLICE_X106Y132_A1 = 1'b1;
  assign CLBLL_R_X71Y132_SLICE_X106Y132_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y132_SLICE_X106Y132_A3 = CLBLL_R_X71Y132_SLICE_X106Y132_AQ;
  assign CLBLL_R_X71Y132_SLICE_X106Y132_A4 = CLBLL_R_X71Y131_SLICE_X106Y131_AQ;
  assign CLBLL_R_X71Y132_SLICE_X106Y132_A5 = CLBLL_R_X71Y125_SLICE_X107Y125_CO6;
  assign CLBLL_R_X71Y132_SLICE_X106Y132_A6 = 1'b1;
  assign CLBLM_R_X67Y110_SLICE_X100Y110_D3 = CLBLM_R_X67Y110_SLICE_X100Y110_AQ;
  assign CLBLL_R_X71Y132_SLICE_X106Y132_B1 = CLBLL_R_X71Y132_SLICE_X107Y132_DQ;
  assign CLBLL_R_X71Y132_SLICE_X106Y132_B2 = CLBLL_R_X71Y132_SLICE_X106Y132_BQ;
  assign CLBLL_R_X71Y132_SLICE_X106Y132_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y132_SLICE_X106Y132_B4 = CLBLM_L_X72Y133_SLICE_X109Y133_BQ;
  assign CLBLL_R_X71Y132_SLICE_X106Y132_B5 = 1'b1;
  assign CLBLL_R_X71Y132_SLICE_X106Y132_B6 = CLBLL_R_X71Y132_SLICE_X106Y132_AO5;
  assign CLBLL_R_X71Y132_SLICE_X106Y132_C1 = CLBLL_R_X71Y125_SLICE_X107Y125_CO6;
  assign CLBLL_R_X71Y132_SLICE_X106Y132_C2 = CLBLL_R_X71Y132_SLICE_X106Y132_CQ;
  assign CLBLL_R_X71Y132_SLICE_X106Y132_C3 = CLBLL_R_X71Y132_SLICE_X106Y132_BQ;
  assign CLBLL_R_X71Y132_SLICE_X106Y132_C4 = CLBLL_R_X71Y131_SLICE_X107Y131_A5Q;
  assign CLBLL_R_X71Y132_SLICE_X106Y132_C5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y132_SLICE_X106Y132_C6 = CLBLL_R_X71Y131_SLICE_X106Y131_AQ;
  assign CLBLL_R_X71Y132_SLICE_X106Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X71Y132_SLICE_X106Y132_D1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y132_SLICE_X106Y132_D2 = CLBLM_L_X72Y133_SLICE_X108Y133_AQ;
  assign CLBLL_R_X71Y132_SLICE_X106Y132_D3 = CLBLL_R_X71Y132_SLICE_X106Y132_DQ;
  assign CLBLL_R_X71Y132_SLICE_X106Y132_D4 = CLBLL_R_X73Y132_SLICE_X110Y132_BO6;
  assign CLBLL_R_X71Y132_SLICE_X106Y132_D5 = CLBLL_R_X71Y133_SLICE_X106Y133_DQ;
  assign CLBLL_R_X71Y132_SLICE_X106Y132_D6 = CLBLM_L_X72Y133_SLICE_X108Y133_A5Q;
  assign CLBLM_L_X72Y109_SLICE_X108Y109_C5 = 1'b1;
  assign CLBLM_L_X72Y109_SLICE_X108Y109_C6 = 1'b1;
  assign CLBLL_R_X71Y132_SLICE_X106Y132_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1 = CLBLM_R_X67Y105_SLICE_X101Y105_AO6;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1 = 1'b1;
  assign CLBLM_L_X72Y109_SLICE_X108Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X71Y132_SLICE_X107Y132_A1 = CLBLM_L_X72Y132_SLICE_X109Y132_AQ;
  assign CLBLL_R_X71Y132_SLICE_X107Y132_A2 = CLBLL_R_X73Y132_SLICE_X110Y132_BO6;
  assign CLBLL_R_X71Y132_SLICE_X107Y132_A3 = CLBLL_R_X71Y132_SLICE_X107Y132_AQ;
  assign CLBLL_R_X71Y132_SLICE_X107Y132_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y132_SLICE_X107Y132_A5 = CLBLM_L_X72Y133_SLICE_X108Y133_AQ;
  assign CLBLL_R_X71Y132_SLICE_X107Y132_A6 = 1'b1;
  assign CLBLL_R_X71Y132_SLICE_X107Y132_B1 = CLBLL_R_X71Y131_SLICE_X107Y131_DO6;
  assign CLBLL_R_X71Y132_SLICE_X107Y132_B2 = CLBLL_R_X71Y132_SLICE_X107Y132_BQ;
  assign CLBLL_R_X71Y132_SLICE_X107Y132_B3 = CLBLL_R_X71Y125_SLICE_X107Y125_CO6;
  assign CLBLL_R_X71Y132_SLICE_X107Y132_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y132_SLICE_X107Y132_B5 = CLBLL_R_X71Y132_SLICE_X107Y132_AO6;
  assign CLBLL_R_X71Y132_SLICE_X107Y132_B6 = CLBLM_L_X72Y132_SLICE_X108Y132_BQ;
  assign CLBLM_R_X67Y115_SLICE_X101Y115_A1 = 1'b1;
  assign CLBLM_R_X67Y115_SLICE_X101Y115_A2 = 1'b1;
  assign CLBLL_R_X71Y132_SLICE_X107Y132_C1 = CLBLM_L_X72Y132_SLICE_X109Y132_BO6;
  assign CLBLL_R_X71Y132_SLICE_X107Y132_C2 = CLBLL_R_X71Y132_SLICE_X107Y132_CQ;
  assign CLBLL_R_X71Y132_SLICE_X107Y132_C3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y132_SLICE_X107Y132_C4 = 1'b1;
  assign CLBLL_R_X71Y132_SLICE_X107Y132_C5 = CLBLL_R_X71Y131_SLICE_X107Y131_A5Q;
  assign CLBLL_R_X71Y132_SLICE_X107Y132_C6 = CLBLL_R_X71Y125_SLICE_X107Y125_CO6;
  assign CLBLM_R_X67Y115_SLICE_X101Y115_A3 = 1'b1;
  assign CLBLL_R_X71Y132_SLICE_X107Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X67Y115_SLICE_X101Y115_A4 = 1'b1;
  assign CLBLM_R_X67Y115_SLICE_X101Y115_A5 = 1'b1;
  assign CLBLL_R_X71Y132_SLICE_X107Y132_D1 = CLBLL_R_X71Y132_SLICE_X106Y132_AQ;
  assign CLBLL_R_X71Y132_SLICE_X107Y132_D2 = CLBLL_R_X71Y132_SLICE_X107Y132_CQ;
  assign CLBLL_R_X71Y132_SLICE_X107Y132_D3 = CLBLL_R_X71Y132_SLICE_X107Y132_DQ;
  assign CLBLL_R_X71Y132_SLICE_X107Y132_D4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y132_SLICE_X107Y132_D5 = CLBLL_R_X71Y131_SLICE_X106Y131_AQ;
  assign CLBLL_R_X71Y132_SLICE_X107Y132_D6 = CLBLL_R_X71Y125_SLICE_X107Y125_CO6;
  assign CLBLM_L_X74Y104_SLICE_X113Y104_A4 = 1'b1;
  assign CLBLM_L_X72Y109_SLICE_X108Y109_D4 = 1'b1;
  assign CLBLL_R_X71Y132_SLICE_X107Y132_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y104_SLICE_X113Y104_A5 = 1'b1;
  assign CLBLL_R_X79Y128_SLICE_X122Y128_A1 = CLBLL_R_X77Y125_SLICE_X118Y125_BO5;
  assign CLBLL_R_X79Y128_SLICE_X122Y128_A2 = CLBLL_R_X83Y132_SLICE_X130Y132_AQ;
  assign CLBLL_R_X79Y128_SLICE_X122Y128_A3 = CLBLL_R_X79Y128_SLICE_X122Y128_AQ;
  assign CLBLL_R_X79Y128_SLICE_X122Y128_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X79Y128_SLICE_X122Y128_A5 = CLBLL_R_X79Y128_SLICE_X122Y128_CQ;
  assign CLBLL_R_X79Y128_SLICE_X122Y128_A6 = 1'b1;
  assign CLBLM_L_X72Y109_SLICE_X108Y109_D5 = 1'b1;
  assign CLBLM_L_X74Y104_SLICE_X113Y104_A6 = 1'b1;
  assign CLBLL_R_X79Y128_SLICE_X122Y128_B1 = CLBLL_R_X77Y125_SLICE_X118Y125_BO5;
  assign CLBLL_R_X79Y128_SLICE_X122Y128_B2 = CLBLL_R_X79Y128_SLICE_X122Y128_BQ;
  assign CLBLL_R_X79Y128_SLICE_X122Y128_B3 = CLBLL_R_X79Y128_SLICE_X122Y128_DQ;
  assign CLBLL_R_X79Y128_SLICE_X122Y128_B4 = 1'b1;
  assign CLBLL_R_X79Y128_SLICE_X122Y128_B5 = CLBLL_R_X83Y130_SLICE_X130Y130_BQ;
  assign CLBLL_R_X79Y128_SLICE_X122Y128_B6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_B2 = CLBLM_L_X64Y98_SLICE_X96Y98_AO6;
  assign CLBLM_R_X67Y115_SLICE_X101Y115_B1 = 1'b1;
  assign CLBLL_R_X79Y128_SLICE_X122Y128_C1 = CLBLL_R_X79Y127_SLICE_X122Y127_AQ;
  assign CLBLL_R_X79Y128_SLICE_X122Y128_C2 = CLBLL_R_X79Y128_SLICE_X122Y128_CQ;
  assign CLBLL_R_X79Y128_SLICE_X122Y128_C3 = CLBLL_R_X77Y125_SLICE_X118Y125_BO5;
  assign CLBLL_R_X79Y128_SLICE_X122Y128_C4 = CLBLM_L_X82Y130_SLICE_X128Y130_AQ;
  assign CLBLL_R_X79Y128_SLICE_X122Y128_C5 = 1'b1;
  assign CLBLL_R_X79Y128_SLICE_X122Y128_C6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y115_SLICE_X101Y115_B2 = 1'b1;
  assign CLBLL_R_X79Y128_SLICE_X122Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X67Y115_SLICE_X101Y115_B3 = 1'b1;
  assign CLBLM_L_X74Y104_SLICE_X113Y104_B2 = 1'b1;
  assign CLBLM_L_X78Y131_SLICE_X121Y131_A1 = 1'b1;
  assign CLBLM_L_X78Y131_SLICE_X121Y131_A2 = 1'b1;
  assign CLBLM_L_X78Y131_SLICE_X121Y131_A3 = 1'b1;
  assign CLBLL_R_X79Y128_SLICE_X122Y128_D1 = CLBLL_R_X83Y130_SLICE_X130Y130_AQ;
  assign CLBLL_R_X79Y128_SLICE_X122Y128_D2 = CLBLL_R_X79Y128_SLICE_X122Y128_AQ;
  assign CLBLL_R_X79Y128_SLICE_X122Y128_D3 = CLBLL_R_X79Y128_SLICE_X122Y128_DQ;
  assign CLBLL_R_X79Y128_SLICE_X122Y128_D4 = 1'b1;
  assign CLBLL_R_X79Y128_SLICE_X122Y128_D5 = CLBLL_R_X77Y125_SLICE_X118Y125_BO5;
  assign CLBLL_R_X79Y128_SLICE_X122Y128_D6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y104_SLICE_X113Y104_B3 = 1'b1;
  assign CLBLM_L_X74Y104_SLICE_X113Y104_B4 = 1'b1;
  assign CLBLL_R_X79Y128_SLICE_X122Y128_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y104_SLICE_X113Y104_B5 = 1'b1;
  assign CLBLM_L_X78Y131_SLICE_X121Y131_B1 = 1'b1;
  assign CLBLM_L_X78Y131_SLICE_X121Y131_B2 = 1'b1;
  assign CLBLM_L_X78Y131_SLICE_X121Y131_B3 = 1'b1;
  assign CLBLM_L_X74Y104_SLICE_X113Y104_B6 = 1'b1;
  assign CLBLM_L_X78Y131_SLICE_X121Y131_B4 = 1'b1;
  assign CLBLM_L_X78Y131_SLICE_X121Y131_B5 = 1'b1;
  assign CLBLM_L_X78Y131_SLICE_X121Y131_B6 = 1'b1;
  assign CLBLM_L_X78Y131_SLICE_X121Y131_C1 = 1'b1;
  assign CLBLM_L_X78Y131_SLICE_X121Y131_C2 = 1'b1;
  assign CLBLM_L_X78Y131_SLICE_X121Y131_C3 = 1'b1;
  assign CLBLM_L_X78Y131_SLICE_X121Y131_C4 = 1'b1;
  assign CLBLM_L_X78Y131_SLICE_X121Y131_C5 = 1'b1;
  assign CLBLM_L_X78Y131_SLICE_X121Y131_C6 = 1'b1;
  assign CLBLM_L_X78Y131_SLICE_X121Y131_D1 = 1'b1;
  assign CLBLM_L_X78Y131_SLICE_X121Y131_D2 = 1'b1;
  assign CLBLM_L_X78Y131_SLICE_X121Y131_D3 = 1'b1;
  assign CLBLM_L_X78Y131_SLICE_X121Y131_D4 = 1'b1;
  assign CLBLL_R_X79Y128_SLICE_X123Y128_A1 = 1'b1;
  assign CLBLL_R_X79Y128_SLICE_X123Y128_A2 = 1'b1;
  assign CLBLL_R_X79Y128_SLICE_X123Y128_A3 = 1'b1;
  assign CLBLL_R_X79Y128_SLICE_X123Y128_A4 = 1'b1;
  assign CLBLL_R_X79Y128_SLICE_X123Y128_A5 = 1'b1;
  assign CLBLL_R_X79Y128_SLICE_X123Y128_A6 = 1'b1;
  assign CLBLM_L_X78Y131_SLICE_X121Y131_D5 = 1'b1;
  assign CLBLM_L_X78Y131_SLICE_X121Y131_D6 = 1'b1;
  assign CLBLM_L_X72Y107_SLICE_X109Y107_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X79Y128_SLICE_X123Y128_B1 = 1'b1;
  assign CLBLL_R_X79Y128_SLICE_X123Y128_B2 = 1'b1;
  assign CLBLL_R_X79Y128_SLICE_X123Y128_B3 = 1'b1;
  assign CLBLL_R_X79Y128_SLICE_X123Y128_B4 = 1'b1;
  assign CLBLL_R_X79Y128_SLICE_X123Y128_B5 = 1'b1;
  assign CLBLL_R_X79Y128_SLICE_X123Y128_B6 = 1'b1;
  assign CLBLM_L_X72Y107_SLICE_X109Y107_A2 = CLBLM_L_X72Y108_SLICE_X109Y108_CO5;
  assign CLBLM_L_X72Y107_SLICE_X109Y107_A3 = CLBLM_L_X72Y107_SLICE_X109Y107_AQ;
  assign CLBLM_L_X72Y107_SLICE_X109Y107_A4 = CLBLM_L_X72Y108_SLICE_X108Y108_BO6;
  assign CLBLL_R_X79Y128_SLICE_X123Y128_C1 = 1'b1;
  assign CLBLL_R_X79Y128_SLICE_X123Y128_C2 = 1'b1;
  assign CLBLL_R_X79Y128_SLICE_X123Y128_C3 = 1'b1;
  assign CLBLL_R_X79Y128_SLICE_X123Y128_C4 = 1'b1;
  assign CLBLL_R_X79Y128_SLICE_X123Y128_C5 = 1'b1;
  assign CLBLL_R_X79Y128_SLICE_X123Y128_C6 = 1'b1;
  assign CLBLM_L_X72Y107_SLICE_X109Y107_AX = CLBLM_L_X62Y92_SLICE_X92Y92_AQ;
  assign CLBLM_L_X72Y107_SLICE_X109Y107_B1 = CLBLL_R_X73Y108_SLICE_X110Y108_A5Q;
  assign CLBLM_L_X72Y107_SLICE_X109Y107_B2 = CLBLL_R_X71Y107_SLICE_X106Y107_CQ;
  assign CLBLM_L_X72Y107_SLICE_X109Y107_B3 = CLBLM_L_X72Y107_SLICE_X109Y107_AQ;
  assign CLBLM_L_X72Y107_SLICE_X109Y107_B4 = CLBLL_R_X71Y107_SLICE_X106Y107_C5Q;
  assign CLBLM_L_X72Y107_SLICE_X109Y107_B5 = CLBLM_L_X72Y106_SLICE_X108Y106_AQ;
  assign CLBLM_L_X72Y107_SLICE_X109Y107_B6 = 1'b1;
  assign CLBLM_L_X68Y95_SLICE_X103Y95_A2 = 1'b1;
  assign CLBLM_L_X68Y95_SLICE_X103Y95_A3 = 1'b1;
  assign CLBLM_L_X68Y95_SLICE_X103Y95_A1 = 1'b1;
  assign CLBLL_R_X79Y128_SLICE_X123Y128_D1 = 1'b1;
  assign CLBLL_R_X79Y128_SLICE_X123Y128_D2 = 1'b1;
  assign CLBLL_R_X79Y128_SLICE_X123Y128_D3 = 1'b1;
  assign CLBLL_R_X79Y128_SLICE_X123Y128_D4 = 1'b1;
  assign CLBLL_R_X79Y128_SLICE_X123Y128_D5 = 1'b1;
  assign CLBLL_R_X79Y128_SLICE_X123Y128_D6 = 1'b1;
  assign CLBLM_L_X68Y95_SLICE_X103Y95_A4 = 1'b1;
  assign CLBLM_L_X68Y95_SLICE_X103Y95_A5 = 1'b1;
  assign CLBLM_L_X68Y95_SLICE_X103Y95_A6 = 1'b1;
  assign CLBLM_L_X68Y95_SLICE_X103Y95_B1 = 1'b1;
  assign CLBLM_L_X68Y95_SLICE_X103Y95_B2 = 1'b1;
  assign CLBLM_L_X68Y95_SLICE_X103Y95_B3 = 1'b1;
  assign CLBLM_L_X68Y95_SLICE_X103Y95_B4 = 1'b1;
  assign CLBLM_L_X68Y95_SLICE_X103Y95_B5 = 1'b1;
  assign CLBLM_L_X68Y95_SLICE_X103Y95_B6 = 1'b1;
  assign CLBLM_L_X68Y95_SLICE_X103Y95_C1 = 1'b1;
  assign CLBLM_L_X68Y95_SLICE_X103Y95_C2 = 1'b1;
  assign CLBLM_L_X68Y95_SLICE_X103Y95_C3 = 1'b1;
  assign CLBLM_L_X68Y95_SLICE_X103Y95_C4 = 1'b1;
  assign CLBLM_L_X68Y95_SLICE_X103Y95_C5 = 1'b1;
  assign CLBLM_L_X68Y95_SLICE_X103Y95_C6 = 1'b1;
  assign CLBLM_L_X72Y107_SLICE_X108Y107_A1 = CLBLL_R_X71Y109_SLICE_X106Y109_CO6;
  assign CLBLM_L_X72Y107_SLICE_X108Y107_A2 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X72Y107_SLICE_X108Y107_A3 = CLBLM_L_X72Y107_SLICE_X108Y107_AQ;
  assign CLBLM_L_X72Y107_SLICE_X108Y107_A4 = CLBLM_L_X72Y108_SLICE_X109Y108_A5Q;
  assign CLBLM_L_X72Y107_SLICE_X108Y107_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y107_SLICE_X108Y107_A6 = CLBLM_L_X72Y108_SLICE_X108Y108_CQ;
  assign CLBLM_L_X68Y95_SLICE_X103Y95_D1 = 1'b1;
  assign CLBLM_L_X68Y95_SLICE_X103Y95_D2 = 1'b1;
  assign CLBLM_L_X68Y95_SLICE_X103Y95_D3 = 1'b1;
  assign CLBLM_L_X68Y95_SLICE_X103Y95_D4 = 1'b1;
  assign CLBLM_L_X68Y95_SLICE_X103Y95_D5 = 1'b1;
  assign CLBLM_L_X68Y95_SLICE_X103Y95_D6 = 1'b1;
  assign CLBLM_L_X72Y107_SLICE_X108Y107_AX = CLBLM_L_X72Y107_SLICE_X109Y107_BQ;
  assign CLBLM_L_X72Y107_SLICE_X108Y107_B1 = CLBLL_R_X71Y107_SLICE_X106Y107_C5Q;
  assign CLBLM_L_X72Y107_SLICE_X108Y107_B2 = CLBLL_R_X71Y107_SLICE_X106Y107_CQ;
  assign CLBLM_L_X72Y107_SLICE_X108Y107_B3 = CLBLM_L_X72Y107_SLICE_X108Y107_AQ;
  assign CLBLM_L_X72Y107_SLICE_X108Y107_B4 = CLBLL_R_X73Y108_SLICE_X110Y108_A5Q;
  assign CLBLM_L_X72Y107_SLICE_X108Y107_B5 = CLBLM_L_X72Y107_SLICE_X108Y107_CQ;
  assign CLBLM_L_X68Y95_SLICE_X102Y95_A1 = CLBLM_L_X60Y94_SLICE_X90Y94_CQ;
  assign CLBLM_L_X68Y95_SLICE_X102Y95_A2 = CLBLM_L_X62Y95_SLICE_X92Y95_BQ;
  assign CLBLM_L_X68Y95_SLICE_X102Y95_A3 = CLBLM_L_X68Y95_SLICE_X102Y95_AQ;
  assign CLBLM_L_X68Y95_SLICE_X102Y95_A4 = CLBLM_L_X68Y95_SLICE_X102Y95_BO6;
  assign CLBLM_L_X68Y95_SLICE_X102Y95_A5 = CLBLM_L_X60Y94_SLICE_X90Y94_BQ;
  assign CLBLM_L_X68Y95_SLICE_X102Y95_A6 = CLBLM_L_X68Y95_SLICE_X102Y95_A5Q;
  assign CLBLM_L_X72Y107_SLICE_X108Y107_C1 = CLBLL_R_X71Y107_SLICE_X106Y107_BO5;
  assign CLBLM_L_X72Y107_SLICE_X108Y107_C2 = CLBLM_L_X72Y107_SLICE_X108Y107_BO5;
  assign CLBLM_L_X72Y107_SLICE_X108Y107_C3 = CLBLM_L_X72Y107_SLICE_X109Y107_BO6;
  assign CLBLM_L_X68Y95_SLICE_X102Y95_AX = CLBLM_L_X68Y95_SLICE_X102Y95_AQ;
  assign CLBLM_L_X72Y107_SLICE_X108Y107_C4 = CLBLM_L_X72Y108_SLICE_X108Y108_DQ;
  assign CLBLM_L_X68Y95_SLICE_X102Y95_B1 = CLBLM_L_X60Y94_SLICE_X90Y94_CQ;
  assign CLBLM_L_X68Y95_SLICE_X102Y95_B2 = CLBLM_L_X62Y95_SLICE_X92Y95_BQ;
  assign CLBLM_L_X68Y95_SLICE_X102Y95_B3 = CLBLM_L_X68Y95_SLICE_X102Y95_AQ;
  assign CLBLM_L_X68Y95_SLICE_X102Y95_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y95_SLICE_X102Y95_B5 = CLBLM_L_X68Y99_SLICE_X102Y99_AQ;
  assign CLBLM_L_X68Y95_SLICE_X102Y95_B6 = CLBLM_L_X68Y95_SLICE_X102Y95_A5Q;
  assign CLBLM_L_X72Y107_SLICE_X108Y107_CX = CLBLM_L_X72Y107_SLICE_X108Y107_BQ;
  assign CLBLM_L_X72Y107_SLICE_X108Y107_D1 = CLBLM_L_X72Y106_SLICE_X108Y106_AQ;
  assign CLBLM_L_X72Y107_SLICE_X108Y107_D2 = CLBLL_R_X73Y107_SLICE_X110Y107_AQ;
  assign CLBLM_L_X72Y107_SLICE_X108Y107_D3 = CLBLM_L_X72Y107_SLICE_X108Y107_A5Q;
  assign CLBLM_L_X68Y95_SLICE_X102Y95_C1 = 1'b1;
  assign CLBLM_L_X68Y95_SLICE_X102Y95_C2 = 1'b1;
  assign CLBLM_L_X68Y95_SLICE_X102Y95_C3 = 1'b1;
  assign CLBLM_L_X68Y95_SLICE_X102Y95_C4 = 1'b1;
  assign CLBLM_L_X68Y95_SLICE_X102Y95_C5 = 1'b1;
  assign CLBLM_L_X68Y95_SLICE_X102Y95_C6 = 1'b1;
  assign CLBLM_L_X72Y107_SLICE_X108Y107_D6 = CLBLL_R_X73Y108_SLICE_X110Y108_A5Q;
  assign CLBLM_L_X72Y107_SLICE_X108Y107_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X68Y95_SLICE_X102Y95_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X74Y104_SLICE_X113Y104_D6 = 1'b1;
  assign CLBLM_L_X68Y95_SLICE_X102Y95_D1 = 1'b1;
  assign CLBLM_L_X68Y95_SLICE_X102Y95_D2 = 1'b1;
  assign CLBLM_L_X68Y95_SLICE_X102Y95_D3 = 1'b1;
  assign CLBLM_L_X68Y95_SLICE_X102Y95_D4 = 1'b1;
  assign CLBLM_L_X68Y95_SLICE_X102Y95_D5 = 1'b1;
  assign CLBLL_R_X71Y133_SLICE_X106Y133_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y133_SLICE_X106Y133_A2 = CLBLM_L_X70Y135_SLICE_X105Y135_AQ;
  assign CLBLL_R_X71Y133_SLICE_X106Y133_A3 = CLBLL_R_X71Y133_SLICE_X106Y133_AQ;
  assign CLBLL_R_X71Y133_SLICE_X106Y133_A4 = CLBLM_L_X72Y133_SLICE_X109Y133_CO6;
  assign CLBLL_R_X71Y133_SLICE_X106Y133_A5 = CLBLM_L_X70Y132_SLICE_X105Y132_AQ;
  assign CLBLL_R_X71Y133_SLICE_X106Y133_A6 = 1'b1;
  assign CLBLM_L_X68Y95_SLICE_X102Y95_D6 = 1'b1;
  assign CLBLM_L_X68Y95_SLICE_X102Y95_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X71Y133_SLICE_X106Y133_B1 = CLBLM_L_X70Y124_SLICE_X105Y124_AO6;
  assign CLBLL_R_X71Y133_SLICE_X106Y133_B2 = CLBLL_R_X71Y133_SLICE_X106Y133_BQ;
  assign CLBLL_R_X71Y133_SLICE_X106Y133_B3 = CLBLM_L_X70Y133_SLICE_X105Y133_AQ;
  assign CLBLL_R_X71Y133_SLICE_X106Y133_B4 = CLBLM_L_X70Y133_SLICE_X105Y133_DQ;
  assign CLBLL_R_X71Y133_SLICE_X106Y133_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y133_SLICE_X106Y133_B6 = CLBLM_L_X70Y133_SLICE_X104Y133_AQ;
  assign CLBLM_R_X67Y115_SLICE_X100Y115_A1 = RIOB33_X105Y53_IOB_X1Y54_I;
  assign CLBLL_R_X71Y133_SLICE_X106Y133_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y133_SLICE_X106Y133_C2 = CLBLL_R_X71Y133_SLICE_X106Y133_CQ;
  assign CLBLL_R_X71Y133_SLICE_X106Y133_C3 = CLBLM_L_X72Y133_SLICE_X108Y133_A5Q;
  assign CLBLL_R_X71Y133_SLICE_X106Y133_C4 = CLBLL_R_X71Y132_SLICE_X106Y132_CQ;
  assign CLBLL_R_X71Y133_SLICE_X106Y133_C5 = CLBLM_L_X72Y133_SLICE_X108Y133_AQ;
  assign CLBLL_R_X71Y133_SLICE_X106Y133_C6 = CLBLL_R_X73Y132_SLICE_X110Y132_BO6;
  assign CLBLM_R_X67Y115_SLICE_X100Y115_A2 = 1'b1;
  assign CLBLM_R_X67Y115_SLICE_X100Y115_A3 = CLBLM_R_X67Y115_SLICE_X100Y115_AQ;
  assign CLBLL_R_X71Y133_SLICE_X106Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X67Y115_SLICE_X100Y115_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y133_SLICE_X106Y133_D1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y133_SLICE_X106Y133_D2 = CLBLL_R_X71Y133_SLICE_X106Y133_CQ;
  assign CLBLL_R_X71Y133_SLICE_X106Y133_D3 = CLBLL_R_X71Y133_SLICE_X106Y133_DQ;
  assign CLBLL_R_X71Y133_SLICE_X106Y133_D4 = CLBLL_R_X71Y132_SLICE_X106Y132_CQ;
  assign CLBLL_R_X71Y133_SLICE_X106Y133_D5 = CLBLM_L_X72Y133_SLICE_X108Y133_BO5;
  assign CLBLL_R_X71Y133_SLICE_X106Y133_D6 = 1'b1;
  assign CLBLM_R_X67Y115_SLICE_X100Y115_A5 = RIOB33_X105Y53_IOB_X1Y53_I;
  assign CLBLM_R_X67Y115_SLICE_X100Y115_A6 = 1'b1;
  assign CLBLL_R_X71Y133_SLICE_X106Y133_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y130_SLICE_X109Y130_D5 = 1'b1;
  assign CLBLM_L_X72Y130_SLICE_X109Y130_D6 = 1'b1;
  assign CLBLL_R_X71Y133_SLICE_X107Y133_A1 = CLBLM_L_X70Y124_SLICE_X105Y124_AO6;
  assign CLBLL_R_X71Y133_SLICE_X107Y133_A2 = CLBLM_L_X70Y133_SLICE_X104Y133_AQ;
  assign CLBLL_R_X71Y133_SLICE_X107Y133_A3 = CLBLL_R_X71Y133_SLICE_X107Y133_AQ;
  assign CLBLL_R_X71Y133_SLICE_X107Y133_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y133_SLICE_X107Y133_A5 = CLBLM_L_X70Y133_SLICE_X105Y133_AQ;
  assign CLBLL_R_X71Y133_SLICE_X107Y133_A6 = CLBLL_R_X71Y134_SLICE_X107Y134_CQ;
  assign CLBLM_R_X67Y115_SLICE_X100Y115_B1 = 1'b1;
  assign CLBLM_R_X67Y115_SLICE_X100Y115_B2 = 1'b1;
  assign CLBLL_R_X71Y133_SLICE_X107Y133_B1 = 1'b1;
  assign CLBLL_R_X71Y133_SLICE_X107Y133_B2 = CLBLL_R_X71Y133_SLICE_X107Y133_BQ;
  assign CLBLL_R_X71Y133_SLICE_X107Y133_B3 = CLBLL_R_X71Y133_SLICE_X107Y133_AQ;
  assign CLBLL_R_X71Y133_SLICE_X107Y133_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y133_SLICE_X107Y133_B5 = CLBLL_R_X71Y133_SLICE_X107Y133_CO6;
  assign CLBLL_R_X71Y133_SLICE_X107Y133_B6 = CLBLL_R_X71Y134_SLICE_X107Y134_CQ;
  assign CLBLM_R_X67Y115_SLICE_X100Y115_B3 = 1'b1;
  assign CLBLM_L_X72Y130_SLICE_X109Y130_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X71Y133_SLICE_X107Y133_C1 = CLBLM_L_X70Y133_SLICE_X105Y133_AQ;
  assign CLBLL_R_X71Y133_SLICE_X107Y133_C2 = CLBLM_L_X70Y133_SLICE_X104Y133_AQ;
  assign CLBLL_R_X71Y133_SLICE_X107Y133_C3 = CLBLM_L_X70Y124_SLICE_X105Y124_AO6;
  assign CLBLL_R_X71Y133_SLICE_X107Y133_C4 = 1'b1;
  assign CLBLL_R_X71Y133_SLICE_X107Y133_C5 = 1'b1;
  assign CLBLL_R_X71Y133_SLICE_X107Y133_C6 = 1'b1;
  assign CLBLM_R_X67Y115_SLICE_X100Y115_B5 = 1'b1;
  assign CLBLM_R_X67Y115_SLICE_X100Y115_B6 = 1'b1;
  assign CLBLL_R_X71Y133_SLICE_X107Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1 = CLBLM_L_X74Y129_SLICE_X113Y129_BO6;
  assign CLBLL_R_X71Y133_SLICE_X107Y133_D1 = 1'b1;
  assign CLBLL_R_X71Y133_SLICE_X107Y133_D2 = 1'b1;
  assign CLBLL_R_X71Y133_SLICE_X107Y133_D3 = 1'b1;
  assign CLBLL_R_X71Y133_SLICE_X107Y133_D4 = 1'b1;
  assign CLBLL_R_X71Y133_SLICE_X107Y133_D5 = 1'b1;
  assign CLBLL_R_X71Y133_SLICE_X107Y133_D6 = 1'b1;
  assign CLBLM_L_X72Y130_SLICE_X108Y130_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1 = 1'b1;
  assign CLBLL_R_X71Y133_SLICE_X107Y133_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y130_SLICE_X108Y130_A2 = CLBLL_R_X71Y130_SLICE_X107Y130_AQ;
  assign CLBLM_L_X72Y130_SLICE_X108Y130_A3 = CLBLM_L_X72Y130_SLICE_X108Y130_AQ;
  assign CLBLM_L_X72Y130_SLICE_X108Y130_A4 = CLBLM_L_X72Y133_SLICE_X109Y133_DO6;
  assign CLBLM_R_X67Y115_SLICE_X100Y115_C1 = 1'b1;
  assign CLBLM_L_X72Y130_SLICE_X108Y130_A5 = CLBLM_L_X72Y131_SLICE_X108Y131_AQ;
  assign CLBLM_R_X67Y115_SLICE_X100Y115_C2 = 1'b1;
  assign RIOB33_X105Y115_IOB_X1Y115_O = CLBLM_L_X62Y100_SLICE_X92Y100_AQ;
  assign RIOB33_X105Y115_IOB_X1Y116_O = CLBLM_L_X68Y95_SLICE_X102Y95_AQ;
  assign CLBLM_L_X72Y130_SLICE_X108Y130_A6 = 1'b1;
  assign CLBLM_R_X67Y115_SLICE_X100Y115_C3 = 1'b1;
  assign CLBLM_L_X74Y104_SLICE_X112Y104_C2 = CLBLM_L_X74Y104_SLICE_X112Y104_CQ;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_B5 = 1'b1;
  assign CLBLM_R_X67Y115_SLICE_X100Y115_C4 = 1'b1;
  assign CLBLM_L_X74Y104_SLICE_X112Y104_C3 = CLBLL_R_X73Y104_SLICE_X110Y104_DO5;
  assign CLBLM_R_X67Y115_SLICE_X100Y115_C5 = 1'b1;
  assign CLBLM_L_X74Y104_SLICE_X112Y104_C4 = CLBLM_L_X74Y104_SLICE_X112Y104_BQ;
  assign CLBLM_R_X67Y115_SLICE_X100Y115_C6 = 1'b1;
  assign CLBLM_L_X74Y104_SLICE_X112Y104_C5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y104_SLICE_X112Y104_C6 = CLBLM_L_X72Y103_SLICE_X108Y103_DO6;
  assign CLBLM_L_X72Y130_SLICE_X108Y130_B1 = CLBLM_L_X72Y129_SLICE_X108Y129_AQ;
  assign CLBLM_L_X72Y130_SLICE_X108Y130_B2 = CLBLM_L_X72Y130_SLICE_X108Y130_BQ;
  assign CLBLM_R_X67Y115_SLICE_X100Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X72Y130_SLICE_X108Y130_B3 = CLBLL_R_X71Y130_SLICE_X106Y130_BQ;
  assign CLBLM_L_X74Y104_SLICE_X112Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X72Y130_SLICE_X108Y130_B4 = CLBLM_L_X72Y129_SLICE_X108Y129_BQ;
  assign CLBLM_L_X72Y130_SLICE_X108Y130_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y130_SLICE_X108Y130_B6 = CLBLL_R_X71Y125_SLICE_X107Y125_BO6;
  assign CLBLM_L_X72Y108_SLICE_X109Y108_A1 = 1'b1;
  assign CLBLM_L_X72Y108_SLICE_X109Y108_A2 = CLBLM_L_X72Y108_SLICE_X109Y108_A5Q;
  assign CLBLM_L_X72Y108_SLICE_X109Y108_A3 = CLBLM_L_X72Y108_SLICE_X109Y108_AQ;
  assign CLBLM_L_X72Y108_SLICE_X109Y108_A4 = CLBLL_R_X71Y111_SLICE_X106Y111_AQ;
  assign CLBLM_L_X72Y108_SLICE_X109Y108_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y108_SLICE_X109Y108_A6 = 1'b1;
  assign CLBLM_R_X67Y115_SLICE_X100Y115_D1 = 1'b1;
  assign CLBLM_L_X72Y108_SLICE_X109Y108_B1 = 1'b1;
  assign CLBLM_L_X72Y108_SLICE_X109Y108_B2 = 1'b1;
  assign CLBLM_L_X72Y108_SLICE_X109Y108_B3 = CLBLM_L_X72Y108_SLICE_X109Y108_AQ;
  assign CLBLM_L_X72Y108_SLICE_X109Y108_B4 = 1'b1;
  assign CLBLM_L_X72Y108_SLICE_X109Y108_B5 = CLBLL_R_X71Y111_SLICE_X106Y111_AQ;
  assign CLBLM_L_X72Y108_SLICE_X109Y108_B6 = 1'b1;
  assign CLBLM_L_X74Y104_SLICE_X112Y104_D1 = 1'b1;
  assign CLBLM_L_X74Y104_SLICE_X112Y104_D2 = 1'b1;
  assign CLBLM_L_X72Y108_SLICE_X109Y108_C1 = 1'b1;
  assign CLBLM_L_X72Y108_SLICE_X109Y108_C2 = CLBLM_L_X72Y108_SLICE_X109Y108_AQ;
  assign CLBLM_L_X72Y108_SLICE_X109Y108_C3 = CLBLL_R_X71Y111_SLICE_X106Y111_AQ;
  assign CLBLM_L_X72Y108_SLICE_X109Y108_C4 = CLBLM_L_X72Y108_SLICE_X109Y108_A5Q;
  assign CLBLM_L_X68Y96_SLICE_X103Y96_A1 = CLBLM_L_X68Y98_SLICE_X103Y98_A5Q;
  assign CLBLM_L_X68Y96_SLICE_X103Y96_A2 = CLBLM_L_X68Y95_SLICE_X102Y95_AQ;
  assign CLBLM_L_X68Y96_SLICE_X103Y96_A3 = CLBLM_L_X68Y98_SLICE_X102Y98_DQ;
  assign CLBLM_L_X68Y96_SLICE_X103Y96_A4 = CLBLM_L_X60Y94_SLICE_X90Y94_BQ;
  assign CLBLM_L_X68Y96_SLICE_X103Y96_A5 = CLBLM_L_X68Y99_SLICE_X103Y99_CQ;
  assign CLBLM_L_X68Y96_SLICE_X103Y96_A6 = CLBLM_L_X68Y99_SLICE_X103Y99_C5Q;
  assign CLBLM_L_X72Y108_SLICE_X109Y108_C5 = 1'b1;
  assign CLBLM_L_X72Y108_SLICE_X109Y108_C6 = 1'b1;
  assign CLBLM_L_X72Y108_SLICE_X109Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X68Y96_SLICE_X103Y96_B1 = CLBLM_L_X68Y95_SLICE_X102Y95_A5Q;
  assign CLBLM_L_X68Y96_SLICE_X103Y96_B2 = CLBLM_L_X68Y95_SLICE_X102Y95_AQ;
  assign CLBLM_L_X68Y96_SLICE_X103Y96_B3 = 1'b1;
  assign CLBLM_L_X68Y96_SLICE_X103Y96_B4 = CLBLM_L_X62Y95_SLICE_X92Y95_BQ;
  assign CLBLM_L_X68Y96_SLICE_X103Y96_B5 = CLBLM_L_X60Y94_SLICE_X90Y94_BQ;
  assign CLBLM_L_X68Y96_SLICE_X103Y96_B6 = 1'b1;
  assign CLBLM_L_X72Y108_SLICE_X109Y108_D1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y108_SLICE_X109Y108_D2 = CLBLL_R_X73Y108_SLICE_X110Y108_BQ;
  assign CLBLM_L_X68Y96_SLICE_X103Y96_C1 = 1'b1;
  assign CLBLM_L_X68Y96_SLICE_X103Y96_C2 = 1'b1;
  assign CLBLM_L_X68Y96_SLICE_X103Y96_C3 = 1'b1;
  assign CLBLM_L_X68Y96_SLICE_X103Y96_C4 = 1'b1;
  assign CLBLM_L_X68Y96_SLICE_X103Y96_C5 = 1'b1;
  assign CLBLM_L_X68Y96_SLICE_X103Y96_C6 = 1'b1;
  assign CLBLM_L_X72Y108_SLICE_X108Y108_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y108_SLICE_X108Y108_A2 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X72Y108_SLICE_X108Y108_A3 = CLBLM_L_X72Y108_SLICE_X109Y108_CO5;
  assign CLBLM_L_X72Y108_SLICE_X108Y108_A4 = CLBLM_L_X72Y108_SLICE_X108Y108_AQ;
  assign CLBLM_L_X72Y108_SLICE_X108Y108_A5 = CLBLL_R_X71Y109_SLICE_X106Y109_BQ;
  assign CLBLM_L_X72Y108_SLICE_X108Y108_A6 = CLBLL_R_X71Y109_SLICE_X106Y109_B5Q;
  assign CLBLM_L_X68Y96_SLICE_X103Y96_D1 = 1'b1;
  assign CLBLM_L_X68Y96_SLICE_X103Y96_D2 = 1'b1;
  assign CLBLM_L_X68Y96_SLICE_X103Y96_D3 = 1'b1;
  assign CLBLM_L_X68Y96_SLICE_X103Y96_D4 = 1'b1;
  assign CLBLM_L_X68Y96_SLICE_X103Y96_D5 = 1'b1;
  assign CLBLM_L_X68Y96_SLICE_X103Y96_D6 = 1'b1;
  assign CLBLM_L_X72Y108_SLICE_X108Y108_B1 = CLBLL_R_X71Y109_SLICE_X106Y109_B5Q;
  assign CLBLM_L_X72Y108_SLICE_X108Y108_B2 = 1'b1;
  assign CLBLM_L_X72Y108_SLICE_X108Y108_B3 = CLBLL_R_X71Y109_SLICE_X106Y109_BQ;
  assign CLBLM_L_X72Y108_SLICE_X108Y108_B4 = 1'b1;
  assign CLBLM_L_X72Y108_SLICE_X108Y108_B5 = 1'b1;
  assign CLBLM_L_X72Y108_SLICE_X108Y108_B6 = 1'b1;
  assign CLBLM_L_X68Y96_SLICE_X102Y96_A1 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X68Y96_SLICE_X102Y96_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y96_SLICE_X102Y96_A3 = CLBLM_L_X68Y96_SLICE_X102Y96_AQ;
  assign CLBLM_L_X68Y96_SLICE_X102Y96_A4 = CLBLM_L_X68Y98_SLICE_X102Y98_CQ;
  assign CLBLM_L_X68Y96_SLICE_X102Y96_A5 = CLBLM_R_X67Y98_SLICE_X101Y98_BO6;
  assign CLBLM_L_X68Y96_SLICE_X102Y96_A6 = CLBLM_R_X67Y98_SLICE_X100Y98_CO6;
  assign CLBLM_L_X72Y108_SLICE_X108Y108_C1 = CLBLM_L_X72Y108_SLICE_X109Y108_CO6;
  assign CLBLM_L_X72Y108_SLICE_X108Y108_C2 = CLBLM_L_X72Y108_SLICE_X108Y108_CQ;
  assign CLBLM_L_X72Y108_SLICE_X108Y108_C3 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X72Y108_SLICE_X108Y108_C4 = CLBLL_R_X71Y107_SLICE_X107Y107_BQ;
  assign CLBLM_L_X68Y96_SLICE_X102Y96_B1 = CLBLM_L_X68Y98_SLICE_X103Y98_A5Q;
  assign CLBLM_L_X68Y96_SLICE_X102Y96_B2 = CLBLM_L_X60Y94_SLICE_X90Y94_BQ;
  assign CLBLM_L_X68Y96_SLICE_X102Y96_B3 = CLBLM_L_X68Y99_SLICE_X103Y99_CQ;
  assign CLBLM_L_X68Y96_SLICE_X102Y96_B4 = CLBLM_L_X68Y99_SLICE_X103Y99_C5Q;
  assign CLBLM_L_X68Y96_SLICE_X102Y96_B5 = CLBLM_R_X67Y96_SLICE_X101Y96_CQ;
  assign CLBLM_L_X68Y96_SLICE_X102Y96_B6 = CLBLM_L_X68Y95_SLICE_X102Y95_AQ;
  assign CLBLM_L_X72Y108_SLICE_X108Y108_D1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y108_SLICE_X108Y108_D2 = CLBLL_R_X71Y109_SLICE_X106Y109_CO5;
  assign CLBLM_L_X72Y108_SLICE_X108Y108_D3 = CLBLM_L_X72Y108_SLICE_X108Y108_DQ;
  assign CLBLM_L_X68Y96_SLICE_X102Y96_C1 = CLBLM_L_X62Y95_SLICE_X92Y95_BQ;
  assign CLBLM_L_X68Y96_SLICE_X102Y96_C2 = CLBLM_R_X67Y97_SLICE_X100Y97_AQ;
  assign CLBLM_L_X68Y96_SLICE_X102Y96_C3 = CLBLM_R_X67Y98_SLICE_X101Y98_DQ;
  assign CLBLM_L_X68Y96_SLICE_X102Y96_C4 = CLBLM_L_X68Y95_SLICE_X102Y95_A5Q;
  assign CLBLM_L_X68Y96_SLICE_X102Y96_C5 = CLBLM_L_X68Y99_SLICE_X103Y99_CQ;
  assign CLBLM_L_X68Y96_SLICE_X102Y96_C6 = CLBLM_L_X68Y99_SLICE_X103Y99_C5Q;
  assign CLBLM_L_X72Y108_SLICE_X108Y108_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X68Y96_SLICE_X102Y96_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLL_R_X71Y134_SLICE_X106Y134_A1 = CLBLM_L_X70Y136_SLICE_X105Y136_BO5;
  assign CLBLL_R_X71Y134_SLICE_X106Y134_A2 = CLBLL_R_X75Y134_SLICE_X114Y134_CO6;
  assign CLBLL_R_X71Y134_SLICE_X106Y134_A3 = CLBLL_R_X71Y134_SLICE_X106Y134_AQ;
  assign CLBLL_R_X71Y134_SLICE_X106Y134_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y134_SLICE_X106Y134_A5 = CLBLM_L_X60Y92_SLICE_X90Y92_AQ;
  assign CLBLL_R_X71Y134_SLICE_X106Y134_A6 = CLBLM_L_X60Y94_SLICE_X90Y94_AQ;
  assign CLBLM_L_X68Y96_SLICE_X102Y96_D1 = CLBLM_L_X68Y96_SLICE_X102Y96_CO6;
  assign CLBLM_L_X68Y96_SLICE_X102Y96_D2 = CLBLM_L_X68Y96_SLICE_X103Y96_AO6;
  assign CLBLM_L_X68Y96_SLICE_X102Y96_D3 = CLBLM_L_X68Y96_SLICE_X102Y96_AQ;
  assign CLBLL_R_X71Y134_SLICE_X106Y134_B1 = CLBLM_L_X70Y135_SLICE_X105Y135_A5Q;
  assign CLBLL_R_X71Y134_SLICE_X106Y134_B2 = CLBLL_R_X71Y134_SLICE_X106Y134_BQ;
  assign CLBLL_R_X71Y134_SLICE_X106Y134_B3 = CLBLM_L_X72Y133_SLICE_X109Y133_CO6;
  assign CLBLL_R_X71Y134_SLICE_X106Y134_B4 = CLBLM_L_X72Y134_SLICE_X109Y134_BO6;
  assign CLBLL_R_X71Y134_SLICE_X106Y134_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y134_SLICE_X106Y134_B6 = CLBLM_L_X70Y135_SLICE_X105Y135_AQ;
  assign CLBLM_L_X68Y96_SLICE_X102Y96_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_B3 = 1'b1;
  assign CLBLL_R_X71Y134_SLICE_X106Y134_C1 = 1'b1;
  assign CLBLL_R_X71Y134_SLICE_X106Y134_C2 = 1'b1;
  assign CLBLL_R_X71Y134_SLICE_X106Y134_C3 = 1'b1;
  assign CLBLL_R_X71Y134_SLICE_X106Y134_C4 = 1'b1;
  assign CLBLL_R_X71Y134_SLICE_X106Y134_C5 = 1'b1;
  assign CLBLL_R_X71Y134_SLICE_X106Y134_C6 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_B4 = 1'b1;
  assign CLBLL_R_X71Y134_SLICE_X106Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X76Y111_SLICE_X117Y111_D1 = 1'b1;
  assign RIOI3_X105Y77_OLOGIC_X1Y77_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1 = 1'b1;
  assign CLBLM_L_X76Y111_SLICE_X117Y111_D2 = 1'b1;
  assign CLBLL_R_X71Y134_SLICE_X106Y134_D1 = 1'b1;
  assign CLBLL_R_X71Y134_SLICE_X106Y134_D2 = 1'b1;
  assign CLBLL_R_X71Y134_SLICE_X106Y134_D3 = 1'b1;
  assign CLBLL_R_X71Y134_SLICE_X106Y134_D4 = 1'b1;
  assign CLBLL_R_X71Y134_SLICE_X106Y134_D5 = 1'b1;
  assign CLBLL_R_X71Y134_SLICE_X106Y134_D6 = 1'b1;
  assign CLBLM_L_X76Y111_SLICE_X117Y111_D3 = 1'b1;
  assign CLBLL_R_X71Y134_SLICE_X106Y134_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X76Y111_SLICE_X117Y111_D4 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1 = CLBLL_R_X75Y133_SLICE_X114Y133_BQ;
  assign CLBLM_L_X76Y111_SLICE_X117Y111_D5 = 1'b1;
  assign CLBLM_L_X76Y111_SLICE_X117Y111_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_C2 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_C3 = 1'b1;
  assign CLBLL_R_X71Y134_SLICE_X107Y134_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y134_SLICE_X107Y134_A2 = CLBLM_L_X70Y135_SLICE_X105Y135_AQ;
  assign CLBLL_R_X71Y134_SLICE_X107Y134_A3 = CLBLL_R_X71Y134_SLICE_X107Y134_AQ;
  assign CLBLL_R_X71Y134_SLICE_X107Y134_A4 = CLBLL_R_X71Y133_SLICE_X106Y133_BQ;
  assign CLBLL_R_X71Y134_SLICE_X107Y134_A5 = CLBLM_L_X72Y133_SLICE_X109Y133_CO6;
  assign CLBLL_R_X71Y134_SLICE_X107Y134_A6 = CLBLM_L_X70Y135_SLICE_X105Y135_A5Q;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_C6 = 1'b1;
  assign CLBLL_R_X71Y134_SLICE_X107Y134_B1 = 1'b1;
  assign CLBLL_R_X71Y134_SLICE_X107Y134_B2 = CLBLL_R_X71Y134_SLICE_X107Y134_BQ;
  assign CLBLL_R_X71Y134_SLICE_X107Y134_B3 = CLBLL_R_X71Y134_SLICE_X107Y134_AQ;
  assign CLBLL_R_X71Y134_SLICE_X107Y134_B4 = CLBLL_R_X71Y133_SLICE_X106Y133_BQ;
  assign CLBLL_R_X71Y134_SLICE_X107Y134_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y134_SLICE_X107Y134_B6 = CLBLM_L_X70Y134_SLICE_X105Y134_DO6;
  assign CLBLL_R_X71Y134_SLICE_X107Y134_C1 = CLBLM_L_X72Y133_SLICE_X109Y133_CO6;
  assign CLBLL_R_X71Y134_SLICE_X107Y134_C2 = CLBLL_R_X71Y134_SLICE_X107Y134_CQ;
  assign CLBLL_R_X71Y134_SLICE_X107Y134_C3 = CLBLM_L_X70Y135_SLICE_X105Y135_A5Q;
  assign CLBLL_R_X71Y134_SLICE_X107Y134_C4 = CLBLL_R_X71Y134_SLICE_X107Y134_BQ;
  assign CLBLL_R_X71Y134_SLICE_X107Y134_C5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X71Y134_SLICE_X107Y134_C6 = CLBLM_L_X70Y135_SLICE_X105Y135_AQ;
  assign CLBLM_L_X76Y111_SLICE_X116Y111_A1 = 1'b1;
  assign CLBLL_R_X71Y134_SLICE_X107Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_C4 = 1'b1;
  assign CLBLM_L_X76Y111_SLICE_X116Y111_A2 = 1'b1;
  assign CLBLL_R_X71Y134_SLICE_X107Y134_D1 = 1'b1;
  assign CLBLL_R_X71Y134_SLICE_X107Y134_D2 = 1'b1;
  assign CLBLL_R_X71Y134_SLICE_X107Y134_D3 = 1'b1;
  assign CLBLL_R_X71Y134_SLICE_X107Y134_D4 = 1'b1;
  assign CLBLL_R_X71Y134_SLICE_X107Y134_D5 = 1'b1;
  assign CLBLL_R_X71Y134_SLICE_X107Y134_D6 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_C5 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_A1 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_A2 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_A3 = CLBLL_R_X71Y124_SLICE_X106Y124_A5Q;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_A4 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_A5 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_A6 = 1'b1;
  assign CLBLL_R_X71Y134_SLICE_X107Y134_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X76Y111_SLICE_X116Y111_A5 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_B1 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_B2 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_B3 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_B4 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_B5 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_B6 = 1'b1;
  assign CLBLM_L_X76Y111_SLICE_X116Y111_A6 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_C1 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_C2 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_C3 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_C4 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_C5 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_C6 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_A6 = 1'b1;
  assign CLBLM_L_X76Y111_SLICE_X116Y111_AX = CLBLM_R_X65Y111_SLICE_X98Y111_AQ;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_D1 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_D2 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_D3 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_D4 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_D5 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_D6 = 1'b1;
  assign CLBLM_L_X76Y111_SLICE_X116Y111_B1 = 1'b1;
  assign CLBLM_L_X76Y111_SLICE_X116Y111_B2 = 1'b1;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X76Y111_SLICE_X116Y111_B3 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_D1 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_B2 = CLBLM_L_X64Y99_SLICE_X96Y99_A5Q;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1 = 1'b1;
  assign CLBLM_L_X76Y111_SLICE_X116Y111_B4 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_D2 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_B3 = CLBLM_R_X65Y101_SLICE_X99Y101_AQ;
  assign CLBLM_L_X76Y111_SLICE_X116Y111_B5 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_D3 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_B4 = CLBLM_L_X64Y99_SLICE_X96Y99_BQ;
  assign CLBLM_L_X76Y111_SLICE_X116Y111_B6 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_D4 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_D5 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_A1 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_A2 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_A3 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_A4 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_A5 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_A6 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_D6 = 1'b1;
  assign RIOI3_X105Y77_ILOGIC_X1Y78_D = RIOB33_X105Y77_IOB_X1Y78_I;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_B1 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_B2 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_B3 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_B4 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_B5 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_B6 = 1'b1;
  assign CLBLM_L_X76Y111_SLICE_X116Y111_BX = CLBLM_L_X62Y99_SLICE_X93Y99_AQ;
  assign CLBLM_L_X78Y130_SLICE_X121Y130_A1 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_C1 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_C2 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_C3 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_C4 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_C5 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_C6 = 1'b1;
  assign CLBLM_L_X72Y109_SLICE_X109Y109_A1 = RIOB33_X105Y57_IOB_X1Y57_I;
  assign CLBLM_L_X72Y109_SLICE_X109Y109_A2 = CLBLM_L_X72Y111_SLICE_X109Y111_BQ;
  assign CLBLM_L_X72Y109_SLICE_X109Y109_A3 = 1'b1;
  assign CLBLM_L_X72Y109_SLICE_X109Y109_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y109_SLICE_X109Y109_A5 = CLBLM_L_X72Y109_SLICE_X108Y109_AQ;
  assign CLBLM_L_X72Y109_SLICE_X109Y109_A6 = 1'b1;
  assign CLBLM_L_X72Y109_SLICE_X109Y109_B1 = CLBLM_L_X72Y109_SLICE_X109Y109_AQ;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_D1 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_D2 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_D3 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_D4 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_D5 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_D6 = 1'b1;
  assign CLBLM_L_X72Y109_SLICE_X109Y109_B2 = CLBLM_L_X72Y109_SLICE_X109Y109_A5Q;
  assign CLBLM_L_X72Y109_SLICE_X109Y109_B3 = RIOB33_X105Y57_IOB_X1Y58_I;
  assign CLBLM_L_X72Y109_SLICE_X109Y109_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y109_SLICE_X109Y109_B5 = 1'b1;
  assign CLBLM_L_X72Y109_SLICE_X109Y109_B6 = 1'b1;
  assign CLBLM_L_X68Y97_SLICE_X103Y97_A1 = CLBLM_R_X67Y96_SLICE_X101Y96_DQ;
  assign CLBLM_L_X68Y97_SLICE_X103Y97_A2 = CLBLM_L_X62Y95_SLICE_X92Y95_CQ;
  assign CLBLM_L_X68Y97_SLICE_X103Y97_A3 = CLBLM_L_X68Y99_SLICE_X103Y99_CQ;
  assign CLBLM_L_X68Y97_SLICE_X103Y97_A4 = CLBLM_L_X68Y99_SLICE_X103Y99_C5Q;
  assign CLBLM_L_X68Y97_SLICE_X103Y97_A5 = CLBLM_R_X67Y96_SLICE_X101Y96_AQ;
  assign CLBLM_L_X68Y97_SLICE_X103Y97_A6 = CLBLM_L_X60Y94_SLICE_X90Y94_CQ;
  assign CLBLM_L_X72Y109_SLICE_X109Y109_C2 = RIOB33_X105Y59_IOB_X1Y59_I;
  assign CLBLM_L_X72Y109_SLICE_X109Y109_C3 = 1'b1;
  assign CLBLM_L_X68Y97_SLICE_X103Y97_AX = CLBLM_L_X68Y99_SLICE_X102Y99_AQ;
  assign CLBLM_L_X72Y109_SLICE_X109Y109_C5 = CLBLM_L_X72Y109_SLICE_X109Y109_B5Q;
  assign CLBLM_L_X68Y97_SLICE_X103Y97_B1 = CLBLM_L_X68Y99_SLICE_X103Y99_CQ;
  assign CLBLM_L_X68Y97_SLICE_X103Y97_B2 = CLBLM_R_X67Y96_SLICE_X101Y96_BQ;
  assign CLBLM_L_X68Y97_SLICE_X103Y97_B3 = CLBLM_L_X68Y99_SLICE_X103Y99_C5Q;
  assign CLBLM_L_X68Y97_SLICE_X103Y97_B4 = CLBLM_L_X68Y99_SLICE_X102Y99_AQ;
  assign CLBLM_L_X68Y97_SLICE_X103Y97_B5 = CLBLM_L_X68Y97_SLICE_X102Y97_AQ;
  assign CLBLM_L_X68Y97_SLICE_X103Y97_B6 = CLBLM_R_X67Y97_SLICE_X101Y97_AQ;
  assign CLBLM_L_X72Y109_SLICE_X109Y109_D3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y109_SLICE_X109Y109_D4 = CLBLM_L_X72Y109_SLICE_X109Y109_BQ;
  assign CLBLM_L_X72Y109_SLICE_X109Y109_D5 = CLBLM_L_X72Y109_SLICE_X109Y109_AQ;
  assign CLBLM_L_X68Y97_SLICE_X103Y97_C1 = CLBLM_L_X68Y97_SLICE_X103Y97_AO6;
  assign CLBLM_L_X68Y97_SLICE_X103Y97_C2 = CLBLM_L_X68Y98_SLICE_X103Y98_DO6;
  assign CLBLM_L_X68Y97_SLICE_X103Y97_C3 = CLBLM_L_X68Y97_SLICE_X102Y97_BO6;
  assign CLBLM_L_X68Y97_SLICE_X103Y97_C4 = CLBLM_L_X68Y97_SLICE_X102Y97_AO6;
  assign CLBLM_L_X68Y97_SLICE_X103Y97_C5 = CLBLM_L_X68Y97_SLICE_X103Y97_DO6;
  assign CLBLM_L_X68Y97_SLICE_X103Y97_C6 = CLBLM_L_X68Y97_SLICE_X103Y97_BO6;
  assign CLBLM_L_X72Y109_SLICE_X108Y109_A1 = CLBLM_L_X72Y109_SLICE_X109Y109_BQ;
  assign CLBLM_L_X72Y109_SLICE_X108Y109_A2 = CLBLM_L_X72Y111_SLICE_X108Y111_CQ;
  assign CLBLM_L_X68Y97_SLICE_X103Y97_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X72Y109_SLICE_X108Y109_A3 = 1'b1;
  assign CLBLM_L_X72Y109_SLICE_X108Y109_A4 = CLBLM_L_X72Y111_SLICE_X109Y111_BQ;
  assign CLBLM_L_X72Y109_SLICE_X108Y109_A5 = CLBLM_L_X72Y109_SLICE_X109Y109_AQ;
  assign CLBLM_L_X72Y109_SLICE_X108Y109_A6 = CLBLM_L_X72Y109_SLICE_X109Y109_CQ;
  assign CLBLM_L_X72Y109_SLICE_X108Y109_AX = CLBLM_L_X70Y109_SLICE_X105Y109_AQ;
  assign CLBLM_L_X68Y97_SLICE_X103Y97_D1 = CLBLM_L_X68Y99_SLICE_X103Y99_C5Q;
  assign CLBLM_L_X68Y97_SLICE_X103Y97_D2 = CLBLM_L_X62Y95_SLICE_X92Y95_CQ;
  assign CLBLM_L_X68Y97_SLICE_X103Y97_D3 = CLBLM_L_X68Y98_SLICE_X103Y98_A5Q;
  assign CLBLM_L_X68Y97_SLICE_X103Y97_D4 = CLBLM_L_X68Y99_SLICE_X103Y99_CQ;
  assign CLBLM_L_X68Y97_SLICE_X103Y97_D5 = 1'b1;
  assign CLBLM_L_X68Y97_SLICE_X103Y97_D6 = CLBLM_L_X68Y99_SLICE_X103Y99_BQ;
  assign CLBLM_L_X72Y109_SLICE_X108Y109_B1 = 1'b1;
  assign CLBLM_L_X72Y109_SLICE_X108Y109_B2 = 1'b1;
  assign CLBLM_L_X68Y97_SLICE_X103Y97_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y109_SLICE_X108Y109_B3 = CLBLL_R_X71Y109_SLICE_X106Y109_BQ;
  assign CLBLM_L_X72Y109_SLICE_X108Y109_B4 = 1'b1;
  assign CLBLM_L_X72Y109_SLICE_X108Y109_B5 = 1'b1;
  assign CLBLM_L_X68Y97_SLICE_X102Y97_A1 = CLBLM_L_X68Y98_SLICE_X103Y98_A5Q;
  assign CLBLM_L_X68Y97_SLICE_X102Y97_A2 = CLBLM_L_X60Y97_SLICE_X90Y97_DQ;
  assign CLBLM_L_X68Y97_SLICE_X102Y97_A3 = CLBLM_L_X68Y99_SLICE_X103Y99_C5Q;
  assign CLBLM_L_X68Y97_SLICE_X102Y97_A4 = CLBLM_R_X67Y97_SLICE_X101Y97_DQ;
  assign CLBLM_L_X68Y97_SLICE_X102Y97_A5 = CLBLM_L_X68Y99_SLICE_X103Y99_CQ;
  assign CLBLM_L_X68Y97_SLICE_X102Y97_A6 = 1'b1;
  assign CLBLM_L_X72Y109_SLICE_X108Y109_C1 = 1'b1;
  assign CLBLM_L_X72Y109_SLICE_X108Y109_C2 = 1'b1;
  assign CLBLM_L_X72Y109_SLICE_X108Y109_C3 = 1'b1;
  assign CLBLM_L_X68Y97_SLICE_X102Y97_AX = CLBLM_L_X62Y95_SLICE_X92Y95_CQ;
  assign CLBLM_L_X72Y109_SLICE_X108Y109_C4 = 1'b1;
  assign CLBLM_L_X68Y97_SLICE_X102Y97_B1 = CLBLM_R_X67Y97_SLICE_X101Y97_CQ;
  assign CLBLM_L_X68Y97_SLICE_X102Y97_B2 = CLBLM_L_X68Y95_SLICE_X102Y95_AQ;
  assign CLBLM_L_X68Y97_SLICE_X102Y97_B3 = CLBLM_R_X67Y97_SLICE_X101Y97_BQ;
  assign CLBLM_L_X68Y97_SLICE_X102Y97_B4 = CLBLM_L_X68Y99_SLICE_X103Y99_C5Q;
  assign CLBLM_L_X68Y97_SLICE_X102Y97_B5 = CLBLM_L_X68Y99_SLICE_X103Y99_CQ;
  assign CLBLM_L_X68Y97_SLICE_X102Y97_B6 = CLBLM_L_X68Y97_SLICE_X103Y97_AQ;
  assign CLBLM_L_X72Y109_SLICE_X108Y109_D1 = 1'b1;
  assign CLBLM_L_X72Y109_SLICE_X108Y109_D2 = 1'b1;
  assign CLBLM_L_X72Y109_SLICE_X108Y109_D3 = 1'b1;
  assign CLBLM_L_X68Y97_SLICE_X102Y97_C1 = CLBLM_L_X70Y106_SLICE_X104Y106_CO6;
  assign CLBLM_L_X68Y97_SLICE_X102Y97_C2 = CLBLM_L_X68Y97_SLICE_X103Y97_CO6;
  assign CLBLM_L_X68Y97_SLICE_X102Y97_C3 = CLBLM_L_X68Y99_SLICE_X102Y99_CO6;
  assign CLBLM_L_X68Y97_SLICE_X102Y97_C4 = CLBLM_L_X68Y97_SLICE_X102Y97_AO5;
  assign CLBLM_L_X68Y97_SLICE_X102Y97_C5 = CLBLM_L_X68Y97_SLICE_X102Y97_DO6;
  assign CLBLM_L_X68Y97_SLICE_X102Y97_C6 = CLBLM_L_X68Y96_SLICE_X102Y96_DO6;
  assign CLBLM_L_X72Y109_SLICE_X108Y109_D6 = 1'b1;
  assign CLBLM_L_X72Y109_SLICE_X108Y109_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X68Y97_SLICE_X102Y97_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_B5 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_B6 = CLBLM_L_X74Y127_SLICE_X112Y127_BQ;
  assign CLBLM_L_X76Y111_SLICE_X116Y111_D5 = 1'b1;
  assign CLBLM_L_X76Y111_SLICE_X116Y111_D6 = 1'b1;
  assign CLBLM_L_X68Y97_SLICE_X102Y97_D1 = CLBLM_L_X68Y95_SLICE_X102Y95_A5Q;
  assign CLBLM_L_X68Y97_SLICE_X102Y97_D2 = CLBLM_L_X68Y98_SLICE_X103Y98_CQ;
  assign CLBLM_L_X68Y97_SLICE_X102Y97_D3 = CLBLM_L_X60Y97_SLICE_X90Y97_DQ;
  assign CLBLM_L_X68Y97_SLICE_X102Y97_D4 = CLBLM_L_X68Y95_SLICE_X102Y95_AQ;
  assign CLBLM_L_X68Y97_SLICE_X102Y97_D5 = CLBLM_L_X68Y98_SLICE_X103Y98_A5Q;
  assign CLBLM_L_X68Y97_SLICE_X102Y97_D6 = CLBLM_L_X68Y98_SLICE_X102Y98_CQ;
  assign CLBLM_L_X68Y97_SLICE_X102Y97_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X76Y111_SLICE_X116Y111_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_C1 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_C2 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_C3 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_C4 = 1'b1;
  assign LIOI3_X0Y95_OLOGIC_X0Y96_D1 = CLBLM_R_X63Y97_SLICE_X95Y97_AQ;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_C5 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_C6 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_CE = CLBLM_L_X76Y109_SLICE_X116Y109_AO6;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X78Y130_SLICE_X121Y130_D4 = 1'b1;
  assign CLBLM_L_X78Y130_SLICE_X121Y130_D5 = 1'b1;
  assign RIOB33_X105Y119_IOB_X1Y119_O = CLBLM_L_X76Y128_SLICE_X116Y128_CQ;
  assign RIOB33_X105Y119_IOB_X1Y120_O = CLBLM_L_X62Y106_SLICE_X93Y106_AQ;
  assign CLBLM_L_X78Y130_SLICE_X121Y130_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_T1 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_D1 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_D2 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_D3 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_D4 = 1'b1;
  assign CLBLM_L_X78Y130_SLICE_X120Y130_A1 = CLBLM_L_X78Y130_SLICE_X120Y130_DO6;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_D5 = 1'b1;
  assign CLBLM_L_X78Y130_SLICE_X120Y130_A2 = CLBLL_R_X77Y130_SLICE_X119Y130_AQ;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_D4 = CLBLM_R_X65Y103_SLICE_X98Y103_A5Q;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_D6 = 1'b1;
  assign CLBLM_L_X78Y130_SLICE_X120Y130_A3 = CLBLM_L_X78Y130_SLICE_X120Y130_AQ;
  assign CLBLM_L_X78Y130_SLICE_X120Y130_A4 = CLBLL_R_X77Y130_SLICE_X118Y130_AQ;
  assign CLBLM_L_X78Y130_SLICE_X120Y130_A5 = CLBLL_R_X77Y128_SLICE_X118Y128_AQ;
  assign CLBLM_L_X78Y130_SLICE_X120Y130_A6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_D5 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X78Y130_SLICE_X120Y130_B1 = CLBLM_L_X78Y130_SLICE_X120Y130_DO6;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_D6 = CLBLM_L_X64Y103_SLICE_X96Y103_AQ;
  assign CLBLM_L_X78Y130_SLICE_X120Y130_B2 = CLBLM_L_X78Y130_SLICE_X120Y130_BQ;
  assign CLBLM_L_X78Y130_SLICE_X120Y130_B3 = CLBLM_L_X78Y130_SLICE_X120Y130_AQ;
  assign CLBLM_L_X78Y130_SLICE_X120Y130_B4 = CLBLL_R_X77Y130_SLICE_X119Y130_AQ;
  assign CLBLM_L_X78Y130_SLICE_X120Y130_B5 = CLBLL_R_X77Y128_SLICE_X118Y128_AQ;
  assign CLBLM_L_X72Y109_SLICE_X109Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X78Y130_SLICE_X120Y130_B6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign LIOB33_X0Y57_IOB_X0Y58_O = CLBLM_L_X72Y107_SLICE_X108Y107_BQ;
  assign LIOB33_X0Y57_IOB_X0Y57_O = CLBLM_L_X62Y95_SLICE_X92Y95_AQ;
  assign CLBLM_L_X68Y98_SLICE_X103Y98_A1 = CLBLM_L_X68Y98_SLICE_X103Y98_A5Q;
  assign CLBLM_L_X68Y98_SLICE_X103Y98_A2 = CLBLM_L_X68Y96_SLICE_X103Y96_BO6;
  assign CLBLM_L_X68Y98_SLICE_X103Y98_A3 = CLBLM_L_X68Y97_SLICE_X102Y97_AQ;
  assign CLBLM_L_X68Y98_SLICE_X103Y98_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y98_SLICE_X103Y98_A5 = CLBLM_L_X72Y98_SLICE_X108Y98_BQ;
  assign CLBLM_L_X68Y98_SLICE_X103Y98_A6 = 1'b1;
  assign CLBLM_L_X78Y130_SLICE_X120Y130_C1 = CLBLM_L_X78Y130_SLICE_X120Y130_BQ;
  assign CLBLM_L_X78Y130_SLICE_X120Y130_C2 = CLBLL_R_X77Y131_SLICE_X119Y131_AQ;
  assign CLBLM_L_X68Y98_SLICE_X103Y98_B1 = CLBLM_R_X67Y98_SLICE_X101Y98_AO5;
  assign CLBLM_L_X68Y98_SLICE_X103Y98_B2 = CLBLM_L_X68Y98_SLICE_X103Y98_BQ;
  assign CLBLM_L_X68Y98_SLICE_X103Y98_B3 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X68Y98_SLICE_X103Y98_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y98_SLICE_X103Y98_B5 = CLBLM_L_X68Y98_SLICE_X102Y98_AQ;
  assign CLBLM_L_X68Y98_SLICE_X103Y98_B6 = CLBLM_R_X67Y98_SLICE_X101Y98_BO5;
  assign CLBLM_L_X78Y130_SLICE_X120Y130_C3 = CLBLL_R_X77Y130_SLICE_X118Y130_BQ;
  assign CLBLM_L_X78Y130_SLICE_X120Y130_C4 = CLBLL_R_X77Y130_SLICE_X118Y130_AQ;
  assign CLBLM_L_X68Y98_SLICE_X103Y98_C1 = CLBLM_R_X67Y98_SLICE_X100Y98_CO6;
  assign CLBLM_L_X68Y98_SLICE_X103Y98_C2 = CLBLM_L_X68Y98_SLICE_X103Y98_CQ;
  assign CLBLM_L_X68Y98_SLICE_X103Y98_C3 = CLBLM_L_X68Y98_SLICE_X103Y98_BQ;
  assign CLBLM_L_X68Y98_SLICE_X103Y98_C4 = CLBLM_R_X67Y98_SLICE_X101Y98_BO5;
  assign CLBLM_L_X68Y98_SLICE_X103Y98_C5 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X68Y98_SLICE_X103Y98_C6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X78Y130_SLICE_X120Y130_C5 = CLBLL_R_X77Y130_SLICE_X119Y130_AO5;
  assign CLBLM_L_X78Y130_SLICE_X120Y130_C6 = CLBLL_R_X77Y130_SLICE_X119Y130_AO6;
  assign CLBLM_L_X68Y98_SLICE_X103Y98_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X68Y98_SLICE_X103Y98_D1 = CLBLM_L_X68Y98_SLICE_X102Y98_AQ;
  assign CLBLM_L_X68Y98_SLICE_X103Y98_D2 = CLBLM_L_X68Y99_SLICE_X103Y99_C5Q;
  assign CLBLM_L_X68Y98_SLICE_X103Y98_D3 = CLBLM_L_X68Y99_SLICE_X103Y99_CQ;
  assign CLBLM_L_X68Y98_SLICE_X103Y98_D4 = CLBLM_L_X68Y98_SLICE_X103Y98_BQ;
  assign CLBLM_L_X68Y98_SLICE_X103Y98_D5 = CLBLM_L_X68Y99_SLICE_X102Y99_AQ;
  assign CLBLM_L_X68Y98_SLICE_X103Y98_D6 = CLBLM_L_X68Y97_SLICE_X103Y97_AQ;
  assign CLBLL_R_X75Y103_SLICE_X114Y103_A1 = CLBLM_L_X72Y104_SLICE_X109Y104_B5Q;
  assign CLBLL_R_X75Y103_SLICE_X114Y103_A2 = CLBLM_L_X74Y104_SLICE_X112Y104_BQ;
  assign CLBLL_R_X75Y103_SLICE_X114Y103_A3 = CLBLL_R_X79Y104_SLICE_X122Y104_A5Q;
  assign CLBLL_R_X75Y103_SLICE_X114Y103_A4 = CLBLM_L_X72Y104_SLICE_X109Y104_BQ;
  assign CLBLL_R_X75Y103_SLICE_X114Y103_A5 = CLBLL_R_X75Y103_SLICE_X115Y103_AQ;
  assign CLBLL_R_X75Y103_SLICE_X114Y103_A6 = CLBLL_R_X73Y104_SLICE_X110Y104_A5Q;
  assign CLBLM_L_X68Y98_SLICE_X102Y98_A1 = CLBLM_R_X67Y98_SLICE_X100Y98_A5Q;
  assign CLBLM_L_X68Y98_SLICE_X102Y98_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y98_SLICE_X102Y98_A3 = CLBLM_L_X68Y98_SLICE_X102Y98_AQ;
  assign CLBLL_R_X75Y103_SLICE_X114Y103_B1 = CLBLM_L_X72Y104_SLICE_X109Y104_B5Q;
  assign CLBLL_R_X75Y103_SLICE_X114Y103_B2 = 1'b1;
  assign CLBLL_R_X75Y103_SLICE_X114Y103_B3 = CLBLL_R_X73Y103_SLICE_X111Y103_A5Q;
  assign CLBLL_R_X75Y103_SLICE_X114Y103_B4 = CLBLM_L_X72Y104_SLICE_X109Y104_BQ;
  assign CLBLL_R_X75Y103_SLICE_X114Y103_B5 = CLBLL_R_X75Y103_SLICE_X114Y103_AO6;
  assign CLBLL_R_X75Y103_SLICE_X114Y103_B6 = CLBLM_L_X74Y104_SLICE_X112Y104_CQ;
  assign CLBLM_L_X68Y98_SLICE_X102Y98_A4 = CLBLM_L_X68Y101_SLICE_X102Y101_BQ;
  assign CLBLM_L_X68Y98_SLICE_X102Y98_A5 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X68Y98_SLICE_X102Y98_A6 = CLBLM_R_X67Y98_SLICE_X101Y98_AO6;
  assign CLBLL_R_X75Y103_SLICE_X114Y103_C1 = 1'b1;
  assign CLBLL_R_X75Y103_SLICE_X114Y103_C2 = 1'b1;
  assign CLBLL_R_X75Y103_SLICE_X114Y103_C3 = 1'b1;
  assign CLBLL_R_X75Y103_SLICE_X114Y103_C4 = 1'b1;
  assign CLBLL_R_X75Y103_SLICE_X114Y103_C5 = 1'b1;
  assign CLBLL_R_X75Y103_SLICE_X114Y103_C6 = 1'b1;
  assign CLBLM_L_X68Y98_SLICE_X102Y98_B2 = CLBLM_L_X68Y98_SLICE_X102Y98_BQ;
  assign CLBLM_L_X68Y98_SLICE_X102Y98_B3 = CLBLM_L_X68Y99_SLICE_X103Y99_AQ;
  assign CLBLM_L_X68Y98_SLICE_X102Y98_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y98_SLICE_X102Y98_B5 = CLBLM_R_X67Y98_SLICE_X101Y98_BO6;
  assign CLBLM_L_X68Y98_SLICE_X102Y98_B6 = CLBLM_R_X67Y98_SLICE_X101Y98_AO6;
  assign CLBLM_L_X68Y98_SLICE_X102Y98_C1 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X68Y98_SLICE_X102Y98_C2 = CLBLM_L_X68Y98_SLICE_X102Y98_CQ;
  assign CLBLL_R_X75Y103_SLICE_X114Y103_D1 = 1'b1;
  assign CLBLL_R_X75Y103_SLICE_X114Y103_D2 = 1'b1;
  assign CLBLL_R_X75Y103_SLICE_X114Y103_D3 = 1'b1;
  assign CLBLL_R_X75Y103_SLICE_X114Y103_D4 = 1'b1;
  assign CLBLL_R_X75Y103_SLICE_X114Y103_D5 = 1'b1;
  assign CLBLL_R_X75Y103_SLICE_X114Y103_D6 = 1'b1;
  assign CLBLM_L_X68Y98_SLICE_X102Y98_C5 = CLBLM_R_X67Y98_SLICE_X101Y98_AO5;
  assign CLBLM_L_X68Y98_SLICE_X102Y98_D1 = CLBLM_R_X67Y97_SLICE_X100Y97_AQ;
  assign CLBLM_L_X68Y98_SLICE_X102Y98_D2 = CLBLM_R_X67Y98_SLICE_X101Y98_CO5;
  assign CLBLM_L_X68Y98_SLICE_X102Y98_D3 = CLBLM_L_X68Y98_SLICE_X102Y98_DQ;
  assign CLBLM_L_X68Y98_SLICE_X102Y98_D4 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X68Y98_SLICE_X102Y98_D5 = CLBLM_R_X67Y98_SLICE_X100Y98_CO5;
  assign CLBLM_L_X68Y98_SLICE_X102Y98_D6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X78Y130_SLICE_X120Y130_D2 = CLBLL_R_X77Y130_SLICE_X118Y130_BQ;
  assign CLBLM_L_X78Y130_SLICE_X120Y130_D3 = CLBLL_R_X77Y131_SLICE_X119Y131_AQ;
  assign CLBLM_L_X68Y98_SLICE_X102Y98_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X78Y130_SLICE_X120Y130_D4 = CLBLM_L_X78Y131_SLICE_X120Y131_AQ;
  assign CLBLM_L_X78Y130_SLICE_X120Y130_D5 = CLBLL_R_X77Y130_SLICE_X118Y130_AQ;
  assign CLBLM_L_X78Y130_SLICE_X120Y130_D6 = CLBLL_R_X77Y130_SLICE_X119Y130_AO6;
  assign CLBLL_R_X75Y103_SLICE_X115Y103_A1 = CLBLL_R_X75Y103_SLICE_X115Y103_AQ;
  assign CLBLL_R_X75Y103_SLICE_X115Y103_A2 = CLBLM_L_X62Y95_SLICE_X92Y95_AQ;
  assign CLBLL_R_X75Y103_SLICE_X115Y103_A3 = CLBLL_R_X73Y103_SLICE_X111Y103_A5Q;
  assign CLBLL_R_X75Y103_SLICE_X115Y103_A4 = CLBLL_R_X75Y103_SLICE_X115Y103_BO6;
  assign CLBLL_R_X75Y103_SLICE_X115Y103_A5 = CLBLM_L_X60Y101_SLICE_X90Y101_AQ;
  assign CLBLL_R_X75Y103_SLICE_X115Y103_A6 = CLBLL_R_X79Y104_SLICE_X122Y104_A5Q;
  assign CLBLL_R_X75Y103_SLICE_X115Y103_B1 = CLBLL_R_X75Y103_SLICE_X115Y103_AQ;
  assign CLBLL_R_X75Y103_SLICE_X115Y103_B2 = CLBLL_R_X79Y104_SLICE_X122Y104_A5Q;
  assign CLBLL_R_X75Y103_SLICE_X115Y103_B3 = CLBLL_R_X73Y103_SLICE_X111Y103_A5Q;
  assign CLBLL_R_X75Y103_SLICE_X115Y103_B4 = CLBLL_R_X73Y103_SLICE_X110Y103_A5Q;
  assign CLBLL_R_X75Y103_SLICE_X115Y103_B5 = CLBLM_L_X60Y101_SLICE_X90Y101_AQ;
  assign CLBLL_R_X75Y103_SLICE_X115Y103_B6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign RIOB33_X105Y121_IOB_X1Y122_O = CLBLM_R_X63Y98_SLICE_X94Y98_AQ;
  assign RIOB33_X105Y121_IOB_X1Y121_O = CLBLM_L_X70Y100_SLICE_X104Y100_A5Q;
  assign CLBLL_R_X75Y103_SLICE_X115Y103_C1 = 1'b1;
  assign CLBLL_R_X75Y103_SLICE_X115Y103_C2 = 1'b1;
  assign CLBLL_R_X75Y103_SLICE_X115Y103_C3 = 1'b1;
  assign CLBLL_R_X75Y103_SLICE_X115Y103_C4 = 1'b1;
  assign CLBLL_R_X75Y103_SLICE_X115Y103_C5 = 1'b1;
  assign CLBLL_R_X75Y103_SLICE_X115Y103_C6 = 1'b1;
  assign CLBLL_R_X75Y103_SLICE_X115Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X72Y109_SLICE_X109Y109_D1 = CLBLM_L_X72Y116_SLICE_X108Y116_AQ;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_D1 = CLBLL_R_X71Y119_SLICE_X106Y119_AQ;
  assign CLBLL_R_X75Y103_SLICE_X115Y103_D1 = 1'b1;
  assign CLBLL_R_X75Y103_SLICE_X115Y103_D2 = 1'b1;
  assign CLBLL_R_X75Y103_SLICE_X115Y103_D3 = 1'b1;
  assign CLBLL_R_X75Y103_SLICE_X115Y103_D4 = 1'b1;
  assign CLBLL_R_X75Y103_SLICE_X115Y103_D5 = 1'b1;
  assign CLBLL_R_X75Y103_SLICE_X115Y103_D6 = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_T1 = 1'b1;
  assign CLBLL_R_X75Y103_SLICE_X115Y103_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_D1 = CLBLM_R_X67Y116_SLICE_X100Y116_AQ;
  assign CLBLM_L_X72Y109_SLICE_X109Y109_D2 = CLBLM_L_X72Y109_SLICE_X109Y109_CQ;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_T1 = 1'b1;
  assign RIOI3_X105Y79_OLOGIC_X1Y80_D1 = 1'b0;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_A1 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_A2 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_A3 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_A4 = CLBLL_R_X73Y125_SLICE_X111Y125_A5Q;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_A5 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_A6 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_B1 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_B2 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_B3 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_B4 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_B5 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_B6 = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_D1 = CLBLL_L_X2Y131_SLICE_X0Y131_AO6;
  assign RIOI3_X105Y79_OLOGIC_X1Y80_T1 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_C1 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_C2 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_C3 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_C4 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_C5 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_C6 = 1'b1;
  assign RIOI3_X105Y79_OLOGIC_X1Y79_D1 = CLBLL_R_X83Y94_SLICE_X130Y94_A5Q;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1 = CLBLM_L_X76Y129_SLICE_X116Y129_CQ;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_D1 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_D2 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_D3 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_D4 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_D5 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_D6 = 1'b1;
  assign RIOI3_X105Y79_OLOGIC_X1Y79_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1 = 1'b0;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_A1 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_A2 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_A3 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_A4 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_A5 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_A6 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_B1 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_B2 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_B3 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_B4 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_B5 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_B6 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_C1 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_C2 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_C3 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_C4 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_C5 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_C6 = 1'b1;
  assign CLBLM_L_X72Y111_SLICE_X109Y111_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_D1 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_D2 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_D3 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_D4 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_D5 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_D6 = 1'b1;
  assign CLBLM_L_X72Y111_SLICE_X109Y111_A2 = CLBLM_L_X70Y111_SLICE_X104Y111_BQ;
  assign CLBLM_L_X72Y111_SLICE_X109Y111_A3 = CLBLM_L_X72Y111_SLICE_X109Y111_AQ;
  assign CLBLM_L_X72Y111_SLICE_X109Y111_A4 = CLBLM_L_X72Y111_SLICE_X109Y111_CQ;
  assign CLBLM_L_X72Y111_SLICE_X109Y111_A5 = CLBLM_L_X72Y111_SLICE_X109Y111_A5Q;
  assign CLBLM_L_X72Y111_SLICE_X109Y111_A6 = 1'b1;
  assign CLBLM_L_X72Y111_SLICE_X109Y111_B1 = 1'b1;
  assign CLBLM_L_X72Y111_SLICE_X109Y111_B2 = 1'b1;
  assign CLBLM_L_X72Y111_SLICE_X109Y111_B3 = 1'b1;
  assign CLBLM_L_X72Y111_SLICE_X109Y111_B4 = 1'b1;
  assign CLBLM_L_X72Y111_SLICE_X109Y111_B5 = 1'b1;
  assign CLBLM_L_X72Y111_SLICE_X109Y111_B6 = 1'b1;
  assign CLBLM_L_X72Y111_SLICE_X109Y111_BX = CLBLM_L_X72Y113_SLICE_X108Y113_BQ;
  assign CLBLM_L_X72Y111_SLICE_X109Y111_C1 = 1'b1;
  assign CLBLM_L_X72Y111_SLICE_X109Y111_C2 = 1'b1;
  assign CLBLM_L_X68Y99_SLICE_X103Y99_A1 = CLBLM_R_X67Y98_SLICE_X100Y98_B5Q;
  assign CLBLM_L_X68Y99_SLICE_X103Y99_A2 = CLBLM_L_X68Y99_SLICE_X103Y99_BQ;
  assign CLBLM_L_X68Y99_SLICE_X103Y99_A3 = CLBLM_L_X68Y99_SLICE_X103Y99_AQ;
  assign CLBLM_L_X68Y99_SLICE_X103Y99_A4 = CLBLM_R_X67Y98_SLICE_X101Y98_BO5;
  assign CLBLM_L_X68Y99_SLICE_X103Y99_A5 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X68Y99_SLICE_X103Y99_A6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y111_SLICE_X109Y111_C3 = 1'b1;
  assign CLBLM_L_X72Y111_SLICE_X109Y111_C4 = 1'b1;
  assign CLBLM_L_X72Y111_SLICE_X109Y111_C5 = 1'b1;
  assign CLBLM_L_X68Y99_SLICE_X103Y99_B1 = CLBLM_L_X68Y98_SLICE_X103Y98_CQ;
  assign CLBLM_L_X68Y99_SLICE_X103Y99_B2 = CLBLM_L_X68Y99_SLICE_X103Y99_BQ;
  assign CLBLM_L_X68Y99_SLICE_X103Y99_B3 = CLBLM_R_X67Y98_SLICE_X100Y98_CO5;
  assign CLBLM_L_X68Y99_SLICE_X103Y99_B4 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X68Y99_SLICE_X103Y99_B5 = CLBLM_R_X67Y98_SLICE_X101Y98_BO5;
  assign CLBLM_L_X68Y99_SLICE_X103Y99_B6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y111_SLICE_X109Y111_CX = CLBLM_L_X72Y111_SLICE_X108Y111_AO5;
  assign CLBLM_L_X72Y111_SLICE_X109Y111_D1 = 1'b1;
  assign CLBLM_L_X72Y111_SLICE_X109Y111_D2 = 1'b1;
  assign CLBLM_L_X68Y99_SLICE_X103Y99_C1 = CLBLM_L_X68Y99_SLICE_X103Y99_C5Q;
  assign CLBLM_L_X68Y99_SLICE_X103Y99_C2 = CLBLM_L_X68Y99_SLICE_X103Y99_CQ;
  assign CLBLM_L_X68Y99_SLICE_X103Y99_C3 = CLBLM_L_X70Y106_SLICE_X104Y106_CO6;
  assign CLBLM_L_X68Y99_SLICE_X103Y99_C4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y99_SLICE_X103Y99_C5 = CLBLM_L_X68Y99_SLICE_X103Y99_D5Q;
  assign CLBLM_L_X68Y99_SLICE_X103Y99_C6 = 1'b1;
  assign CLBLM_L_X72Y111_SLICE_X108Y111_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y111_SLICE_X108Y111_A2 = CLBLM_L_X72Y111_SLICE_X109Y111_CQ;
  assign CLBLM_L_X68Y99_SLICE_X103Y99_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X72Y111_SLICE_X108Y111_A3 = CLBLM_L_X72Y111_SLICE_X108Y111_DQ;
  assign CLBLM_L_X72Y111_SLICE_X108Y111_A4 = CLBLM_L_X70Y111_SLICE_X104Y111_BQ;
  assign CLBLM_L_X72Y111_SLICE_X108Y111_A5 = CLBLM_L_X72Y111_SLICE_X109Y111_AQ;
  assign CLBLM_L_X72Y111_SLICE_X108Y111_A6 = 1'b1;
  assign CLBLM_L_X68Y99_SLICE_X103Y99_D1 = CLBLM_L_X68Y98_SLICE_X103Y98_A5Q;
  assign CLBLM_L_X68Y99_SLICE_X103Y99_D2 = CLBLM_L_X68Y96_SLICE_X103Y96_BO6;
  assign CLBLM_L_X68Y99_SLICE_X103Y99_D3 = CLBLM_L_X68Y99_SLICE_X103Y99_DQ;
  assign CLBLM_L_X68Y99_SLICE_X103Y99_D4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y99_SLICE_X103Y99_D5 = CLBLM_L_X68Y99_SLICE_X103Y99_D5Q;
  assign CLBLM_L_X68Y99_SLICE_X103Y99_D6 = 1'b1;
  assign CLBLM_L_X72Y111_SLICE_X108Y111_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y99_SLICE_X103Y99_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y111_SLICE_X108Y111_B2 = CLBLM_L_X72Y111_SLICE_X108Y111_BQ;
  assign CLBLM_L_X72Y111_SLICE_X108Y111_B3 = CLBLM_L_X72Y109_SLICE_X108Y109_AO6;
  assign CLBLM_L_X72Y111_SLICE_X108Y111_B4 = 1'b1;
  assign CLBLM_L_X68Y99_SLICE_X102Y99_A1 = CLBLM_L_X70Y106_SLICE_X104Y106_CO6;
  assign CLBLM_L_X68Y99_SLICE_X102Y99_A2 = CLBLM_L_X68Y98_SLICE_X103Y98_A5Q;
  assign CLBLM_L_X68Y99_SLICE_X102Y99_A3 = CLBLM_L_X68Y99_SLICE_X103Y99_C5Q;
  assign CLBLM_L_X68Y99_SLICE_X102Y99_A4 = CLBLM_L_X60Y94_SLICE_X90Y94_CQ;
  assign CLBLM_L_X68Y99_SLICE_X102Y99_A5 = CLBLM_L_X68Y99_SLICE_X103Y99_CQ;
  assign CLBLM_L_X68Y99_SLICE_X102Y99_A6 = 1'b1;
  assign CLBLM_L_X72Y111_SLICE_X108Y111_C1 = CLBLM_L_X72Y109_SLICE_X108Y109_AO6;
  assign CLBLM_L_X72Y111_SLICE_X108Y111_C2 = CLBLM_L_X78Y123_SLICE_X121Y123_A5Q;
  assign CLBLM_L_X72Y109_SLICE_X109Y109_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X68Y99_SLICE_X102Y99_AX = CLBLM_L_X60Y94_SLICE_X90Y94_CQ;
  assign CLBLM_L_X72Y111_SLICE_X108Y111_C4 = CLBLM_L_X70Y112_SLICE_X104Y112_CQ;
  assign CLBLM_L_X68Y99_SLICE_X102Y99_B1 = CLBLM_L_X68Y95_SLICE_X102Y95_AQ;
  assign CLBLM_L_X68Y99_SLICE_X102Y99_B2 = CLBLM_L_X68Y98_SLICE_X103Y98_A5Q;
  assign CLBLM_L_X68Y99_SLICE_X102Y99_B3 = CLBLM_L_X68Y99_SLICE_X103Y99_C5Q;
  assign CLBLM_L_X68Y99_SLICE_X102Y99_B4 = CLBLM_L_X68Y98_SLICE_X102Y98_BQ;
  assign CLBLM_L_X68Y99_SLICE_X102Y99_B5 = CLBLM_L_X68Y99_SLICE_X103Y99_CQ;
  assign CLBLM_L_X68Y99_SLICE_X102Y99_B6 = 1'b1;
  assign CLBLM_L_X72Y111_SLICE_X108Y111_D1 = CLBLM_L_X72Y111_SLICE_X109Y111_AQ;
  assign CLBLM_L_X72Y111_SLICE_X108Y111_D2 = CLBLM_L_X72Y111_SLICE_X109Y111_A5Q;
  assign CLBLM_L_X72Y111_SLICE_X108Y111_D3 = CLBLM_L_X72Y111_SLICE_X108Y111_DQ;
  assign CLBLM_L_X68Y99_SLICE_X102Y99_C1 = CLBLM_L_X68Y99_SLICE_X102Y99_AO6;
  assign CLBLM_L_X68Y99_SLICE_X102Y99_C2 = CLBLM_L_X68Y99_SLICE_X103Y99_AQ;
  assign CLBLM_L_X68Y99_SLICE_X102Y99_C3 = CLBLM_L_X68Y97_SLICE_X102Y97_AQ;
  assign CLBLM_L_X68Y99_SLICE_X102Y99_C4 = CLBLM_L_X68Y98_SLICE_X103Y98_A5Q;
  assign CLBLM_L_X68Y99_SLICE_X102Y99_C5 = CLBLM_L_X68Y99_SLICE_X102Y99_BO5;
  assign CLBLM_L_X68Y99_SLICE_X102Y99_C6 = CLBLM_L_X68Y99_SLICE_X102Y99_DO6;
  assign CLBLM_L_X72Y111_SLICE_X108Y111_D6 = CLBLM_L_X70Y111_SLICE_X104Y111_BQ;
  assign CLBLM_L_X72Y111_SLICE_X108Y111_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X68Y99_SLICE_X102Y99_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X68Y99_SLICE_X102Y99_D1 = CLBLM_L_X68Y98_SLICE_X103Y98_A5Q;
  assign CLBLM_L_X68Y99_SLICE_X102Y99_D2 = CLBLM_L_X68Y101_SLICE_X102Y101_CQ;
  assign CLBLM_L_X68Y99_SLICE_X102Y99_D3 = CLBLM_L_X68Y99_SLICE_X103Y99_C5Q;
  assign CLBLM_L_X68Y99_SLICE_X102Y99_D4 = CLBLM_L_X68Y99_SLICE_X103Y99_CQ;
  assign CLBLM_L_X68Y99_SLICE_X102Y99_D5 = 1'b1;
  assign CLBLM_L_X68Y99_SLICE_X102Y99_D6 = CLBLM_L_X60Y94_SLICE_X90Y94_CQ;
  assign CLBLM_L_X68Y99_SLICE_X102Y99_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign RIOB33_X105Y123_IOB_X1Y124_O = CLBLM_L_X68Y99_SLICE_X102Y99_AQ;
  assign RIOB33_X105Y123_IOB_X1Y123_O = CLBLM_R_X63Y101_SLICE_X94Y101_AQ;
  assign CLBLM_L_X68Y100_SLICE_X103Y100_A1 = CLBLM_L_X68Y105_SLICE_X103Y105_BQ;
  assign CLBLM_L_X68Y100_SLICE_X103Y100_A2 = CLBLM_L_X70Y106_SLICE_X104Y106_CO6;
  assign CLBLM_L_X68Y100_SLICE_X103Y100_A3 = CLBLM_L_X68Y99_SLICE_X103Y99_D5Q;
  assign CLBLM_L_X68Y100_SLICE_X103Y100_A4 = CLBLM_L_X68Y99_SLICE_X103Y99_C5Q;
  assign CLBLM_L_X68Y100_SLICE_X103Y100_A5 = CLBLM_L_X68Y99_SLICE_X103Y99_DQ;
  assign CLBLM_L_X68Y100_SLICE_X103Y100_A6 = CLBLM_L_X68Y99_SLICE_X103Y99_CQ;
  assign CLBLM_L_X68Y100_SLICE_X103Y100_B1 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X103Y100_B2 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X103Y100_B3 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X103Y100_B4 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X103Y100_B5 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X103Y100_B6 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X103Y100_C1 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X103Y100_C2 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X103Y100_C3 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X103Y100_C4 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X103Y100_C5 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X103Y100_C6 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X103Y100_D1 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X103Y100_D2 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X103Y100_D3 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X103Y100_D4 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X103Y100_D5 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X103Y100_D6 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X102Y100_A1 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X102Y100_A2 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X102Y100_A3 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X102Y100_A4 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X102Y100_A5 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X102Y100_A6 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X102Y100_B1 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X102Y100_B2 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X102Y100_B3 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X102Y100_B4 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X102Y100_B5 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X102Y100_B6 = 1'b1;
  assign RIOB33_X105Y125_IOB_X1Y126_O = CLBLM_L_X76Y127_SLICE_X116Y127_AQ;
  assign CLBLM_L_X62Y90_SLICE_X93Y90_D1 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X102Y100_C1 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X102Y100_C2 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X102Y100_C3 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X102Y100_C4 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X102Y100_C5 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X102Y100_C6 = 1'b1;
  assign RIOB33_X105Y125_IOB_X1Y125_O = CLBLM_L_X74Y129_SLICE_X112Y129_BQ;
  assign CLBLM_L_X68Y100_SLICE_X102Y100_D1 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X102Y100_D2 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X102Y100_D3 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X102Y100_D4 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X102Y100_D5 = 1'b1;
  assign CLBLM_L_X68Y100_SLICE_X102Y100_D6 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X93Y90_D5 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_D3 = CLBLM_L_X72Y131_SLICE_X109Y131_DQ;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_D5 = CLBLM_L_X72Y131_SLICE_X108Y131_A5Q;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_D6 = CLBLM_L_X72Y133_SLICE_X109Y133_DO6;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_A2 = CLBLM_L_X72Y133_SLICE_X109Y133_DO6;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_A3 = CLBLM_L_X72Y131_SLICE_X108Y131_AQ;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_A4 = CLBLM_L_X72Y130_SLICE_X108Y130_AQ;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_A5 = CLBLM_L_X72Y131_SLICE_X108Y131_A5Q;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_A6 = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_D1 = CLBLL_R_X71Y124_SLICE_X106Y124_AQ;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_B1 = CLBLM_L_X72Y134_SLICE_X109Y134_AO5;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_T1 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_B2 = CLBLM_L_X72Y130_SLICE_X108Y130_AQ;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_B3 = CLBLM_L_X72Y131_SLICE_X109Y131_AO6;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_D1 = CLBLM_L_X70Y110_SLICE_X104Y110_CQ;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_B4 = CLBLM_L_X72Y131_SLICE_X109Y131_BQ;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_T1 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X109Y113_A1 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X109Y113_A2 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X109Y113_A3 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X109Y113_A4 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X109Y113_A5 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X109Y113_A6 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_B6 = CLBLM_L_X72Y131_SLICE_X108Y131_BQ;
  assign CLBLM_L_X76Y134_SLICE_X116Y134_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y113_SLICE_X109Y113_B1 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X109Y113_B2 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X109Y113_B3 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X109Y113_B4 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X109Y113_B5 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X109Y113_B6 = 1'b1;
  assign RIOI3_X105Y83_OLOGIC_X1Y84_D1 = CLBLM_L_X72Y118_SLICE_X108Y118_D5Q;
  assign CLBLM_L_X72Y113_SLICE_X109Y113_C1 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X109Y113_C2 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X109Y113_C3 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X109Y113_C4 = 1'b1;
  assign CLBLM_L_X68Y101_SLICE_X103Y101_A1 = 1'b1;
  assign CLBLM_L_X68Y101_SLICE_X103Y101_A2 = 1'b1;
  assign CLBLM_L_X68Y101_SLICE_X103Y101_A3 = 1'b1;
  assign CLBLM_L_X68Y101_SLICE_X103Y101_A4 = 1'b1;
  assign CLBLM_L_X68Y101_SLICE_X103Y101_A5 = 1'b1;
  assign CLBLM_L_X68Y101_SLICE_X103Y101_A6 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X109Y113_C5 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X109Y113_C6 = 1'b1;
  assign CLBLM_L_X68Y101_SLICE_X103Y101_B1 = 1'b1;
  assign CLBLM_L_X68Y101_SLICE_X103Y101_B2 = 1'b1;
  assign CLBLM_L_X68Y101_SLICE_X103Y101_B3 = 1'b1;
  assign CLBLM_L_X68Y101_SLICE_X103Y101_B4 = 1'b1;
  assign CLBLM_L_X68Y101_SLICE_X103Y101_B5 = 1'b1;
  assign CLBLM_L_X68Y101_SLICE_X103Y101_B6 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X92Y90_D2 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X109Y113_D1 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X109Y113_D2 = 1'b1;
  assign CLBLM_L_X68Y101_SLICE_X103Y101_C1 = 1'b1;
  assign CLBLM_L_X68Y101_SLICE_X103Y101_C2 = 1'b1;
  assign CLBLM_L_X68Y101_SLICE_X103Y101_C3 = 1'b1;
  assign CLBLM_L_X68Y101_SLICE_X103Y101_C4 = 1'b1;
  assign CLBLM_L_X68Y101_SLICE_X103Y101_C5 = 1'b1;
  assign CLBLM_L_X68Y101_SLICE_X103Y101_C6 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X108Y113_A1 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X108Y113_A2 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X108Y113_A3 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X108Y113_A4 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X108Y113_A5 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X108Y113_A6 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_C5 = CLBLM_L_X72Y131_SLICE_X108Y131_DO6;
  assign CLBLM_L_X72Y113_SLICE_X108Y113_AX = CLBLM_L_X70Y108_SLICE_X105Y108_AO5;
  assign CLBLM_L_X68Y101_SLICE_X103Y101_D1 = 1'b1;
  assign CLBLM_L_X68Y101_SLICE_X103Y101_D2 = 1'b1;
  assign CLBLM_L_X68Y101_SLICE_X103Y101_D3 = 1'b1;
  assign CLBLM_L_X68Y101_SLICE_X103Y101_D4 = 1'b1;
  assign CLBLM_L_X68Y101_SLICE_X103Y101_D5 = 1'b1;
  assign CLBLM_L_X68Y101_SLICE_X103Y101_D6 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X108Y113_B1 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X108Y113_B2 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X108Y113_B3 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X108Y113_B4 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X108Y113_B5 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X108Y113_B6 = 1'b1;
  assign CLBLM_L_X68Y101_SLICE_X102Y101_A1 = 1'b1;
  assign CLBLM_L_X68Y101_SLICE_X102Y101_A2 = CLBLM_L_X68Y105_SLICE_X102Y105_AQ;
  assign CLBLM_L_X68Y101_SLICE_X102Y101_A3 = CLBLM_L_X68Y101_SLICE_X102Y101_AQ;
  assign CLBLM_L_X68Y101_SLICE_X102Y101_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y101_SLICE_X102Y101_A5 = CLBLM_L_X64Y101_SLICE_X96Y101_AQ;
  assign CLBLM_L_X68Y101_SLICE_X102Y101_A6 = CLBLM_L_X68Y101_SLICE_X102Y101_A5Q;
  assign CLBLM_L_X72Y113_SLICE_X108Y113_C1 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X108Y113_C2 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X108Y113_C3 = 1'b1;
  assign CLBLM_L_X68Y101_SLICE_X102Y101_AX = CLBLM_L_X68Y105_SLICE_X102Y105_AQ;
  assign CLBLM_L_X72Y113_SLICE_X108Y113_C4 = 1'b1;
  assign CLBLM_L_X68Y101_SLICE_X102Y101_B1 = CLBLM_R_X67Y98_SLICE_X100Y98_B5Q;
  assign CLBLM_L_X68Y101_SLICE_X102Y101_B2 = CLBLM_L_X68Y101_SLICE_X102Y101_BQ;
  assign CLBLM_L_X68Y101_SLICE_X102Y101_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y101_SLICE_X102Y101_B4 = CLBLM_R_X67Y98_SLICE_X100Y98_A5Q;
  assign CLBLM_L_X68Y101_SLICE_X102Y101_B5 = 1'b1;
  assign CLBLM_L_X68Y101_SLICE_X102Y101_B6 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X108Y113_D1 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X108Y113_D2 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X108Y113_D3 = 1'b1;
  assign CLBLM_L_X68Y101_SLICE_X102Y101_C1 = 1'b1;
  assign CLBLM_L_X68Y101_SLICE_X102Y101_C2 = CLBLM_L_X68Y101_SLICE_X102Y101_CQ;
  assign CLBLM_L_X68Y101_SLICE_X102Y101_C3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y101_SLICE_X102Y101_C4 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X68Y101_SLICE_X102Y101_C5 = CLBLM_L_X68Y101_SLICE_X102Y101_BO5;
  assign CLBLM_L_X68Y101_SLICE_X102Y101_C6 = CLBLM_L_X68Y98_SLICE_X102Y98_DQ;
  assign CLBLM_L_X72Y113_SLICE_X108Y113_D6 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X108Y113_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X68Y101_SLICE_X102Y101_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X68Y101_SLICE_X102Y101_D1 = 1'b1;
  assign CLBLM_L_X68Y101_SLICE_X102Y101_D2 = 1'b1;
  assign CLBLM_L_X68Y101_SLICE_X102Y101_D3 = 1'b1;
  assign CLBLM_L_X68Y101_SLICE_X102Y101_D4 = 1'b1;
  assign CLBLM_L_X68Y101_SLICE_X102Y101_D5 = 1'b1;
  assign CLBLM_L_X68Y101_SLICE_X102Y101_D6 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_D1 = CLBLM_L_X72Y130_SLICE_X108Y130_AQ;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_D2 = 1'b1;
  assign CLBLM_L_X68Y101_SLICE_X102Y101_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_D3 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_D4 = CLBLM_L_X72Y131_SLICE_X108Y131_A5Q;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_D5 = CLBLM_L_X72Y133_SLICE_X109Y133_DO6;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_D6 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X79Y135_SLICE_X122Y135_A1 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X122Y135_A2 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X122Y135_A3 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X122Y135_A4 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X122Y135_A5 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X122Y135_A6 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_C1 = CLBLM_L_X74Y126_SLICE_X113Y126_BQ;
  assign CLBLL_R_X79Y135_SLICE_X122Y135_AX = CLBLL_R_X75Y133_SLICE_X114Y133_BQ;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_C2 = CLBLM_L_X74Y126_SLICE_X113Y126_CQ;
  assign CLBLL_R_X79Y135_SLICE_X122Y135_B1 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X122Y135_B2 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X122Y135_B3 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X122Y135_B4 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X122Y135_B5 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X122Y135_B6 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_C3 = CLBLM_L_X74Y126_SLICE_X113Y126_AQ;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_C4 = CLBLM_L_X74Y126_SLICE_X113Y126_A5Q;
  assign CLBLL_R_X79Y135_SLICE_X122Y135_C1 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X122Y135_C2 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X122Y135_C3 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X122Y135_C4 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X122Y135_C5 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X122Y135_C6 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_C5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X79Y135_SLICE_X122Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_C6 = CLBLL_R_X75Y128_SLICE_X115Y128_AO6;
  assign CLBLL_R_X79Y135_SLICE_X122Y135_D1 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X122Y135_D2 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X122Y135_D3 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X122Y135_D4 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X122Y135_D5 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X122Y135_D6 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X122Y135_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X79Y135_SLICE_X123Y135_A1 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X123Y135_A2 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X123Y135_A3 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X123Y135_A4 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X123Y135_A5 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X123Y135_A6 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_D1 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X123Y135_B1 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X123Y135_B2 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X123Y135_B3 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X123Y135_B4 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X123Y135_B5 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X123Y135_B6 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_D2 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_D3 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X123Y135_C1 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X123Y135_C2 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X123Y135_C3 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X123Y135_C4 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X123Y135_C5 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X123Y135_C6 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_D4 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_D5 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X123Y135_D1 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X123Y135_D2 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X123Y135_D3 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X123Y135_D4 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X123Y135_D5 = 1'b1;
  assign CLBLL_R_X79Y135_SLICE_X123Y135_D6 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_D6 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X78Y131_SLICE_X121Y131_A4 = 1'b1;
  assign CLBLM_L_X78Y131_SLICE_X121Y131_A5 = 1'b1;
  assign CLBLM_L_X78Y131_SLICE_X121Y131_A6 = 1'b1;
  assign CLBLM_L_X68Y102_SLICE_X103Y102_A1 = 1'b1;
  assign CLBLM_L_X68Y102_SLICE_X103Y102_A2 = 1'b1;
  assign CLBLM_L_X68Y102_SLICE_X103Y102_A3 = 1'b1;
  assign CLBLM_L_X68Y102_SLICE_X103Y102_A4 = 1'b1;
  assign CLBLM_L_X68Y102_SLICE_X103Y102_A5 = 1'b1;
  assign CLBLM_L_X68Y102_SLICE_X103Y102_A6 = 1'b1;
  assign RIOB33_X105Y129_IOB_X1Y129_O = CLBLM_L_X78Y106_SLICE_X120Y106_AQ;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_A1 = CLBLL_R_X75Y128_SLICE_X114Y128_AO6;
  assign RIOB33_X105Y129_IOB_X1Y130_O = CLBLL_R_X73Y103_SLICE_X110Y103_B5Q;
  assign CLBLM_L_X68Y102_SLICE_X103Y102_B1 = 1'b1;
  assign CLBLM_L_X68Y102_SLICE_X103Y102_B2 = 1'b1;
  assign CLBLM_L_X68Y102_SLICE_X103Y102_B3 = 1'b1;
  assign CLBLM_L_X68Y102_SLICE_X103Y102_B4 = 1'b1;
  assign CLBLM_L_X68Y102_SLICE_X103Y102_B5 = 1'b1;
  assign CLBLM_L_X68Y102_SLICE_X103Y102_B6 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_A2 = CLBLM_L_X74Y126_SLICE_X112Y126_A5Q;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_A3 = CLBLM_L_X74Y126_SLICE_X112Y126_AQ;
  assign CLBLM_L_X68Y102_SLICE_X103Y102_C1 = 1'b1;
  assign CLBLM_L_X68Y102_SLICE_X103Y102_C2 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X114Y107_A1 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X114Y107_A2 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X93Y90_A1 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X93Y90_A2 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X93Y90_A3 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X93Y90_A4 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X93Y90_A5 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X93Y90_A6 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X114Y107_A3 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X114Y107_A4 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X114Y107_A5 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X93Y90_B1 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X93Y90_B2 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X93Y90_B3 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X93Y90_B4 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X93Y90_B5 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X93Y90_B6 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X114Y107_B1 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X114Y107_B2 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X114Y107_B3 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X93Y90_C1 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X93Y90_C2 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X93Y90_C3 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X93Y90_C4 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X93Y90_C5 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X93Y90_C6 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X114Y107_C1 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X114Y107_C2 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X114Y107_C3 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X114Y107_C4 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X114Y107_C5 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X114Y107_C6 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X114Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X75Y107_SLICE_X114Y107_D1 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X114Y107_D2 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X114Y107_D3 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X114Y107_D4 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X114Y107_D5 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X93Y90_D6 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X114Y107_D6 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X114Y107_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X62Y90_SLICE_X93Y90_D2 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X93Y90_D3 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X93Y90_D4 = 1'b1;
  assign CLBLM_L_X68Y102_SLICE_X102Y102_C3 = CLBLM_L_X68Y102_SLICE_X102Y102_AQ;
  assign CLBLM_L_X68Y102_SLICE_X102Y102_C4 = CLBLM_L_X68Y99_SLICE_X102Y99_AO5;
  assign CLBLM_L_X62Y90_SLICE_X92Y90_A1 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X92Y90_A2 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X92Y90_A3 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X92Y90_A4 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X92Y90_A5 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X92Y90_A6 = 1'b1;
  assign CLBLM_L_X68Y102_SLICE_X102Y102_C6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X62Y90_SLICE_X92Y90_AX = CLBLM_L_X72Y106_SLICE_X108Y106_A5Q;
  assign CLBLM_L_X68Y102_SLICE_X102Y102_C5 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X92Y90_B1 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X92Y90_B2 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X92Y90_B3 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X92Y90_B4 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X92Y90_B5 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X92Y90_B6 = 1'b1;
  assign CLBLM_L_X68Y102_SLICE_X102Y102_D2 = CLBLM_R_X67Y98_SLICE_X100Y98_A5Q;
  assign CLBLM_L_X68Y102_SLICE_X102Y102_D3 = CLBLM_L_X68Y102_SLICE_X102Y102_DQ;
  assign CLBLM_L_X68Y102_SLICE_X102Y102_D4 = CLBLL_R_X79Y99_SLICE_X122Y99_AO6;
  assign CLBLL_R_X75Y107_SLICE_X115Y107_A1 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X115Y107_A2 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X115Y107_A3 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X115Y107_A4 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X92Y90_C3 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X92Y90_C4 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X92Y90_C5 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X92Y90_C6 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X115Y107_A5 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X115Y107_A6 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X92Y90_C1 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X92Y90_C2 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X115Y107_B1 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X115Y107_B2 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X115Y107_B3 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X115Y107_B4 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X115Y107_B5 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X115Y107_B6 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X92Y90_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X62Y90_SLICE_X92Y90_D1 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X115Y107_C1 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X115Y107_C2 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X115Y107_C3 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X115Y107_C4 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X115Y107_C5 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X115Y107_C6 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X92Y90_D3 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X92Y90_D4 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X92Y90_D5 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X92Y90_D6 = 1'b1;
  assign CLBLM_L_X62Y90_SLICE_X92Y90_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X75Y107_SLICE_X115Y107_D1 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X115Y107_D2 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X115Y107_D3 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X115Y107_D4 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X115Y107_D5 = 1'b1;
  assign CLBLL_R_X75Y107_SLICE_X115Y107_D6 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_C3 = CLBLM_L_X74Y125_SLICE_X112Y125_AQ;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_C4 = CLBLM_L_X74Y126_SLICE_X112Y126_A5Q;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_C5 = CLBLL_R_X75Y128_SLICE_X115Y128_AO6;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_C6 = 1'b1;
  assign LIOB33_X0Y59_IOB_X0Y60_O = CLBLM_L_X72Y106_SLICE_X108Y106_A5Q;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOB33_X0Y59_IOB_X0Y59_O = CLBLM_L_X60Y101_SLICE_X90Y101_AQ;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_D1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_B1 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_D2 = CLBLM_L_X74Y126_SLICE_X112Y126_AQ;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_B2 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_D3 = CLBLL_R_X75Y128_SLICE_X114Y128_AO6;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_B3 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_D4 = CLBLM_L_X74Y126_SLICE_X112Y126_DQ;
  assign CLBLM_L_X78Y131_SLICE_X120Y131_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_D5 = CLBLM_L_X74Y126_SLICE_X112Y126_BO5;
  assign CLBLM_L_X78Y131_SLICE_X120Y131_A2 = CLBLM_L_X78Y130_SLICE_X120Y130_CO6;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_D6 = CLBLL_R_X75Y128_SLICE_X115Y128_AO6;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_B6 = 1'b1;
  assign CLBLM_L_X78Y131_SLICE_X120Y131_A3 = CLBLM_L_X78Y131_SLICE_X120Y131_AQ;
  assign CLBLM_L_X78Y131_SLICE_X120Y131_A4 = CLBLL_R_X77Y130_SLICE_X119Y130_AQ;
  assign CLBLM_L_X78Y131_SLICE_X120Y131_A5 = CLBLL_R_X77Y128_SLICE_X118Y128_BQ;
  assign CLBLM_L_X78Y131_SLICE_X120Y131_A6 = CLBLL_R_X77Y128_SLICE_X118Y128_AQ;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_C1 = 1'b1;
  assign CLBLM_L_X76Y123_SLICE_X116Y123_A5 = CLBLM_L_X76Y122_SLICE_X116Y122_BQ;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_C2 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_C3 = 1'b1;
  assign CLBLM_L_X78Y131_SLICE_X120Y131_B1 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_C6 = 1'b1;
  assign CLBLM_L_X78Y131_SLICE_X120Y131_B2 = 1'b1;
  assign CLBLM_L_X76Y123_SLICE_X116Y123_A6 = CLBLL_R_X75Y123_SLICE_X115Y123_DO6;
  assign CLBLM_L_X78Y131_SLICE_X120Y131_B3 = 1'b1;
  assign CLBLM_L_X78Y131_SLICE_X120Y131_B4 = 1'b1;
  assign RIOB33_X105Y131_IOB_X1Y132_O = CLBLL_R_X79Y104_SLICE_X122Y104_A5Q;
  assign CLBLM_L_X78Y131_SLICE_X120Y131_B5 = 1'b1;
  assign RIOB33_X105Y131_IOB_X1Y131_O = CLBLM_L_X76Y111_SLICE_X116Y111_AQ;
  assign CLBLM_L_X78Y131_SLICE_X120Y131_B6 = 1'b1;
  assign CLBLM_L_X68Y103_SLICE_X103Y103_A1 = 1'b1;
  assign CLBLM_L_X68Y103_SLICE_X103Y103_A2 = 1'b1;
  assign CLBLM_L_X68Y103_SLICE_X103Y103_A3 = 1'b1;
  assign CLBLM_L_X68Y103_SLICE_X103Y103_A4 = 1'b1;
  assign CLBLM_L_X68Y103_SLICE_X103Y103_A5 = 1'b1;
  assign CLBLM_L_X68Y103_SLICE_X103Y103_A6 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_D1 = 1'b1;
  assign CLBLM_L_X68Y103_SLICE_X103Y103_B1 = 1'b1;
  assign CLBLM_L_X68Y103_SLICE_X103Y103_B2 = 1'b1;
  assign CLBLM_L_X68Y103_SLICE_X103Y103_B3 = 1'b1;
  assign CLBLM_L_X68Y103_SLICE_X103Y103_B4 = 1'b1;
  assign CLBLM_L_X68Y103_SLICE_X103Y103_B5 = 1'b1;
  assign CLBLM_L_X68Y103_SLICE_X103Y103_B6 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_D2 = 1'b1;
  assign CLBLM_L_X78Y131_SLICE_X120Y131_C1 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_D3 = 1'b1;
  assign CLBLM_L_X68Y103_SLICE_X103Y103_C1 = 1'b1;
  assign CLBLM_L_X68Y103_SLICE_X103Y103_C2 = 1'b1;
  assign CLBLM_L_X68Y103_SLICE_X103Y103_C3 = 1'b1;
  assign CLBLM_L_X68Y103_SLICE_X103Y103_C4 = 1'b1;
  assign CLBLM_L_X68Y103_SLICE_X103Y103_C5 = 1'b1;
  assign CLBLM_L_X68Y103_SLICE_X103Y103_C6 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_D4 = 1'b1;
  assign CLBLM_L_X78Y131_SLICE_X120Y131_C3 = 1'b1;
  assign CLBLM_L_X78Y131_SLICE_X120Y131_C4 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_D5 = 1'b1;
  assign CLBLM_L_X78Y131_SLICE_X120Y131_C5 = 1'b1;
  assign CLBLM_R_X67Y96_SLICE_X101Y96_A6 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_D6 = 1'b1;
  assign CLBLM_L_X68Y103_SLICE_X103Y103_D1 = 1'b1;
  assign CLBLM_L_X68Y103_SLICE_X103Y103_D2 = 1'b1;
  assign CLBLM_L_X68Y103_SLICE_X103Y103_D3 = 1'b1;
  assign CLBLM_L_X68Y103_SLICE_X103Y103_D4 = 1'b1;
  assign CLBLM_L_X68Y103_SLICE_X103Y103_D5 = 1'b1;
  assign CLBLM_L_X68Y103_SLICE_X103Y103_D6 = 1'b1;
  assign CLBLM_L_X78Y131_SLICE_X120Y131_C6 = 1'b1;
  assign CLBLM_L_X68Y103_SLICE_X102Y103_A1 = 1'b1;
  assign CLBLM_L_X68Y103_SLICE_X102Y103_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y103_SLICE_X102Y103_A3 = CLBLM_L_X68Y103_SLICE_X102Y103_AQ;
  assign CLBLM_L_X68Y103_SLICE_X102Y103_A4 = CLBLM_L_X70Y106_SLICE_X104Y106_CO6;
  assign CLBLM_L_X68Y103_SLICE_X102Y103_A5 = CLBLM_L_X68Y97_SLICE_X102Y97_CO6;
  assign CLBLM_L_X68Y103_SLICE_X102Y103_A6 = CLBLM_L_X68Y101_SLICE_X102Y101_CQ;
  assign CLBLM_L_X78Y131_SLICE_X120Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X67Y96_SLICE_X101Y96_B1 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X68Y103_SLICE_X102Y103_B1 = CLBLM_L_X68Y103_SLICE_X102Y103_B5Q;
  assign CLBLM_L_X68Y103_SLICE_X102Y103_B2 = CLBLM_L_X68Y103_SLICE_X102Y103_BQ;
  assign CLBLM_L_X68Y103_SLICE_X102Y103_B3 = CLBLM_L_X68Y99_SLICE_X102Y99_AO5;
  assign CLBLM_L_X68Y103_SLICE_X102Y103_B4 = CLBLM_R_X67Y103_SLICE_X101Y103_AQ;
  assign CLBLM_L_X68Y103_SLICE_X102Y103_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y103_SLICE_X102Y103_B6 = 1'b1;
  assign CLBLM_R_X67Y96_SLICE_X101Y96_B2 = CLBLM_R_X67Y96_SLICE_X101Y96_BQ;
  assign CLBLM_R_X67Y96_SLICE_X101Y96_B3 = CLBLM_R_X67Y96_SLICE_X101Y96_DQ;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_T1 = 1'b1;
  assign CLBLM_L_X68Y103_SLICE_X102Y103_C1 = CLBLM_L_X68Y101_SLICE_X102Y101_BQ;
  assign CLBLM_L_X68Y103_SLICE_X102Y103_C2 = CLBLM_L_X68Y103_SLICE_X102Y103_CQ;
  assign CLBLM_L_X68Y103_SLICE_X102Y103_C3 = CLBLM_R_X67Y98_SLICE_X100Y98_B5Q;
  assign CLBLM_L_X68Y103_SLICE_X102Y103_C4 = CLBLM_R_X67Y103_SLICE_X100Y103_B5Q;
  assign CLBLM_L_X68Y103_SLICE_X102Y103_C5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y103_SLICE_X102Y103_C6 = CLBLM_R_X67Y98_SLICE_X100Y98_A5Q;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_A1 = CLBLL_R_X75Y134_SLICE_X115Y134_AQ;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_D1 = CLBLL_L_X34Y123_SLICE_X50Y123_AO6;
  assign CLBLM_L_X68Y103_SLICE_X102Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_A3 = CLBLM_L_X76Y133_SLICE_X116Y133_AQ;
  assign CLBLM_L_X68Y103_SLICE_X102Y103_D1 = CLBLM_L_X68Y103_SLICE_X102Y103_DQ;
  assign CLBLM_L_X68Y103_SLICE_X102Y103_D2 = CLBLM_L_X68Y103_SLICE_X102Y103_CQ;
  assign CLBLM_L_X68Y103_SLICE_X102Y103_D3 = CLBLM_L_X68Y101_SLICE_X102Y101_BO5;
  assign CLBLM_L_X68Y103_SLICE_X102Y103_D4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y103_SLICE_X102Y103_D5 = 1'b1;
  assign CLBLM_L_X68Y103_SLICE_X102Y103_D6 = CLBLM_R_X67Y103_SLICE_X100Y103_B5Q;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_A4 = CLBLM_L_X76Y134_SLICE_X117Y134_CO6;
  assign CLBLM_L_X78Y131_SLICE_X120Y131_D1 = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_T1 = 1'b1;
  assign CLBLM_L_X68Y103_SLICE_X102Y103_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_A5 = CLBLL_R_X75Y133_SLICE_X115Y133_BQ;
  assign CLBLM_L_X78Y131_SLICE_X120Y131_D2 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_A6 = CLBLL_R_X75Y133_SLICE_X115Y133_AQ;
  assign CLBLM_L_X78Y131_SLICE_X120Y131_D3 = 1'b1;
  assign RIOI3_X105Y85_OLOGIC_X1Y86_D1 = CLBLM_L_X64Y99_SLICE_X97Y99_A5Q;
  assign CLBLL_R_X77Y121_SLICE_X119Y121_C6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X78Y131_SLICE_X120Y131_D4 = 1'b1;
  assign CLBLM_L_X78Y131_SLICE_X120Y131_D5 = 1'b1;
  assign RIOI3_X105Y85_OLOGIC_X1Y86_T1 = 1'b1;
  assign CLBLM_L_X78Y131_SLICE_X120Y131_D6 = 1'b1;
  assign CLBLM_R_X67Y96_SLICE_X101Y96_C5 = CLBLM_L_X68Y96_SLICE_X102Y96_AQ;
  assign RIOI3_X105Y85_OLOGIC_X1Y85_D1 = CLBLL_R_X71Y98_SLICE_X106Y98_AQ;
  assign CLBLM_R_X67Y96_SLICE_X101Y96_C6 = CLBLM_R_X67Y98_SLICE_X101Y98_BO6;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_B1 = CLBLM_L_X76Y134_SLICE_X116Y134_DO6;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_B2 = CLBLM_L_X76Y133_SLICE_X116Y133_BQ;
  assign RIOI3_X105Y85_OLOGIC_X1Y85_T1 = 1'b1;
  assign CLBLM_L_X76Y123_SLICE_X116Y123_B2 = CLBLM_L_X76Y123_SLICE_X116Y123_BQ;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X78Y131_SLICE_X120Y131_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X67Y96_SLICE_X101Y96_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_B4 = CLBLL_R_X75Y134_SLICE_X115Y134_AQ;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_B5 = CLBLL_R_X75Y133_SLICE_X115Y133_BQ;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_B6 = CLBLM_L_X74Y132_SLICE_X112Y132_C5Q;
  assign RIOB33_X105Y183_IOB_X1Y184_O = 1'b0;
  assign CLBLM_L_X76Y123_SLICE_X116Y123_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign RIOB33_X105Y183_IOB_X1Y183_O = 1'b0;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_C1 = 1'b1;
  assign CLBLM_L_X76Y123_SLICE_X116Y123_B4 = CLBLL_R_X75Y123_SLICE_X115Y123_AQ;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_C2 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_C3 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_C4 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_C5 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_C6 = 1'b1;
  assign CLBLM_L_X76Y123_SLICE_X116Y123_B5 = CLBLM_L_X74Y123_SLICE_X113Y123_CO5;
  assign CLBLM_L_X72Y111_SLICE_X109Y111_C6 = 1'b1;
  assign CLBLM_R_X67Y96_SLICE_X101Y96_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X72Y111_SLICE_X109Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X76Y123_SLICE_X116Y123_B6 = CLBLL_R_X75Y121_SLICE_X114Y121_BQ;
  assign RIOB33_X105Y133_IOB_X1Y134_O = CLBLL_R_X83Y130_SLICE_X130Y130_BQ;
  assign RIOB33_X105Y133_IOB_X1Y133_O = CLBLL_R_X83Y130_SLICE_X130Y130_AQ;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_D1 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_D2 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_D3 = 1'b1;
  assign CLBLM_L_X72Y111_SLICE_X109Y111_D3 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_D4 = 1'b1;
  assign CLBLM_L_X72Y111_SLICE_X109Y111_D4 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_D5 = 1'b1;
  assign CLBLM_L_X72Y111_SLICE_X109Y111_D5 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_A1 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_A2 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_A3 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_A4 = 1'b1;
  assign CLBLM_L_X72Y111_SLICE_X109Y111_D6 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_A5 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_A6 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_D6 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_B1 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_B2 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_B3 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_B4 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_B5 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_B6 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_C1 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_C2 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_C3 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_C4 = 1'b1;
  assign CLBLM_L_X72Y111_SLICE_X109Y111_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_C5 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_C6 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_D1 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_D2 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_D3 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_D4 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_D5 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_D6 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X93Y92_A1 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X93Y92_A2 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X93Y92_A3 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X93Y92_A4 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X93Y92_A5 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X93Y92_A6 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_A1 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_A2 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_A3 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X93Y92_B1 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X93Y92_B2 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X93Y92_B3 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X93Y92_B4 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X93Y92_B5 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X93Y92_B6 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_AX = CLBLM_L_X72Y116_SLICE_X108Y116_BQ;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_B1 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_B2 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X93Y92_C1 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X93Y92_C2 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X93Y92_C3 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X93Y92_C4 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X93Y92_C5 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X93Y92_C6 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_BX = CLBLM_L_X72Y118_SLICE_X108Y118_BQ;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_C1 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_C2 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_C3 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_C4 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_C5 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_C6 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_CE = CLBLM_L_X76Y109_SLICE_X116Y109_AO6;
  assign CLBLM_L_X62Y92_SLICE_X93Y92_D1 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X93Y92_D2 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X93Y92_D3 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X93Y92_D4 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X93Y92_D5 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X93Y92_D6 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_D1 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_D2 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_D3 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_D4 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_D5 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X92Y92_A1 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X92Y92_A2 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X92Y92_A3 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X92Y92_A4 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X92Y92_A5 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X92Y92_A6 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X62Y92_SLICE_X92Y92_AX = CLBLM_L_X62Y90_SLICE_X92Y90_AQ;
  assign CLBLM_L_X62Y92_SLICE_X92Y92_B1 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X92Y92_B2 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X92Y92_B3 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X92Y92_B4 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X92Y92_B5 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X92Y92_B6 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X92Y92_BX = CLBLM_L_X60Y97_SLICE_X91Y97_AQ;
  assign CLBLM_L_X62Y92_SLICE_X92Y92_C1 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X92Y92_C2 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X92Y92_C3 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X92Y92_C4 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X92Y92_C5 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X92Y92_C6 = 1'b1;
  assign CLBLM_L_X72Y111_SLICE_X108Y111_B5 = CLBLM_L_X72Y111_SLICE_X108Y111_CQ;
  assign CLBLM_L_X72Y111_SLICE_X108Y111_B6 = CLBLM_L_X70Y112_SLICE_X104Y112_CQ;
  assign CLBLM_L_X62Y92_SLICE_X92Y92_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X62Y92_SLICE_X92Y92_D1 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X92Y92_D2 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X92Y92_D3 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X92Y92_D4 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X92Y92_D5 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X92Y92_D6 = 1'b1;
  assign CLBLM_L_X62Y92_SLICE_X92Y92_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y111_SLICE_X108Y111_C3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y104_SLICE_X113Y104_C5 = 1'b1;
  assign CLBLM_L_X72Y111_SLICE_X108Y111_C5 = CLBLL_R_X71Y111_SLICE_X107Y111_CO6;
  assign CLBLM_L_X72Y111_SLICE_X108Y111_C6 = 1'b1;
  assign CLBLM_L_X72Y111_SLICE_X108Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOB33_X105Y135_IOB_X1Y136_O = CLBLL_R_X83Y130_SLICE_X130Y130_DQ;
  assign CLBLM_L_X72Y111_SLICE_X108Y111_D4 = CLBLM_L_X72Y111_SLICE_X109Y111_CQ;
  assign RIOB33_X105Y135_IOB_X1Y135_O = CLBLL_R_X83Y130_SLICE_X130Y130_CQ;
  assign CLBLM_L_X72Y111_SLICE_X108Y111_D5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_A1 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_A2 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_A3 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_A4 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_A5 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_A6 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_B1 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_B2 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_B3 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_B4 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_B5 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_B6 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_C1 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_C2 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_C3 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_C4 = 1'b1;
  assign CLBLM_L_X68Y105_SLICE_X103Y105_A1 = CLBLM_L_X68Y109_SLICE_X103Y109_BQ;
  assign CLBLM_L_X68Y105_SLICE_X103Y105_A2 = CLBLM_L_X68Y105_SLICE_X103Y105_BQ;
  assign CLBLM_L_X68Y105_SLICE_X103Y105_A3 = CLBLM_L_X68Y105_SLICE_X103Y105_AQ;
  assign CLBLM_L_X68Y105_SLICE_X103Y105_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y105_SLICE_X103Y105_A5 = CLBLM_L_X68Y109_SLICE_X103Y109_B5Q;
  assign CLBLM_L_X68Y105_SLICE_X103Y105_A6 = CLBLM_L_X68Y108_SLICE_X103Y108_CO6;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_C5 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_C6 = 1'b1;
  assign CLBLM_L_X68Y105_SLICE_X103Y105_B1 = CLBLM_L_X68Y109_SLICE_X103Y109_BQ;
  assign CLBLM_L_X68Y105_SLICE_X103Y105_B2 = CLBLM_L_X70Y106_SLICE_X104Y106_CO6;
  assign CLBLM_L_X68Y105_SLICE_X103Y105_B3 = CLBLM_L_X68Y100_SLICE_X103Y100_AO6;
  assign CLBLM_L_X68Y105_SLICE_X103Y105_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y105_SLICE_X103Y105_B5 = CLBLM_L_X68Y109_SLICE_X103Y109_B5Q;
  assign CLBLM_L_X68Y105_SLICE_X103Y105_B6 = CLBLM_L_X68Y108_SLICE_X103Y108_CO6;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_D1 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_D2 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_D3 = 1'b1;
  assign CLBLM_L_X68Y105_SLICE_X103Y105_C1 = 1'b1;
  assign CLBLM_L_X68Y105_SLICE_X103Y105_C2 = 1'b1;
  assign CLBLM_L_X68Y105_SLICE_X103Y105_C3 = 1'b1;
  assign CLBLM_L_X68Y105_SLICE_X103Y105_C4 = 1'b1;
  assign CLBLM_L_X68Y105_SLICE_X103Y105_C5 = 1'b1;
  assign CLBLM_L_X68Y105_SLICE_X103Y105_C6 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_A1 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_A2 = 1'b1;
  assign CLBLM_L_X68Y105_SLICE_X103Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_A3 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_A4 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_A5 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_A6 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_AX = CLBLM_L_X72Y118_SLICE_X108Y118_C5Q;
  assign CLBLM_L_X68Y105_SLICE_X103Y105_D1 = 1'b1;
  assign CLBLM_L_X68Y105_SLICE_X103Y105_D2 = 1'b1;
  assign CLBLM_L_X68Y105_SLICE_X103Y105_D3 = 1'b1;
  assign CLBLM_L_X68Y105_SLICE_X103Y105_D4 = 1'b1;
  assign CLBLM_L_X68Y105_SLICE_X103Y105_D5 = 1'b1;
  assign CLBLM_L_X68Y105_SLICE_X103Y105_D6 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_B1 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_B2 = 1'b1;
  assign CLBLM_L_X68Y105_SLICE_X103Y105_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_B3 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_B4 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_B5 = 1'b1;
  assign CLBLM_L_X68Y105_SLICE_X102Y105_A1 = CLBLM_R_X65Y105_SLICE_X98Y105_CQ;
  assign CLBLM_L_X68Y105_SLICE_X102Y105_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y105_SLICE_X102Y105_A3 = CLBLM_L_X70Y104_SLICE_X104Y104_BQ;
  assign CLBLM_L_X68Y105_SLICE_X102Y105_A4 = CLBLM_L_X70Y104_SLICE_X105Y104_D5Q;
  assign CLBLM_L_X68Y105_SLICE_X102Y105_A5 = CLBLM_R_X65Y106_SLICE_X99Y106_C5Q;
  assign CLBLM_L_X68Y105_SLICE_X102Y105_A6 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_C1 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_C2 = 1'b1;
  assign CLBLM_L_X68Y105_SLICE_X102Y105_AX = CLBLM_L_X68Y106_SLICE_X102Y106_AO5;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_C4 = 1'b1;
  assign CLBLM_L_X68Y105_SLICE_X102Y105_B1 = CLBLM_L_X68Y108_SLICE_X103Y108_A5Q;
  assign CLBLM_L_X68Y105_SLICE_X102Y105_B2 = CLBLM_L_X68Y105_SLICE_X102Y105_BQ;
  assign CLBLM_L_X68Y105_SLICE_X102Y105_B3 = CLBLM_L_X68Y105_SLICE_X102Y105_CQ;
  assign CLBLM_L_X68Y105_SLICE_X102Y105_B4 = CLBLM_L_X70Y106_SLICE_X104Y106_BQ;
  assign CLBLM_L_X68Y105_SLICE_X102Y105_B5 = CLBLM_L_X68Y108_SLICE_X103Y108_AQ;
  assign CLBLM_L_X68Y105_SLICE_X102Y105_B6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_D1 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_D2 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_D3 = 1'b1;
  assign CLBLM_L_X68Y105_SLICE_X102Y105_C1 = CLBLM_L_X68Y108_SLICE_X103Y108_AQ;
  assign CLBLM_L_X68Y105_SLICE_X102Y105_C2 = CLBLM_L_X68Y108_SLICE_X103Y108_A5Q;
  assign CLBLM_L_X68Y105_SLICE_X102Y105_C3 = CLBLM_L_X70Y106_SLICE_X104Y106_BQ;
  assign CLBLM_L_X68Y105_SLICE_X102Y105_C4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y105_SLICE_X102Y105_C5 = CLBLM_L_X68Y105_SLICE_X102Y105_BQ;
  assign CLBLM_L_X68Y105_SLICE_X102Y105_C6 = CLBLM_L_X68Y105_SLICE_X102Y105_CQ;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_D6 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X68Y105_SLICE_X102Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X68Y105_SLICE_X102Y105_D1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y105_SLICE_X102Y105_D2 = CLBLM_R_X67Y105_SLICE_X101Y105_CO6;
  assign CLBLM_L_X68Y105_SLICE_X102Y105_D3 = CLBLM_R_X65Y105_SLICE_X98Y105_CQ;
  assign CLBLM_L_X68Y105_SLICE_X102Y105_D4 = CLBLM_L_X68Y105_SLICE_X102Y105_AO5;
  assign CLBLM_L_X68Y105_SLICE_X102Y105_D5 = CLBLM_R_X65Y106_SLICE_X99Y106_C5Q;
  assign CLBLM_L_X68Y105_SLICE_X102Y105_D6 = CLBLM_R_X65Y105_SLICE_X99Y105_BO5;
  assign CLBLM_L_X68Y105_SLICE_X102Y105_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_A1 = CLBLM_L_X64Y105_SLICE_X96Y105_AO5;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_A3 = CLBLM_R_X63Y107_SLICE_X95Y107_AQ;
  assign LIOB33_X0Y51_IOB_X0Y52_O = CLBLM_L_X68Y95_SLICE_X102Y95_A5Q;
  assign LIOB33_X0Y51_IOB_X0Y51_O = CLBLM_L_X62Y101_SLICE_X92Y101_AQ;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_D1 = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_B4 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_T1 = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_D1 = CLBLL_L_X34Y126_SLICE_X50Y126_AO6;
  assign RIOB33_X105Y137_IOB_X1Y138_O = CLBLM_L_X82Y130_SLICE_X128Y130_AQ;
  assign RIOB33_X105Y137_IOB_X1Y137_O = CLBLL_R_X77Y125_SLICE_X118Y125_AQ;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_T1 = 1'b1;
  assign RIOI3_X105Y89_OLOGIC_X1Y90_D1 = CLBLM_L_X72Y119_SLICE_X108Y119_C5Q;
  assign CLBLM_L_X74Y104_SLICE_X113Y104_D5 = 1'b1;
  assign RIOI3_X105Y89_OLOGIC_X1Y90_T1 = 1'b1;
  assign RIOI3_X105Y89_OLOGIC_X1Y89_D1 = CLBLM_L_X64Y101_SLICE_X96Y101_AQ;
  assign RIOI3_X105Y89_OLOGIC_X1Y89_T1 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X122Y96_C4 = 1'b1;
  assign CLBLL_R_X79Y96_SLICE_X122Y96_C6 = 1'b1;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_A1 = CLBLL_R_X83Y94_SLICE_X130Y94_AQ;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_A2 = CLBLL_R_X73Y104_SLICE_X110Y104_BQ;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_A3 = CLBLM_L_X72Y118_SLICE_X109Y118_AQ;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_A5 = CLBLM_L_X72Y119_SLICE_X108Y119_AQ;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_A6 = 1'b1;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_B1 = 1'b1;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_B2 = CLBLL_R_X73Y118_SLICE_X110Y118_AQ;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_B4 = CLBLM_L_X72Y119_SLICE_X108Y119_BQ;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_B5 = CLBLL_R_X73Y118_SLICE_X110Y118_BQ;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_B6 = CLBLM_L_X72Y119_SLICE_X108Y119_A5Q;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_C1 = 1'b1;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_C2 = 1'b1;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_C3 = 1'b1;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_C4 = 1'b1;
  assign CLBLM_L_X68Y106_SLICE_X103Y106_A1 = CLBLM_L_X68Y108_SLICE_X103Y108_A5Q;
  assign CLBLM_L_X68Y106_SLICE_X103Y106_A2 = CLBLM_L_X70Y106_SLICE_X104Y106_BQ;
  assign CLBLM_L_X68Y106_SLICE_X103Y106_A3 = CLBLM_L_X68Y106_SLICE_X103Y106_CQ;
  assign CLBLM_L_X68Y106_SLICE_X103Y106_A4 = CLBLM_L_X68Y108_SLICE_X103Y108_AQ;
  assign CLBLM_L_X68Y106_SLICE_X103Y106_A5 = CLBLM_L_X68Y105_SLICE_X102Y105_CQ;
  assign CLBLM_L_X68Y106_SLICE_X103Y106_A6 = 1'b1;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_C5 = 1'b1;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_C6 = 1'b1;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X68Y106_SLICE_X103Y106_B1 = CLBLM_L_X68Y106_SLICE_X103Y106_B5Q;
  assign CLBLM_L_X68Y106_SLICE_X103Y106_B2 = CLBLM_L_X68Y106_SLICE_X103Y106_BQ;
  assign CLBLM_L_X68Y106_SLICE_X103Y106_B3 = CLBLM_L_X68Y106_SLICE_X103Y106_CQ;
  assign CLBLM_L_X68Y106_SLICE_X103Y106_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y106_SLICE_X103Y106_B5 = CLBLM_L_X68Y106_SLICE_X103Y106_AO5;
  assign CLBLM_L_X68Y106_SLICE_X103Y106_B6 = 1'b1;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_D1 = 1'b1;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_D2 = 1'b1;
  assign CLBLM_L_X68Y106_SLICE_X103Y106_C1 = CLBLM_L_X68Y108_SLICE_X103Y108_AQ;
  assign CLBLM_L_X68Y106_SLICE_X103Y106_C2 = CLBLM_L_X70Y106_SLICE_X104Y106_BQ;
  assign CLBLM_L_X68Y106_SLICE_X103Y106_C3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y106_SLICE_X103Y106_C4 = CLBLM_L_X68Y108_SLICE_X103Y108_A5Q;
  assign CLBLM_L_X68Y106_SLICE_X103Y106_C5 = CLBLM_L_X68Y106_SLICE_X103Y106_CQ;
  assign CLBLM_L_X68Y106_SLICE_X103Y106_C6 = CLBLM_L_X68Y105_SLICE_X102Y105_CQ;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_A1 = CLBLM_L_X72Y121_SLICE_X109Y121_A5Q;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_A2 = CLBLM_L_X72Y118_SLICE_X108Y118_DQ;
  assign CLBLM_L_X68Y106_SLICE_X103Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_A3 = CLBLM_L_X72Y118_SLICE_X108Y118_AQ;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_A4 = CLBLM_L_X74Y119_SLICE_X112Y119_AQ;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_A6 = 1'b1;
  assign CLBLM_L_X68Y106_SLICE_X103Y106_D1 = CLBLM_L_X68Y108_SLICE_X103Y108_AQ;
  assign CLBLM_L_X68Y106_SLICE_X103Y106_D2 = CLBLM_L_X68Y106_SLICE_X103Y106_CQ;
  assign CLBLM_L_X68Y106_SLICE_X103Y106_D3 = CLBLM_L_X68Y106_SLICE_X103Y106_BQ;
  assign CLBLM_L_X68Y106_SLICE_X103Y106_D4 = CLBLM_L_X68Y108_SLICE_X103Y108_A5Q;
  assign CLBLM_L_X68Y106_SLICE_X103Y106_D5 = CLBLM_L_X68Y106_SLICE_X103Y106_B5Q;
  assign CLBLM_L_X68Y106_SLICE_X103Y106_D6 = CLBLM_L_X68Y105_SLICE_X102Y105_CQ;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_B1 = CLBLM_L_X72Y118_SLICE_X108Y118_B5Q;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_B2 = CLBLM_L_X72Y118_SLICE_X108Y118_BQ;
  assign CLBLL_R_X79Y96_SLICE_X122Y96_D5 = 1'b1;
  assign CLBLM_L_X68Y106_SLICE_X103Y106_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_B3 = CLBLM_L_X72Y118_SLICE_X108Y118_DQ;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y106_SLICE_X102Y106_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y106_SLICE_X102Y106_A2 = CLBLM_L_X64Y104_SLICE_X96Y104_CQ;
  assign CLBLM_L_X68Y106_SLICE_X102Y106_A3 = CLBLM_L_X70Y104_SLICE_X105Y104_BQ;
  assign CLBLM_L_X68Y106_SLICE_X102Y106_A4 = CLBLM_R_X65Y100_SLICE_X98Y100_AQ;
  assign CLBLM_L_X68Y106_SLICE_X102Y106_A5 = CLBLM_L_X64Y105_SLICE_X96Y105_C5Q;
  assign CLBLL_R_X79Y96_SLICE_X122Y96_D6 = 1'b1;
  assign CLBLM_L_X68Y106_SLICE_X102Y106_A6 = 1'b1;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_C1 = CLBLM_L_X72Y118_SLICE_X108Y118_C5Q;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_C2 = 1'b1;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_C4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y106_SLICE_X102Y106_B1 = CLBLM_L_X68Y107_SLICE_X102Y107_AO5;
  assign CLBLM_L_X68Y106_SLICE_X102Y106_B2 = CLBLM_L_X64Y104_SLICE_X96Y104_CQ;
  assign CLBLM_L_X68Y106_SLICE_X102Y106_B3 = CLBLM_L_X68Y106_SLICE_X102Y106_DO6;
  assign CLBLM_L_X68Y106_SLICE_X102Y106_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y106_SLICE_X102Y106_B5 = CLBLM_L_X68Y102_SLICE_X102Y102_CQ;
  assign CLBLM_L_X68Y106_SLICE_X102Y106_B6 = CLBLM_L_X68Y106_SLICE_X102Y106_CO6;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_D1 = CLBLM_L_X72Y117_SLICE_X108Y117_BQ;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_D2 = CLBLM_L_X70Y104_SLICE_X104Y104_A5Q;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_D3 = CLBLM_L_X74Y118_SLICE_X112Y118_CQ;
  assign CLBLM_L_X68Y106_SLICE_X102Y106_C1 = CLBLM_R_X65Y100_SLICE_X98Y100_AQ;
  assign CLBLM_L_X68Y106_SLICE_X102Y106_C2 = CLBLL_R_X71Y108_SLICE_X106Y108_BQ;
  assign CLBLM_L_X68Y106_SLICE_X102Y106_C3 = CLBLM_L_X72Y105_SLICE_X108Y105_CQ;
  assign CLBLM_L_X68Y106_SLICE_X102Y106_C4 = CLBLM_R_X67Y109_SLICE_X100Y109_BQ;
  assign CLBLM_L_X68Y106_SLICE_X102Y106_C5 = CLBLM_L_X70Y104_SLICE_X105Y104_BQ;
  assign CLBLM_L_X68Y106_SLICE_X102Y106_C6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_D6 = 1'b1;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X82Y130_SLICE_X129Y130_A4 = 1'b1;
  assign CLBLM_L_X68Y106_SLICE_X102Y106_D1 = CLBLM_L_X64Y104_SLICE_X96Y104_CQ;
  assign CLBLM_L_X68Y106_SLICE_X102Y106_D2 = CLBLM_R_X67Y109_SLICE_X100Y109_BQ;
  assign CLBLM_L_X68Y106_SLICE_X102Y106_D3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y106_SLICE_X102Y106_D4 = CLBLM_L_X68Y102_SLICE_X102Y102_CQ;
  assign CLBLM_L_X68Y106_SLICE_X102Y106_D5 = CLBLM_L_X70Y104_SLICE_X105Y104_BQ;
  assign CLBLM_L_X68Y106_SLICE_X102Y106_D6 = CLBLM_R_X65Y100_SLICE_X98Y100_AQ;
  assign CLBLM_L_X76Y119_SLICE_X116Y119_A6 = 1'b1;
  assign CLBLM_L_X82Y130_SLICE_X129Y130_A5 = 1'b1;
  assign LIOB33_X0Y53_IOB_X0Y54_O = CLBLM_L_X62Y92_SLICE_X92Y92_AQ;
  assign LIOB33_X0Y53_IOB_X0Y53_O = CLBLM_L_X62Y90_SLICE_X92Y90_AQ;
  assign CLBLM_L_X82Y130_SLICE_X129Y130_A6 = 1'b1;
  assign RIOB33_X105Y139_IOB_X1Y140_O = CLBLM_L_X72Y107_SLICE_X109Y107_A5Q;
  assign RIOB33_X105Y139_IOB_X1Y139_O = CLBLL_R_X83Y132_SLICE_X130Y132_AQ;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_D1 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_B2 = 1'b1;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_C3 = CLBLL_R_X75Y128_SLICE_X115Y128_DO6;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_C5 = CLBLM_L_X74Y127_SLICE_X113Y127_BO5;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_C6 = CLBLL_R_X75Y128_SLICE_X114Y128_DO6;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1 = 1'b1;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_T1 = 1'b1;
  assign CLBLM_L_X82Y130_SLICE_X129Y130_B2 = 1'b1;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_A1 = CLBLL_R_X73Y119_SLICE_X110Y119_CO6;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_A3 = CLBLM_L_X72Y119_SLICE_X109Y119_AQ;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_A4 = CLBLM_L_X72Y119_SLICE_X109Y119_DO6;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_A5 = CLBLL_R_X73Y118_SLICE_X110Y118_AQ;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_A6 = CLBLM_L_X72Y113_SLICE_X108Y113_AQ;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_D6 = 1'b1;
  assign CLBLM_L_X76Y119_SLICE_X116Y119_B3 = 1'b1;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_AX = CLBLM_L_X72Y119_SLICE_X108Y119_CQ;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_B1 = CLBLM_L_X70Y119_SLICE_X105Y119_A5Q;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_B2 = CLBLL_R_X73Y118_SLICE_X111Y118_A5Q;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_B3 = CLBLM_L_X72Y119_SLICE_X109Y119_AQ;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_B5 = CLBLM_L_X72Y119_SLICE_X109Y119_CO6;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_B6 = CLBLM_L_X72Y119_SLICE_X109Y119_A5Q;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_BX = CLBLM_L_X72Y119_SLICE_X109Y119_BQ;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_C1 = CLBLM_L_X72Y119_SLICE_X109Y119_A5Q;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_C2 = CLBLM_L_X70Y119_SLICE_X105Y119_A5Q;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_C3 = CLBLM_L_X72Y119_SLICE_X109Y119_BQ;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_C4 = CLBLM_L_X72Y119_SLICE_X108Y119_CQ;
  assign CLBLM_L_X68Y107_SLICE_X103Y107_A1 = CLBLM_L_X64Y104_SLICE_X96Y104_CQ;
  assign CLBLM_L_X68Y107_SLICE_X103Y107_A2 = CLBLM_L_X70Y108_SLICE_X105Y108_AO6;
  assign CLBLM_L_X68Y107_SLICE_X103Y107_A3 = CLBLM_L_X70Y104_SLICE_X105Y104_BQ;
  assign CLBLM_L_X68Y107_SLICE_X103Y107_A4 = CLBLM_L_X68Y107_SLICE_X102Y107_AO6;
  assign CLBLM_L_X68Y107_SLICE_X103Y107_A5 = CLBLM_R_X65Y100_SLICE_X98Y100_AQ;
  assign CLBLM_L_X68Y107_SLICE_X103Y107_A6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_C5 = CLBLM_L_X72Y119_SLICE_X109Y119_B5Q;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_C6 = 1'b1;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X68Y107_SLICE_X103Y107_B1 = CLBLM_L_X68Y107_SLICE_X102Y107_CO6;
  assign CLBLM_L_X68Y107_SLICE_X103Y107_B2 = CLBLL_R_X71Y108_SLICE_X106Y108_BQ;
  assign CLBLM_L_X68Y107_SLICE_X103Y107_B3 = CLBLM_L_X70Y104_SLICE_X105Y104_BQ;
  assign CLBLM_L_X68Y107_SLICE_X103Y107_B4 = CLBLM_R_X67Y109_SLICE_X100Y109_BQ;
  assign CLBLM_L_X68Y107_SLICE_X103Y107_B5 = CLBLM_L_X68Y107_SLICE_X103Y107_CO6;
  assign CLBLM_L_X68Y107_SLICE_X103Y107_B6 = CLBLM_R_X65Y106_SLICE_X98Y106_CQ;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_D1 = 1'b1;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_D2 = CLBLL_R_X73Y118_SLICE_X111Y118_A5Q;
  assign CLBLM_L_X68Y107_SLICE_X103Y107_C1 = CLBLM_L_X68Y102_SLICE_X102Y102_CQ;
  assign CLBLM_L_X68Y107_SLICE_X103Y107_C2 = CLBLM_L_X72Y105_SLICE_X108Y105_CQ;
  assign CLBLM_L_X68Y107_SLICE_X103Y107_C3 = CLBLM_L_X64Y104_SLICE_X96Y104_CQ;
  assign CLBLM_L_X68Y107_SLICE_X103Y107_C4 = CLBLM_L_X74Y109_SLICE_X113Y109_A5Q;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_A1 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_A2 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_A3 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_A4 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_A5 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_A6 = 1'b1;
  assign CLBLM_L_X68Y107_SLICE_X103Y107_C5 = CLBLM_R_X65Y100_SLICE_X98Y100_AQ;
  assign CLBLM_L_X68Y107_SLICE_X103Y107_C6 = CLBLM_L_X72Y118_SLICE_X109Y118_BQ;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_B1 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_B2 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_B3 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_B4 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_B5 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_B6 = 1'b1;
  assign CLBLM_L_X68Y107_SLICE_X103Y107_D1 = CLBLM_L_X68Y106_SLICE_X103Y106_CQ;
  assign CLBLM_L_X68Y107_SLICE_X103Y107_D2 = CLBLM_L_X70Y106_SLICE_X104Y106_BO6;
  assign CLBLM_L_X68Y107_SLICE_X103Y107_D3 = CLBLM_L_X68Y106_SLICE_X103Y106_B5Q;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_C1 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_C2 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_C3 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_C4 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_C5 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_C6 = 1'b1;
  assign CLBLM_L_X68Y107_SLICE_X102Y107_A1 = CLBLM_L_X72Y105_SLICE_X108Y105_CQ;
  assign CLBLM_L_X68Y107_SLICE_X102Y107_A2 = CLBLM_R_X67Y109_SLICE_X100Y109_BQ;
  assign CLBLM_L_X68Y107_SLICE_X102Y107_A3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y107_SLICE_X102Y107_A4 = CLBLL_R_X71Y108_SLICE_X106Y108_BQ;
  assign CLBLM_L_X68Y107_SLICE_X102Y107_A5 = CLBLM_L_X68Y102_SLICE_X102Y102_CQ;
  assign CLBLM_L_X68Y107_SLICE_X102Y107_A6 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_D1 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_D2 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_D3 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_D4 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_D5 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_D6 = 1'b1;
  assign CLBLM_L_X68Y107_SLICE_X102Y107_B1 = CLBLM_L_X72Y118_SLICE_X109Y118_BQ;
  assign CLBLM_L_X68Y107_SLICE_X102Y107_B2 = CLBLM_L_X68Y107_SLICE_X103Y107_BO6;
  assign CLBLM_L_X68Y107_SLICE_X102Y107_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y107_SLICE_X102Y107_B4 = CLBLM_R_X65Y106_SLICE_X98Y106_CQ;
  assign CLBLM_L_X68Y107_SLICE_X102Y107_B5 = CLBLM_L_X68Y106_SLICE_X102Y106_BO6;
  assign CLBLM_L_X68Y107_SLICE_X102Y107_B6 = CLBLM_L_X74Y109_SLICE_X113Y109_A5Q;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_A1 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_A2 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_A3 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_A4 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_A5 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_A6 = 1'b1;
  assign CLBLM_L_X68Y107_SLICE_X102Y107_C1 = CLBLM_L_X68Y106_SLICE_X102Y106_AO6;
  assign CLBLM_L_X68Y107_SLICE_X102Y107_C2 = CLBLM_L_X72Y118_SLICE_X109Y118_BQ;
  assign CLBLM_L_X68Y107_SLICE_X102Y107_C3 = CLBLM_L_X74Y109_SLICE_X113Y109_A5Q;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_AX = CLBLL_R_X73Y103_SLICE_X111Y103_A5Q;
  assign CLBLM_L_X68Y107_SLICE_X102Y107_C4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_B1 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_B2 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_B3 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_B4 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_B5 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_B6 = 1'b1;
  assign CLBLM_L_X68Y107_SLICE_X102Y107_D1 = CLBLM_L_X68Y102_SLICE_X102Y102_CQ;
  assign CLBLM_L_X68Y107_SLICE_X102Y107_D2 = CLBLM_R_X67Y109_SLICE_X100Y109_BQ;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_BX = CLBLM_L_X68Y95_SLICE_X102Y95_A5Q;
  assign CLBLM_L_X68Y107_SLICE_X102Y107_D3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_C1 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_C2 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_C3 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_C4 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_C5 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_C6 = 1'b1;
  assign CLBLM_L_X68Y107_SLICE_X102Y107_D6 = CLBLL_R_X71Y108_SLICE_X106Y108_BQ;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_B6 = CLBLM_L_X72Y127_SLICE_X108Y127_A5Q;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign LIOB33_X0Y55_IOB_X0Y55_O = CLBLM_L_X60Y97_SLICE_X91Y97_AQ;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_CX = CLBLM_L_X60Y97_SLICE_X90Y97_DQ;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_D1 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_D2 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_D3 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_D4 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_D5 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_D6 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X73Y101_SLICE_X110Y101_A1 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLL_R_X73Y101_SLICE_X110Y101_A2 = CLBLM_L_X72Y103_SLICE_X108Y103_CO6;
  assign CLBLL_R_X73Y101_SLICE_X110Y101_A3 = CLBLL_R_X73Y101_SLICE_X110Y101_AQ;
  assign CLBLL_R_X73Y101_SLICE_X110Y101_A4 = CLBLL_R_X73Y103_SLICE_X110Y103_BQ;
  assign CLBLL_R_X73Y101_SLICE_X110Y101_A5 = CLBLM_L_X72Y103_SLICE_X108Y103_DO6;
  assign CLBLL_R_X73Y101_SLICE_X110Y101_A6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y101_SLICE_X110Y101_B1 = 1'b1;
  assign CLBLL_R_X73Y101_SLICE_X110Y101_B2 = 1'b1;
  assign CLBLL_R_X73Y101_SLICE_X110Y101_B3 = 1'b1;
  assign CLBLL_R_X73Y101_SLICE_X110Y101_B4 = 1'b1;
  assign CLBLL_R_X73Y101_SLICE_X110Y101_B5 = 1'b1;
  assign CLBLL_R_X73Y101_SLICE_X110Y101_B6 = 1'b1;
  assign RIOB33_X105Y89_IOB_X1Y90_O = CLBLM_L_X72Y119_SLICE_X108Y119_C5Q;
  assign RIOB33_X105Y141_IOB_X1Y141_O = CLBLM_R_X65Y110_SLICE_X99Y110_AQ;
  assign RIOB33_X105Y141_IOB_X1Y142_O = CLBLL_R_X73Y103_SLICE_X110Y103_A5Q;
  assign CLBLL_R_X73Y101_SLICE_X110Y101_C1 = 1'b1;
  assign CLBLL_R_X73Y101_SLICE_X110Y101_C2 = 1'b1;
  assign CLBLL_R_X73Y101_SLICE_X110Y101_C3 = 1'b1;
  assign CLBLL_R_X73Y101_SLICE_X110Y101_C4 = 1'b1;
  assign CLBLL_R_X73Y101_SLICE_X110Y101_C5 = 1'b1;
  assign CLBLL_R_X73Y101_SLICE_X110Y101_C6 = 1'b1;
  assign RIOB33_X105Y89_IOB_X1Y89_O = CLBLM_L_X64Y101_SLICE_X96Y101_AQ;
  assign CLBLL_R_X73Y101_SLICE_X110Y101_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_CE = CLBLM_L_X76Y109_SLICE_X116Y109_AO6;
  assign CLBLL_R_X73Y101_SLICE_X110Y101_D1 = 1'b1;
  assign CLBLL_R_X73Y101_SLICE_X110Y101_D2 = 1'b1;
  assign CLBLL_R_X73Y101_SLICE_X110Y101_D3 = 1'b1;
  assign CLBLL_R_X73Y101_SLICE_X110Y101_D4 = 1'b1;
  assign CLBLL_R_X73Y101_SLICE_X110Y101_D5 = 1'b1;
  assign CLBLL_R_X73Y101_SLICE_X110Y101_D6 = 1'b1;
  assign CLBLL_R_X73Y101_SLICE_X110Y101_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X73Y101_SLICE_X111Y101_A1 = 1'b1;
  assign CLBLL_R_X73Y101_SLICE_X111Y101_A2 = 1'b1;
  assign CLBLL_R_X73Y101_SLICE_X111Y101_A3 = 1'b1;
  assign CLBLL_R_X73Y101_SLICE_X111Y101_A4 = 1'b1;
  assign CLBLL_R_X73Y101_SLICE_X111Y101_A5 = 1'b1;
  assign CLBLL_R_X73Y101_SLICE_X111Y101_A6 = 1'b1;
  assign CLBLM_L_X76Y119_SLICE_X116Y119_C1 = 1'b1;
  assign CLBLL_R_X73Y101_SLICE_X111Y101_B1 = 1'b1;
  assign CLBLL_R_X73Y101_SLICE_X111Y101_B2 = 1'b1;
  assign CLBLL_R_X73Y101_SLICE_X111Y101_B3 = 1'b1;
  assign CLBLL_R_X73Y101_SLICE_X111Y101_B4 = 1'b1;
  assign CLBLL_R_X73Y101_SLICE_X111Y101_B5 = 1'b1;
  assign CLBLL_R_X73Y101_SLICE_X111Y101_B6 = 1'b1;
  assign CLBLM_L_X76Y134_SLICE_X117Y134_B1 = CLBLM_L_X76Y134_SLICE_X116Y134_CO6;
  assign CLBLL_R_X73Y101_SLICE_X111Y101_C1 = 1'b1;
  assign CLBLL_R_X73Y101_SLICE_X111Y101_C2 = 1'b1;
  assign CLBLL_R_X73Y101_SLICE_X111Y101_C3 = 1'b1;
  assign CLBLL_R_X73Y101_SLICE_X111Y101_C4 = 1'b1;
  assign CLBLL_R_X73Y101_SLICE_X111Y101_C5 = 1'b1;
  assign CLBLL_R_X73Y101_SLICE_X111Y101_C6 = 1'b1;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_D2 = CLBLM_L_X72Y127_SLICE_X108Y127_A5Q;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_D3 = 1'b1;
  assign CLBLM_L_X76Y134_SLICE_X117Y134_B2 = CLBLM_L_X76Y134_SLICE_X117Y134_BQ;
  assign CLBLM_L_X76Y134_SLICE_X117Y134_B3 = CLBLM_L_X76Y134_SLICE_X117Y134_AQ;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_D4 = CLBLM_L_X74Y127_SLICE_X113Y127_CQ;
  assign CLBLM_L_X76Y134_SLICE_X117Y134_B4 = 1'b1;
  assign CLBLM_L_X76Y119_SLICE_X116Y119_C2 = 1'b1;
  assign CLBLL_R_X73Y101_SLICE_X111Y101_D1 = 1'b1;
  assign CLBLL_R_X73Y101_SLICE_X111Y101_D2 = 1'b1;
  assign CLBLL_R_X73Y101_SLICE_X111Y101_D3 = 1'b1;
  assign CLBLL_R_X73Y101_SLICE_X111Y101_D4 = 1'b1;
  assign CLBLL_R_X73Y101_SLICE_X111Y101_D5 = 1'b1;
  assign CLBLL_R_X73Y101_SLICE_X111Y101_D6 = 1'b1;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_D5 = CLBLM_L_X72Y128_SLICE_X108Y128_A5Q;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_D6 = CLBLM_L_X74Y128_SLICE_X112Y128_AQ;
  assign CLBLM_L_X76Y134_SLICE_X117Y134_B6 = CLBLM_L_X76Y134_SLICE_X117Y134_CO6;
  assign CLBLM_L_X76Y119_SLICE_X116Y119_C3 = 1'b1;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X76Y134_SLICE_X117Y134_C1 = CLBLL_R_X75Y134_SLICE_X114Y134_A5Q;
  assign CLBLM_L_X76Y134_SLICE_X117Y134_C2 = CLBLL_R_X75Y134_SLICE_X115Y134_AO6;
  assign CLBLM_L_X76Y134_SLICE_X117Y134_C3 = CLBLM_L_X76Y134_SLICE_X117Y134_AQ;
  assign CLBLM_L_X76Y119_SLICE_X116Y119_C4 = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_D1 = 1'b1;
  assign CLBLM_L_X76Y134_SLICE_X117Y134_C6 = CLBLL_R_X75Y133_SLICE_X115Y133_AQ;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_A1 = 1'b1;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_A2 = 1'b1;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_A3 = 1'b1;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_A4 = 1'b1;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_A5 = 1'b1;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_A6 = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_T1 = 1'b1;
  assign CLBLM_L_X76Y134_SLICE_X117Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_B1 = 1'b1;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_B2 = 1'b1;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_B3 = 1'b1;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_B4 = 1'b1;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_B5 = 1'b1;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_B6 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X114Y113_A1 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X114Y113_A2 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X114Y113_A3 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X114Y113_A4 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X114Y113_A5 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X114Y113_A6 = 1'b1;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_C1 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X114Y113_AX = CLBLM_L_X74Y109_SLICE_X113Y109_AQ;
  assign CLBLM_L_X68Y108_SLICE_X103Y108_A1 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X114Y113_B1 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X114Y113_B2 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X114Y113_B3 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X114Y113_B4 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X114Y113_B5 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X114Y113_B6 = 1'b1;
  assign CLBLM_L_X68Y108_SLICE_X103Y108_A2 = CLBLM_L_X68Y108_SLICE_X103Y108_A5Q;
  assign CLBLM_L_X68Y108_SLICE_X103Y108_A3 = CLBLM_L_X68Y108_SLICE_X103Y108_AQ;
  assign CLBLM_L_X68Y108_SLICE_X103Y108_A4 = CLBLM_L_X70Y106_SLICE_X104Y106_BQ;
  assign CLBLL_R_X75Y113_SLICE_X114Y113_C1 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X114Y113_C2 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X114Y113_C3 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X114Y113_C4 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X114Y113_C5 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X114Y113_C6 = 1'b1;
  assign CLBLM_L_X68Y108_SLICE_X103Y108_B1 = CLBLM_L_X68Y109_SLICE_X103Y109_B5Q;
  assign CLBLM_L_X68Y108_SLICE_X103Y108_B2 = CLBLM_L_X68Y109_SLICE_X103Y109_BQ;
  assign CLBLL_R_X75Y113_SLICE_X114Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X68Y108_SLICE_X103Y108_B3 = CLBLM_L_X68Y108_SLICE_X102Y108_CO6;
  assign CLBLM_L_X68Y108_SLICE_X103Y108_B4 = CLBLM_L_X70Y106_SLICE_X105Y106_DO6;
  assign CLBLM_L_X68Y108_SLICE_X103Y108_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y108_SLICE_X103Y108_B6 = CLBLM_L_X68Y108_SLICE_X103Y108_CO6;
  assign CLBLL_R_X75Y113_SLICE_X114Y113_D1 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X114Y113_D2 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X114Y113_D3 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X114Y113_D4 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X114Y113_D5 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X114Y113_D6 = 1'b1;
  assign CLBLM_L_X68Y108_SLICE_X103Y108_C5 = 1'b1;
  assign CLBLM_L_X68Y108_SLICE_X103Y108_C6 = CLBLM_L_X68Y106_SLICE_X103Y106_CQ;
  assign CLBLL_R_X75Y113_SLICE_X114Y113_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X68Y108_SLICE_X103Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X68Y108_SLICE_X103Y108_D1 = 1'b1;
  assign CLBLM_L_X68Y108_SLICE_X103Y108_D2 = 1'b1;
  assign CLBLM_L_X68Y108_SLICE_X103Y108_D3 = 1'b1;
  assign CLBLM_L_X68Y108_SLICE_X103Y108_D4 = 1'b1;
  assign CLBLM_L_X68Y108_SLICE_X103Y108_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X68Y108_SLICE_X103Y108_D5 = 1'b1;
  assign CLBLM_L_X68Y108_SLICE_X103Y108_D6 = 1'b1;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_B4 = 1'b1;
  assign CLBLM_L_X68Y108_SLICE_X102Y108_A1 = CLBLM_L_X68Y108_SLICE_X102Y108_B5Q;
  assign CLBLM_L_X68Y108_SLICE_X102Y108_A2 = CLBLM_L_X68Y108_SLICE_X102Y108_A5Q;
  assign CLBLM_L_X68Y108_SLICE_X102Y108_A3 = CLBLM_L_X68Y108_SLICE_X102Y108_AQ;
  assign CLBLM_L_X68Y108_SLICE_X102Y108_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y108_SLICE_X102Y108_A5 = CLBLM_L_X70Y106_SLICE_X105Y106_DO6;
  assign CLBLM_L_X68Y108_SLICE_X102Y108_A6 = 1'b1;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_C1 = 1'b1;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_C2 = 1'b1;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_C3 = 1'b1;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_C4 = 1'b1;
  assign CLBLM_L_X68Y108_SLICE_X102Y108_B1 = CLBLM_L_X68Y108_SLICE_X102Y108_B5Q;
  assign CLBLM_L_X68Y108_SLICE_X102Y108_B2 = CLBLM_L_X68Y108_SLICE_X102Y108_BQ;
  assign CLBLM_L_X68Y108_SLICE_X102Y108_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y113_SLICE_X115Y113_A1 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X115Y113_A2 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X115Y113_A3 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X115Y113_A4 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X115Y113_A5 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X115Y113_A6 = 1'b1;
  assign CLBLM_L_X68Y108_SLICE_X102Y108_B4 = CLBLM_L_X68Y109_SLICE_X102Y109_A5Q;
  assign CLBLM_L_X68Y108_SLICE_X102Y108_B5 = CLBLM_R_X67Y109_SLICE_X100Y109_DO5;
  assign CLBLM_L_X68Y108_SLICE_X102Y108_B6 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X115Y113_B1 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X115Y113_B2 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X115Y113_B3 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X115Y113_B4 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X115Y113_B5 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X115Y113_B6 = 1'b1;
  assign CLBLM_L_X68Y108_SLICE_X102Y108_C1 = CLBLM_L_X70Y106_SLICE_X105Y106_DO6;
  assign CLBLM_L_X68Y108_SLICE_X102Y108_C2 = CLBLM_L_X68Y108_SLICE_X102Y108_AQ;
  assign CLBLM_L_X68Y108_SLICE_X102Y108_C3 = CLBLM_L_X68Y108_SLICE_X102Y108_BQ;
  assign CLBLL_R_X75Y113_SLICE_X115Y113_C1 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X115Y113_C2 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X115Y113_C3 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X115Y113_C4 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X115Y113_C5 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X115Y113_C6 = 1'b1;
  assign CLBLM_L_X68Y108_SLICE_X102Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X68Y108_SLICE_X102Y108_D1 = 1'b1;
  assign CLBLM_L_X68Y108_SLICE_X102Y108_D2 = 1'b1;
  assign CLBLM_L_X68Y108_SLICE_X102Y108_D3 = 1'b1;
  assign CLBLM_L_X68Y108_SLICE_X102Y108_D4 = 1'b1;
  assign CLBLM_L_X68Y108_SLICE_X102Y108_D5 = 1'b1;
  assign CLBLM_L_X68Y108_SLICE_X102Y108_D6 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X115Y113_D1 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X115Y113_D2 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X115Y113_D3 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X115Y113_D4 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X115Y113_D5 = 1'b1;
  assign CLBLL_R_X75Y113_SLICE_X115Y113_D6 = 1'b1;
  assign CLBLM_L_X68Y108_SLICE_X102Y108_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X76Y134_SLICE_X116Y134_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X76Y134_SLICE_X116Y134_A5 = CLBLM_L_X76Y133_SLICE_X116Y133_AQ;
  assign CLBLM_L_X76Y134_SLICE_X116Y134_A6 = CLBLL_R_X75Y134_SLICE_X115Y134_AQ;
  assign RIOB33_X105Y143_IOB_X1Y143_O = CLBLM_L_X62Y106_SLICE_X92Y106_BQ;
  assign CLBLM_R_X67Y97_SLICE_X101Y97_C1 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign RIOB33_X105Y143_IOB_X1Y144_O = CLBLM_L_X70Y101_SLICE_X105Y101_AQ;
  assign CLBLM_R_X67Y97_SLICE_X101Y97_C2 = CLBLM_R_X67Y97_SLICE_X101Y97_CQ;
  assign CLBLL_R_X73Y102_SLICE_X110Y102_A1 = CLBLL_R_X73Y102_SLICE_X110Y102_CQ;
  assign CLBLL_R_X73Y102_SLICE_X110Y102_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y102_SLICE_X110Y102_A3 = CLBLL_R_X73Y102_SLICE_X110Y102_AQ;
  assign CLBLL_R_X73Y102_SLICE_X110Y102_A4 = CLBLM_L_X72Y103_SLICE_X108Y103_A5Q;
  assign CLBLL_R_X73Y102_SLICE_X110Y102_A5 = CLBLM_L_X72Y103_SLICE_X108Y103_CO5;
  assign CLBLL_R_X73Y102_SLICE_X110Y102_A6 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X67Y97_SLICE_X101Y97_C3 = CLBLM_R_X67Y98_SLICE_X101Y98_AO5;
  assign CLBLL_R_X73Y102_SLICE_X110Y102_AX = CLBLL_R_X73Y102_SLICE_X111Y102_A5Q;
  assign CLBLM_R_X67Y97_SLICE_X101Y97_C4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y102_SLICE_X110Y102_B1 = CLBLM_L_X72Y103_SLICE_X108Y103_CO5;
  assign CLBLL_R_X73Y102_SLICE_X110Y102_B2 = CLBLL_R_X73Y102_SLICE_X110Y102_BQ;
  assign CLBLL_R_X73Y102_SLICE_X110Y102_B3 = CLBLM_L_X72Y103_SLICE_X108Y103_DO6;
  assign CLBLL_R_X73Y102_SLICE_X110Y102_B4 = CLBLM_L_X72Y103_SLICE_X109Y103_BQ;
  assign CLBLL_R_X73Y102_SLICE_X110Y102_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y102_SLICE_X110Y102_B6 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X67Y97_SLICE_X101Y97_C5 = CLBLM_R_X67Y97_SLICE_X101Y97_AQ;
  assign CLBLM_R_X67Y97_SLICE_X101Y97_C6 = CLBLM_R_X67Y98_SLICE_X101Y98_CO6;
  assign CLBLL_R_X73Y102_SLICE_X110Y102_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y102_SLICE_X110Y102_C2 = CLBLL_R_X73Y102_SLICE_X110Y102_CQ;
  assign CLBLL_R_X73Y102_SLICE_X110Y102_C3 = CLBLM_L_X72Y103_SLICE_X108Y103_CO5;
  assign CLBLL_R_X73Y102_SLICE_X110Y102_C4 = CLBLL_R_X73Y102_SLICE_X110Y102_BQ;
  assign CLBLL_R_X73Y102_SLICE_X110Y102_C5 = CLBLM_L_X72Y103_SLICE_X108Y103_DO5;
  assign CLBLL_R_X73Y102_SLICE_X110Y102_C6 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X76Y134_SLICE_X116Y134_B1 = CLBLM_L_X76Y134_SLICE_X116Y134_AQ;
  assign CLBLM_L_X76Y134_SLICE_X116Y134_B2 = CLBLM_L_X76Y134_SLICE_X116Y134_BQ;
  assign CLBLL_R_X73Y102_SLICE_X110Y102_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X76Y134_SLICE_X116Y134_B3 = CLBLM_L_X76Y134_SLICE_X117Y134_CO6;
  assign CLBLM_R_X67Y97_SLICE_X101Y97_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLL_R_X73Y102_SLICE_X110Y102_D1 = 1'b1;
  assign CLBLL_R_X73Y102_SLICE_X110Y102_D2 = CLBLL_R_X73Y102_SLICE_X111Y102_A5Q;
  assign CLBLL_R_X73Y102_SLICE_X110Y102_D3 = CLBLM_L_X72Y104_SLICE_X109Y104_BQ;
  assign CLBLL_R_X73Y102_SLICE_X110Y102_D4 = CLBLL_R_X73Y104_SLICE_X110Y104_A5Q;
  assign CLBLL_R_X73Y102_SLICE_X110Y102_D5 = CLBLL_R_X73Y102_SLICE_X110Y102_CQ;
  assign CLBLL_R_X73Y102_SLICE_X110Y102_D6 = CLBLM_L_X72Y104_SLICE_X109Y104_B5Q;
  assign CLBLM_L_X76Y134_SLICE_X116Y134_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y102_SLICE_X110Y102_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X76Y134_SLICE_X116Y134_B5 = CLBLL_R_X75Y134_SLICE_X115Y134_DO5;
  assign CLBLM_R_X67Y97_SLICE_X100Y97_B6 = 1'b1;
  assign CLBLM_L_X76Y134_SLICE_X116Y134_B6 = CLBLM_L_X76Y133_SLICE_X116Y133_AQ;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_B2 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_B3 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_B5 = 1'b1;
  assign CLBLL_R_X73Y102_SLICE_X111Y102_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y102_SLICE_X111Y102_A2 = CLBLM_L_X72Y103_SLICE_X108Y103_A5Q;
  assign CLBLL_R_X73Y102_SLICE_X111Y102_A3 = CLBLL_R_X73Y102_SLICE_X111Y102_AQ;
  assign CLBLL_R_X73Y102_SLICE_X111Y102_A4 = CLBLM_L_X74Y102_SLICE_X112Y102_AQ;
  assign CLBLL_R_X73Y102_SLICE_X111Y102_A5 = CLBLM_L_X72Y103_SLICE_X108Y103_CO6;
  assign CLBLL_R_X73Y102_SLICE_X111Y102_A6 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X76Y134_SLICE_X116Y134_C1 = CLBLM_L_X76Y133_SLICE_X116Y133_AQ;
  assign CLBLL_R_X73Y102_SLICE_X111Y102_AX = CLBLL_R_X73Y103_SLICE_X110Y103_B5Q;
  assign CLBLL_R_X73Y102_SLICE_X111Y102_B1 = CLBLM_L_X72Y104_SLICE_X109Y104_BQ;
  assign CLBLL_R_X73Y102_SLICE_X111Y102_B2 = CLBLL_R_X73Y103_SLICE_X111Y103_AQ;
  assign CLBLL_R_X73Y102_SLICE_X111Y102_B3 = CLBLL_R_X73Y102_SLICE_X111Y102_AQ;
  assign CLBLL_R_X73Y102_SLICE_X111Y102_B4 = CLBLM_L_X72Y104_SLICE_X109Y104_B5Q;
  assign CLBLL_R_X73Y102_SLICE_X111Y102_B5 = CLBLL_R_X73Y102_SLICE_X111Y102_A5Q;
  assign CLBLL_R_X73Y102_SLICE_X111Y102_B6 = CLBLM_L_X60Y101_SLICE_X90Y101_AQ;
  assign CLBLM_L_X76Y134_SLICE_X116Y134_C2 = CLBLM_L_X76Y134_SLICE_X117Y134_CO6;
  assign CLBLM_L_X76Y134_SLICE_X116Y134_C3 = CLBLM_L_X76Y134_SLICE_X116Y134_BQ;
  assign CLBLL_R_X73Y102_SLICE_X111Y102_C1 = CLBLM_L_X72Y103_SLICE_X109Y103_DO6;
  assign CLBLL_R_X73Y102_SLICE_X111Y102_C2 = CLBLM_L_X74Y103_SLICE_X112Y103_DO6;
  assign CLBLL_R_X73Y102_SLICE_X111Y102_C3 = CLBLL_R_X73Y102_SLICE_X110Y102_DO6;
  assign CLBLL_R_X73Y102_SLICE_X111Y102_C4 = CLBLM_L_X74Y103_SLICE_X112Y103_CO6;
  assign CLBLL_R_X73Y102_SLICE_X111Y102_C5 = CLBLL_R_X73Y102_SLICE_X111Y102_DO6;
  assign CLBLL_R_X73Y102_SLICE_X111Y102_C6 = CLBLL_R_X73Y102_SLICE_X111Y102_BO6;
  assign CLBLM_L_X76Y134_SLICE_X116Y134_C4 = CLBLL_R_X75Y134_SLICE_X115Y134_AQ;
  assign CLBLM_L_X76Y134_SLICE_X116Y134_C5 = CLBLM_L_X76Y134_SLICE_X116Y134_AQ;
  assign CLBLL_R_X73Y102_SLICE_X111Y102_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X76Y134_SLICE_X116Y134_C6 = CLBLL_R_X75Y133_SLICE_X115Y133_BQ;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_C2 = 1'b1;
  assign CLBLL_R_X73Y102_SLICE_X111Y102_D1 = CLBLL_R_X73Y103_SLICE_X110Y103_B5Q;
  assign CLBLL_R_X73Y102_SLICE_X111Y102_D2 = 1'b1;
  assign CLBLL_R_X73Y102_SLICE_X111Y102_D3 = CLBLL_R_X73Y104_SLICE_X110Y104_A5Q;
  assign CLBLL_R_X73Y102_SLICE_X111Y102_D4 = CLBLM_L_X74Y103_SLICE_X113Y103_BQ;
  assign CLBLL_R_X73Y102_SLICE_X111Y102_D5 = CLBLM_L_X72Y104_SLICE_X109Y104_BQ;
  assign CLBLL_R_X73Y102_SLICE_X111Y102_D6 = CLBLM_L_X72Y104_SLICE_X109Y104_B5Q;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_C3 = 1'b1;
  assign CLBLL_R_X73Y102_SLICE_X111Y102_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_C5 = 1'b1;
  assign CLBLM_L_X76Y134_SLICE_X116Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X76Y134_SLICE_X116Y134_D1 = CLBLM_L_X76Y134_SLICE_X117Y134_AQ;
  assign CLBLM_L_X76Y134_SLICE_X116Y134_D2 = CLBLL_R_X75Y134_SLICE_X114Y134_A5Q;
  assign CLBLM_L_X74Y133_SLICE_X112Y133_B4 = CLBLM_L_X74Y132_SLICE_X112Y132_BO6;
  assign CLBLM_L_X76Y134_SLICE_X116Y134_D3 = CLBLM_L_X76Y134_SLICE_X116Y134_AQ;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_A1 = CLBLM_L_X74Y129_SLICE_X113Y129_BO5;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_D1 = 1'b1;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_A3 = CLBLM_L_X72Y121_SLICE_X109Y121_AQ;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_A4 = CLBLL_R_X73Y132_SLICE_X111Y132_AO6;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_A5 = CLBLM_L_X74Y122_SLICE_X112Y122_BQ;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_D2 = 1'b1;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_A6 = 1'b1;
  assign CLBLM_L_X76Y134_SLICE_X116Y134_D4 = CLBLL_R_X75Y133_SLICE_X115Y133_AQ;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_B1 = 1'b1;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_B2 = 1'b1;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_B3 = 1'b1;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_B4 = 1'b1;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_B5 = 1'b1;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_B6 = 1'b1;
  assign CLBLM_L_X76Y134_SLICE_X116Y134_D6 = CLBLL_R_X75Y134_SLICE_X115Y134_AO6;
  assign CLBLM_R_X103Y75_SLICE_X163Y75_B2 = 1'b1;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_C1 = 1'b1;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_C2 = 1'b1;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_C3 = 1'b1;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_C4 = 1'b1;
  assign CLBLM_L_X68Y109_SLICE_X103Y109_A1 = CLBLM_R_X67Y110_SLICE_X101Y110_DQ;
  assign CLBLM_L_X68Y109_SLICE_X103Y109_A2 = CLBLM_L_X70Y106_SLICE_X105Y106_DO6;
  assign CLBLM_L_X68Y109_SLICE_X103Y109_A3 = CLBLM_L_X68Y109_SLICE_X102Y109_CO6;
  assign CLBLM_L_X68Y109_SLICE_X103Y109_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y109_SLICE_X103Y109_A5 = 1'b1;
  assign CLBLM_L_X68Y109_SLICE_X103Y109_A6 = CLBLM_L_X68Y109_SLICE_X103Y109_AQ;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_C5 = 1'b1;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_C6 = 1'b1;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X68Y109_SLICE_X103Y109_B1 = CLBLM_L_X68Y109_SLICE_X103Y109_B5Q;
  assign CLBLM_L_X68Y109_SLICE_X103Y109_B2 = CLBLM_L_X68Y109_SLICE_X103Y109_BQ;
  assign CLBLM_L_X68Y109_SLICE_X103Y109_B3 = CLBLM_L_X68Y106_SLICE_X103Y106_BQ;
  assign CLBLM_L_X68Y109_SLICE_X103Y109_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y109_SLICE_X103Y109_B5 = CLBLM_L_X68Y106_SLICE_X103Y106_AO5;
  assign CLBLM_L_X68Y109_SLICE_X103Y109_B6 = 1'b1;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_D1 = 1'b1;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_D2 = 1'b1;
  assign CLBLM_L_X68Y109_SLICE_X103Y109_C1 = 1'b1;
  assign CLBLM_L_X68Y109_SLICE_X103Y109_C2 = 1'b1;
  assign CLBLM_L_X68Y109_SLICE_X103Y109_C3 = 1'b1;
  assign CLBLM_L_X68Y109_SLICE_X103Y109_C4 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_A1 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_A2 = CLBLM_R_X63Y99_SLICE_X94Y99_CO6;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_A3 = CLBLM_L_X62Y97_SLICE_X93Y97_AQ;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_A5 = CLBLM_R_X63Y96_SLICE_X94Y96_BQ;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_A6 = CLBLM_L_X64Y97_SLICE_X97Y97_BO6;
  assign CLBLM_L_X68Y109_SLICE_X103Y109_C5 = 1'b1;
  assign CLBLM_L_X68Y109_SLICE_X103Y109_C6 = 1'b1;
  assign CLBLM_L_X68Y109_SLICE_X103Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_B1 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_B2 = CLBLM_L_X62Y97_SLICE_X93Y97_BQ;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_B3 = CLBLM_L_X62Y97_SLICE_X93Y97_AQ;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_B4 = CLBLM_R_X63Y99_SLICE_X94Y99_CO5;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_B6 = CLBLM_L_X64Y97_SLICE_X97Y97_BO6;
  assign CLBLM_L_X68Y109_SLICE_X103Y109_D1 = 1'b1;
  assign CLBLM_L_X68Y109_SLICE_X103Y109_D2 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_C1 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_C2 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_C3 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_C4 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_C5 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_C6 = 1'b1;
  assign CLBLM_L_X68Y109_SLICE_X103Y109_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X68Y109_SLICE_X102Y109_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y109_SLICE_X102Y109_A2 = CLBLM_R_X65Y109_SLICE_X99Y109_A5Q;
  assign CLBLM_L_X68Y109_SLICE_X102Y109_A3 = CLBLM_R_X67Y109_SLICE_X100Y109_DO5;
  assign CLBLM_L_X68Y109_SLICE_X102Y109_A4 = CLBLM_L_X70Y114_SLICE_X104Y114_AQ;
  assign CLBLM_L_X68Y109_SLICE_X102Y109_A5 = CLBLM_L_X68Y109_SLICE_X102Y109_A5Q;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_D1 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_D2 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_D3 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_D4 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_D5 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_D6 = 1'b1;
  assign CLBLM_L_X68Y109_SLICE_X102Y109_B1 = CLBLM_R_X67Y109_SLICE_X101Y109_AQ;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X68Y109_SLICE_X102Y109_B2 = CLBLM_L_X68Y108_SLICE_X102Y108_A5Q;
  assign CLBLM_L_X68Y109_SLICE_X102Y109_B3 = CLBLM_L_X68Y108_SLICE_X102Y108_AQ;
  assign CLBLM_L_X68Y109_SLICE_X102Y109_C2 = CLBLM_L_X68Y109_SLICE_X102Y109_BO5;
  assign CLBLM_L_X68Y109_SLICE_X102Y109_C3 = CLBLM_L_X70Y106_SLICE_X105Y106_DO6;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_A1 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_A2 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_A3 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_A4 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_A5 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_A6 = 1'b1;
  assign CLBLM_L_X68Y109_SLICE_X102Y109_C1 = CLBLM_R_X65Y108_SLICE_X99Y108_AO6;
  assign CLBLM_L_X68Y109_SLICE_X102Y109_C4 = CLBLM_R_X65Y110_SLICE_X99Y110_CO6;
  assign CLBLM_L_X68Y109_SLICE_X102Y109_C5 = CLBLM_L_X68Y109_SLICE_X102Y109_DO6;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_B1 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_B2 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_B3 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_B4 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_B5 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_B6 = 1'b1;
  assign CLBLM_L_X68Y109_SLICE_X102Y109_D4 = CLBLM_L_X68Y109_SLICE_X102Y109_A5Q;
  assign CLBLM_L_X68Y109_SLICE_X102Y109_D5 = CLBLM_R_X65Y111_SLICE_X98Y111_AQ;
  assign CLBLM_L_X68Y109_SLICE_X102Y109_D6 = CLBLM_R_X67Y108_SLICE_X101Y108_AO5;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_C1 = 1'b1;
  assign CLBLM_L_X68Y109_SLICE_X102Y109_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_C2 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_C3 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_C4 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_C5 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_C6 = 1'b1;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_B6 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_D1 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_D2 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_D3 = 1'b1;
  assign CLBLL_R_X73Y103_SLICE_X110Y103_A1 = CLBLM_L_X72Y103_SLICE_X108Y103_BO6;
  assign CLBLL_R_X73Y103_SLICE_X110Y103_A2 = CLBLM_L_X72Y103_SLICE_X108Y103_CO6;
  assign CLBLL_R_X73Y103_SLICE_X110Y103_A3 = CLBLL_R_X73Y103_SLICE_X110Y103_AQ;
  assign CLBLL_R_X73Y103_SLICE_X110Y103_A4 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLL_R_X73Y103_SLICE_X110Y103_A5 = CLBLL_R_X73Y102_SLICE_X110Y102_AQ;
  assign CLBLL_R_X73Y103_SLICE_X110Y103_A6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y102_SLICE_X103Y102_C3 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_D4 = 1'b1;
  assign CLBLL_R_X73Y103_SLICE_X110Y103_AX = CLBLM_L_X60Y101_SLICE_X90Y101_AQ;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_D5 = 1'b1;
  assign CLBLL_R_X73Y103_SLICE_X110Y103_B1 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLL_R_X73Y103_SLICE_X110Y103_B2 = CLBLL_R_X73Y103_SLICE_X110Y103_BQ;
  assign CLBLL_R_X73Y103_SLICE_X110Y103_B3 = CLBLL_R_X73Y103_SLICE_X110Y103_AQ;
  assign CLBLL_R_X73Y103_SLICE_X110Y103_B4 = CLBLM_L_X72Y103_SLICE_X108Y103_BO5;
  assign CLBLL_R_X73Y103_SLICE_X110Y103_B5 = CLBLM_L_X72Y103_SLICE_X108Y103_CO6;
  assign CLBLL_R_X73Y103_SLICE_X110Y103_B6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y102_SLICE_X103Y102_C4 = 1'b1;
  assign CLBLM_L_X68Y102_SLICE_X103Y102_C5 = 1'b1;
  assign CLBLL_R_X73Y103_SLICE_X110Y103_BX = CLBLM_L_X72Y103_SLICE_X109Y103_AQ;
  assign CLBLM_L_X72Y130_SLICE_X108Y130_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y103_SLICE_X110Y103_C1 = CLBLM_L_X72Y104_SLICE_X109Y104_BQ;
  assign CLBLL_R_X73Y103_SLICE_X110Y103_C2 = CLBLL_R_X73Y103_SLICE_X110Y103_AQ;
  assign CLBLL_R_X73Y103_SLICE_X110Y103_C3 = CLBLL_R_X75Y103_SLICE_X115Y103_AQ;
  assign CLBLL_R_X73Y103_SLICE_X110Y103_C4 = CLBLL_R_X73Y104_SLICE_X110Y104_A5Q;
  assign CLBLL_R_X73Y103_SLICE_X110Y103_C5 = CLBLM_L_X72Y104_SLICE_X109Y104_B5Q;
  assign CLBLL_R_X73Y103_SLICE_X110Y103_C6 = 1'b1;
  assign CLBLM_L_X68Y102_SLICE_X103Y102_C6 = 1'b1;
  assign CLBLM_R_X67Y115_SLICE_X101Y115_A6 = 1'b1;
  assign CLBLL_R_X73Y103_SLICE_X110Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X73Y103_SLICE_X110Y103_D1 = CLBLL_R_X73Y102_SLICE_X110Y102_AQ;
  assign CLBLL_R_X73Y103_SLICE_X110Y103_D2 = CLBLL_R_X73Y104_SLICE_X110Y104_A5Q;
  assign CLBLL_R_X73Y103_SLICE_X110Y103_D3 = CLBLL_R_X73Y103_SLICE_X111Y103_DO6;
  assign CLBLL_R_X73Y103_SLICE_X110Y103_D4 = CLBLL_R_X73Y103_SLICE_X110Y103_CO6;
  assign CLBLL_R_X73Y103_SLICE_X110Y103_D5 = CLBLM_L_X72Y103_SLICE_X109Y103_AO5;
  assign CLBLL_R_X73Y103_SLICE_X110Y103_D6 = CLBLL_R_X73Y102_SLICE_X110Y102_A5Q;
  assign CLBLL_R_X73Y103_SLICE_X110Y103_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y130_SLICE_X108Y130_C2 = CLBLM_L_X72Y130_SLICE_X108Y130_CQ;
  assign CLBLM_R_X103Y75_SLICE_X163Y75_BX = CLBLM_R_X103Y75_SLICE_X162Y75_CQ;
  assign CLBLM_L_X72Y130_SLICE_X108Y130_C3 = CLBLM_L_X72Y131_SLICE_X109Y131_DQ;
  assign CLBLL_R_X73Y103_SLICE_X111Y103_A1 = CLBLL_R_X73Y104_SLICE_X110Y104_DO6;
  assign CLBLL_R_X73Y103_SLICE_X111Y103_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y103_SLICE_X111Y103_A3 = CLBLL_R_X73Y103_SLICE_X111Y103_AQ;
  assign CLBLL_R_X73Y103_SLICE_X111Y103_A4 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLL_R_X73Y103_SLICE_X111Y103_A5 = CLBLM_L_X72Y103_SLICE_X108Y103_DO5;
  assign CLBLL_R_X73Y103_SLICE_X111Y103_A6 = CLBLM_L_X74Y103_SLICE_X113Y103_BQ;
  assign CLBLM_L_X68Y102_SLICE_X103Y102_D1 = 1'b1;
  assign CLBLM_L_X68Y102_SLICE_X103Y102_D2 = 1'b1;
  assign CLBLL_R_X73Y103_SLICE_X111Y103_AX = CLBLL_R_X79Y104_SLICE_X122Y104_A5Q;
  assign CLBLL_R_X73Y103_SLICE_X111Y103_B1 = CLBLM_L_X74Y103_SLICE_X113Y103_DO6;
  assign CLBLL_R_X73Y103_SLICE_X111Y103_B2 = CLBLL_R_X73Y103_SLICE_X110Y103_DO6;
  assign CLBLL_R_X73Y103_SLICE_X111Y103_B3 = CLBLM_L_X70Y105_SLICE_X104Y105_BO6;
  assign CLBLL_R_X73Y103_SLICE_X111Y103_B4 = CLBLL_R_X75Y103_SLICE_X114Y103_BO6;
  assign CLBLL_R_X73Y103_SLICE_X111Y103_B5 = CLBLL_R_X73Y102_SLICE_X111Y102_CO6;
  assign CLBLL_R_X73Y103_SLICE_X111Y103_B6 = CLBLL_R_X73Y103_SLICE_X111Y103_CO6;
  assign CLBLM_L_X68Y102_SLICE_X103Y102_D3 = 1'b1;
  assign CLBLM_L_X68Y102_SLICE_X103Y102_D4 = 1'b1;
  assign CLBLL_R_X73Y103_SLICE_X111Y103_C1 = CLBLM_L_X72Y104_SLICE_X109Y104_BQ;
  assign CLBLL_R_X73Y103_SLICE_X111Y103_C2 = CLBLM_L_X72Y104_SLICE_X109Y104_B5Q;
  assign CLBLL_R_X73Y103_SLICE_X111Y103_C3 = CLBLL_R_X73Y104_SLICE_X111Y104_CO6;
  assign CLBLL_R_X73Y103_SLICE_X111Y103_C4 = CLBLL_R_X79Y104_SLICE_X122Y104_A5Q;
  assign CLBLL_R_X73Y103_SLICE_X111Y103_C5 = CLBLL_R_X73Y103_SLICE_X110Y103_CO5;
  assign CLBLL_R_X73Y103_SLICE_X111Y103_C6 = CLBLL_R_X73Y103_SLICE_X110Y103_BQ;
  assign CLBLM_L_X68Y102_SLICE_X103Y102_D5 = 1'b1;
  assign CLBLM_L_X68Y102_SLICE_X103Y102_D6 = 1'b1;
  assign CLBLL_R_X73Y103_SLICE_X111Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X72Y130_SLICE_X108Y130_C4 = CLBLM_L_X72Y129_SLICE_X108Y129_AO5;
  assign CLBLL_R_X73Y103_SLICE_X111Y103_D1 = CLBLM_L_X60Y101_SLICE_X90Y101_AQ;
  assign CLBLL_R_X73Y103_SLICE_X111Y103_D2 = CLBLL_R_X73Y104_SLICE_X110Y104_A5Q;
  assign CLBLL_R_X73Y103_SLICE_X111Y103_D3 = CLBLM_L_X72Y104_SLICE_X109Y104_BQ;
  assign CLBLL_R_X73Y103_SLICE_X111Y103_D4 = 1'b1;
  assign CLBLL_R_X73Y103_SLICE_X111Y103_D5 = CLBLM_L_X72Y104_SLICE_X109Y104_B5Q;
  assign CLBLL_R_X73Y103_SLICE_X111Y103_D6 = CLBLL_R_X73Y104_SLICE_X111Y104_BQ;
  assign CLBLL_R_X73Y103_SLICE_X111Y103_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y130_SLICE_X108Y130_C5 = CLBLM_L_X72Y130_SLICE_X108Y130_BQ;
  assign CLBLM_L_X68Y102_SLICE_X102Y102_A1 = 1'b1;
  assign CLBLM_L_X68Y102_SLICE_X102Y102_A2 = CLBLM_L_X68Y97_SLICE_X102Y97_CO6;
  assign CLBLM_L_X72Y130_SLICE_X108Y130_C6 = 1'b1;
  assign CLBLM_L_X68Y102_SLICE_X102Y102_A3 = CLBLM_L_X68Y102_SLICE_X102Y102_AQ;
  assign CLBLM_L_X68Y102_SLICE_X102Y102_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X103Y75_SLICE_X163Y75_C3 = 1'b1;
  assign CLBLM_L_X68Y102_SLICE_X102Y102_A5 = CLBLM_L_X68Y102_SLICE_X102Y102_BQ;
  assign CLBLM_L_X68Y102_SLICE_X102Y102_A6 = CLBLM_L_X68Y99_SLICE_X102Y99_AO5;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_A1 = CLBLL_R_X71Y124_SLICE_X106Y124_CO6;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_A2 = CLBLM_L_X72Y122_SLICE_X109Y122_BQ;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_A3 = CLBLM_L_X72Y122_SLICE_X109Y122_AQ;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_A4 = CLBLL_R_X73Y123_SLICE_X111Y123_AQ;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_A6 = CLBLM_L_X72Y122_SLICE_X109Y122_A5Q;
  assign CLBLM_R_X103Y75_SLICE_X163Y75_C4 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_AX = CLBLM_L_X72Y122_SLICE_X109Y122_CO5;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_B1 = CLBLL_R_X71Y124_SLICE_X106Y124_CO6;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_B2 = CLBLM_L_X72Y122_SLICE_X109Y122_BQ;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_B3 = CLBLL_R_X73Y121_SLICE_X111Y121_AQ;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_B4 = CLBLL_R_X73Y122_SLICE_X111Y122_AO6;
  assign CLBLM_L_X68Y102_SLICE_X102Y102_B1 = CLBLM_R_X67Y98_SLICE_X100Y98_B5Q;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_B6 = CLBLM_L_X72Y122_SLICE_X109Y122_CO6;
  assign CLBLM_L_X68Y102_SLICE_X102Y102_B2 = CLBLM_L_X68Y102_SLICE_X102Y102_BQ;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_C2 = CLBLL_R_X71Y124_SLICE_X106Y124_CO6;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_C3 = CLBLL_R_X73Y123_SLICE_X111Y123_AQ;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_C4 = CLBLM_L_X72Y122_SLICE_X109Y122_A5Q;
  assign CLBLM_L_X68Y102_SLICE_X102Y102_B3 = CLBLM_L_X68Y102_SLICE_X102Y102_DQ;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_C5 = CLBLL_R_X73Y123_SLICE_X110Y123_CQ;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_C6 = 1'b1;
  assign CLBLM_R_X103Y75_SLICE_X163Y75_C5 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X68Y102_SLICE_X102Y102_B4 = CLBLM_R_X67Y98_SLICE_X100Y98_A5Q;
  assign LIOB33_X0Y61_IOB_X0Y61_O = CLBLM_R_X65Y109_SLICE_X98Y109_A5Q;
  assign LIOB33_X0Y61_IOB_X0Y62_O = CLBLM_R_X65Y110_SLICE_X99Y110_B5Q;
  assign CLBLM_L_X68Y102_SLICE_X102Y102_B5 = CLBLM_L_X68Y101_SLICE_X102Y101_BQ;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_D1 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_D2 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_D3 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_D4 = 1'b1;
  assign CLBLM_L_X68Y102_SLICE_X102Y102_B6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_D5 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_D6 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_A1 = CLBLM_L_X64Y98_SLICE_X96Y98_AO5;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_A2 = CLBLM_L_X64Y98_SLICE_X96Y98_BQ;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_A3 = CLBLM_L_X62Y98_SLICE_X93Y98_AQ;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_A4 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_A5 = CLBLM_R_X63Y99_SLICE_X94Y99_BO5;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_A6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_A1 = CLBLM_L_X72Y122_SLICE_X108Y122_BQ;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_A2 = CLBLM_L_X72Y123_SLICE_X108Y123_BQ;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_A3 = CLBLM_L_X72Y121_SLICE_X108Y121_AO6;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_B2 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_B3 = CLBLM_L_X62Y98_SLICE_X93Y98_AQ;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_B4 = CLBLM_R_X63Y99_SLICE_X94Y99_CO6;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_B5 = CLBLM_L_X62Y98_SLICE_X93Y98_BQ;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_B6 = CLBLM_L_X64Y98_SLICE_X96Y98_AO5;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_AX = CLBLM_L_X72Y121_SLICE_X108Y121_A5Q;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_B1 = 1'b1;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_C1 = CLBLM_L_X62Y98_SLICE_X93Y98_BQ;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_C2 = CLBLM_L_X62Y98_SLICE_X93Y98_CQ;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_C3 = CLBLM_R_X63Y99_SLICE_X94Y99_CO5;
  assign CLBLM_L_X68Y102_SLICE_X102Y102_C1 = CLBLM_L_X68Y102_SLICE_X102Y102_BQ;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_C4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_C5 = CLBLM_L_X64Y98_SLICE_X96Y98_AO5;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_C6 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X68Y102_SLICE_X102Y102_C2 = CLBLM_L_X68Y102_SLICE_X102Y102_CQ;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_BX = CLBLM_L_X72Y122_SLICE_X108Y122_AQ;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_C1 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_C2 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_C3 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_C4 = 1'b1;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_D1 = 1'b1;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_D2 = 1'b1;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_D3 = 1'b1;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_D4 = 1'b1;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_D5 = 1'b1;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_D6 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_CX = CLBLM_L_X72Y122_SLICE_X108Y122_BQ;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_D1 = 1'b1;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_D2 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_D3 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_D4 = 1'b1;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_A1 = 1'b1;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_A2 = 1'b1;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_A3 = 1'b1;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_A4 = 1'b1;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_A5 = 1'b1;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_A6 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X67Y115_SLICE_X101Y115_B6 = 1'b1;
  assign CLBLM_R_X67Y118_SLICE_X101Y118_D2 = 1'b1;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_B1 = 1'b1;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_B2 = 1'b1;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_B3 = 1'b1;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_B4 = 1'b1;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_B5 = 1'b1;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_B6 = 1'b1;
  assign CLBLM_R_X67Y118_SLICE_X101Y118_D3 = 1'b1;
  assign CLBLM_R_X67Y118_SLICE_X101Y118_D4 = 1'b1;
  assign CLBLM_L_X68Y102_SLICE_X102Y102_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X67Y118_SLICE_X101Y118_D5 = 1'b1;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_C1 = 1'b1;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_C2 = 1'b1;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_C3 = 1'b1;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_C4 = 1'b1;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_C5 = 1'b1;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_C6 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_D3 = 1'b1;
  assign CLBLM_R_X67Y118_SLICE_X101Y118_D6 = 1'b1;
  assign CLBLM_R_X103Y75_SLICE_X163Y75_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_D1 = CLBLM_L_X68Y107_SLICE_X102Y107_BO6;
  assign CLBLL_R_X73Y104_SLICE_X110Y104_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y104_SLICE_X110Y104_A2 = CLBLL_R_X73Y104_SLICE_X111Y104_DO6;
  assign CLBLL_R_X73Y104_SLICE_X110Y104_A3 = CLBLL_R_X73Y111_SLICE_X110Y111_AQ;
  assign CLBLL_R_X73Y104_SLICE_X110Y104_A4 = CLBLL_R_X73Y102_SLICE_X110Y102_A5Q;
  assign CLBLL_R_X73Y104_SLICE_X110Y104_A5 = CLBLL_R_X73Y104_SLICE_X110Y104_A5Q;
  assign CLBLL_R_X73Y104_SLICE_X110Y104_A6 = 1'b1;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_D1 = 1'b1;
  assign CLBLL_R_X73Y104_SLICE_X110Y104_B1 = CLBLM_L_X72Y104_SLICE_X109Y104_A5Q;
  assign CLBLL_R_X73Y104_SLICE_X110Y104_B2 = CLBLL_R_X73Y104_SLICE_X110Y104_BQ;
  assign CLBLL_R_X73Y104_SLICE_X110Y104_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y104_SLICE_X110Y104_B4 = CLBLM_L_X72Y103_SLICE_X108Y103_A5Q;
  assign CLBLL_R_X73Y104_SLICE_X110Y104_B5 = 1'b1;
  assign CLBLL_R_X73Y104_SLICE_X110Y104_B6 = 1'b1;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_D6 = 1'b1;
  assign CLBLM_L_X68Y102_SLICE_X102Y102_D1 = CLBLM_L_X68Y101_SLICE_X102Y101_BQ;
  assign CLBLL_R_X73Y104_SLICE_X110Y104_C1 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLL_R_X73Y104_SLICE_X110Y104_C2 = CLBLL_R_X73Y104_SLICE_X110Y104_CQ;
  assign CLBLL_R_X73Y104_SLICE_X110Y104_C3 = CLBLL_R_X73Y104_SLICE_X110Y104_BQ;
  assign CLBLL_R_X73Y104_SLICE_X110Y104_C4 = CLBLM_L_X72Y103_SLICE_X108Y103_BO6;
  assign CLBLL_R_X73Y104_SLICE_X110Y104_C5 = CLBLM_L_X72Y104_SLICE_X109Y104_A5Q;
  assign CLBLL_R_X73Y104_SLICE_X110Y104_C6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y133_SLICE_X109Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X73Y104_SLICE_X110Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_X0Y51_OLOGIC_X0Y51_D1 = CLBLM_L_X62Y101_SLICE_X92Y101_AQ;
  assign CLBLM_L_X76Y111_SLICE_X117Y111_C1 = 1'b1;
  assign CLBLL_R_X73Y104_SLICE_X110Y104_D1 = 1'b1;
  assign CLBLL_R_X73Y104_SLICE_X110Y104_D2 = 1'b1;
  assign CLBLL_R_X73Y104_SLICE_X110Y104_D3 = CLBLM_L_X72Y104_SLICE_X109Y104_A5Q;
  assign CLBLL_R_X73Y104_SLICE_X110Y104_D4 = CLBLL_R_X73Y104_SLICE_X110Y104_BQ;
  assign CLBLL_R_X73Y104_SLICE_X110Y104_D5 = 1'b1;
  assign CLBLL_R_X73Y104_SLICE_X110Y104_D6 = 1'b1;
  assign CLBLM_L_X68Y102_SLICE_X102Y102_D5 = CLBLM_R_X67Y98_SLICE_X100Y98_B5Q;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_D5 = 1'b1;
  assign CLBLL_R_X73Y104_SLICE_X110Y104_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X68Y102_SLICE_X102Y102_D6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign LIOI3_X0Y51_OLOGIC_X0Y51_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y58_T1 = 1'b1;
  assign CLBLM_R_X67Y118_SLICE_X100Y118_A6 = 1'b1;
  assign CLBLM_L_X76Y111_SLICE_X117Y111_C2 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y57_D1 = CLBLM_L_X62Y95_SLICE_X92Y95_AQ;
  assign CLBLM_L_X68Y102_SLICE_X102Y102_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X73Y104_SLICE_X111Y104_A1 = CLBLM_L_X74Y104_SLICE_X112Y104_CQ;
  assign CLBLL_R_X73Y104_SLICE_X111Y104_A2 = CLBLL_R_X73Y104_SLICE_X110Y104_DO5;
  assign CLBLL_R_X73Y104_SLICE_X111Y104_A3 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLL_R_X73Y104_SLICE_X111Y104_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y104_SLICE_X111Y104_A5 = CLBLM_L_X72Y103_SLICE_X108Y103_DO5;
  assign CLBLL_R_X73Y104_SLICE_X111Y104_A6 = CLBLL_R_X73Y104_SLICE_X111Y104_AQ;
  assign CLBLM_L_X72Y133_SLICE_X109Y133_D4 = CLBLL_R_X73Y133_SLICE_X111Y133_CO6;
  assign CLBLM_L_X72Y133_SLICE_X109Y133_D5 = CLBLL_R_X73Y133_SLICE_X110Y133_A5Q;
  assign LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y57_T1 = 1'b1;
  assign CLBLL_R_X73Y104_SLICE_X111Y104_B1 = CLBLL_R_X73Y104_SLICE_X111Y104_AQ;
  assign CLBLL_R_X73Y104_SLICE_X111Y104_B2 = CLBLL_R_X73Y104_SLICE_X111Y104_BQ;
  assign CLBLL_R_X73Y104_SLICE_X111Y104_B3 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLL_R_X73Y104_SLICE_X111Y104_B4 = CLBLL_R_X73Y104_SLICE_X110Y104_BO5;
  assign CLBLL_R_X73Y104_SLICE_X111Y104_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y104_SLICE_X111Y104_B6 = 1'b1;
  assign CLBLM_L_X72Y133_SLICE_X109Y133_D6 = CLBLM_L_X74Y134_SLICE_X113Y134_A5Q;
  assign CLBLM_L_X76Y111_SLICE_X117Y111_C3 = 1'b1;
  assign CLBLL_R_X73Y104_SLICE_X111Y104_C1 = CLBLL_R_X73Y102_SLICE_X110Y102_BQ;
  assign CLBLL_R_X73Y104_SLICE_X111Y104_C2 = CLBLL_R_X73Y104_SLICE_X110Y104_A5Q;
  assign CLBLL_R_X73Y104_SLICE_X111Y104_C3 = CLBLM_L_X62Y95_SLICE_X92Y95_AQ;
  assign CLBLL_R_X73Y104_SLICE_X111Y104_C4 = CLBLL_R_X73Y104_SLICE_X111Y104_AQ;
  assign CLBLL_R_X73Y104_SLICE_X111Y104_C5 = CLBLL_R_X73Y103_SLICE_X110Y103_B5Q;
  assign CLBLL_R_X73Y104_SLICE_X111Y104_C6 = CLBLL_R_X75Y103_SLICE_X115Y103_AQ;
  assign CLBLM_L_X74Y107_SLICE_X112Y107_B1 = CLBLM_L_X72Y108_SLICE_X108Y108_BO6;
  assign CLBLL_R_X73Y104_SLICE_X111Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X67Y115_SLICE_X101Y115_C1 = 1'b1;
  assign CLBLM_L_X72Y133_SLICE_X109Y133_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X67Y118_SLICE_X100Y118_B5 = 1'b1;
  assign CLBLL_R_X73Y104_SLICE_X111Y104_D1 = 1'b1;
  assign CLBLL_R_X73Y104_SLICE_X111Y104_D2 = CLBLL_R_X79Y104_SLICE_X122Y104_A5Q;
  assign CLBLL_R_X73Y104_SLICE_X111Y104_D3 = CLBLM_L_X62Y95_SLICE_X92Y95_AQ;
  assign CLBLL_R_X73Y104_SLICE_X111Y104_D4 = CLBLL_R_X73Y103_SLICE_X111Y103_A5Q;
  assign CLBLL_R_X73Y104_SLICE_X111Y104_D5 = 1'b1;
  assign CLBLL_R_X73Y104_SLICE_X111Y104_D6 = CLBLL_R_X75Y103_SLICE_X115Y103_AQ;
  assign CLBLM_L_X74Y107_SLICE_X112Y107_B4 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X76Y111_SLICE_X117Y111_C4 = 1'b1;
  assign CLBLL_R_X73Y104_SLICE_X111Y104_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X67Y118_SLICE_X100Y118_B6 = 1'b1;
  assign CLBLM_R_X67Y115_SLICE_X101Y115_C2 = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_D1 = 1'b1;
  assign CLBLM_L_X76Y111_SLICE_X117Y111_C5 = 1'b1;
  assign CLBLM_R_X67Y115_SLICE_X101Y115_C3 = 1'b1;
  assign CLBLM_L_X74Y107_SLICE_X112Y107_C3 = CLBLL_R_X73Y107_SLICE_X111Y107_DQ;
  assign CLBLM_L_X76Y111_SLICE_X117Y111_C6 = 1'b1;
  assign CLBLM_R_X67Y118_SLICE_X100Y118_C5 = 1'b1;
  assign CLBLM_L_X74Y107_SLICE_X112Y107_C4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X67Y118_SLICE_X100Y118_C6 = 1'b1;
  assign CLBLM_L_X74Y107_SLICE_X112Y107_C5 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X67Y115_SLICE_X101Y115_C4 = 1'b1;
  assign LIOB33_X0Y63_IOB_X0Y64_O = CLBLL_R_X73Y103_SLICE_X111Y103_A5Q;
  assign LIOB33_X0Y63_IOB_X0Y63_O = CLBLL_R_X73Y102_SLICE_X111Y102_A5Q;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_A1 = CLBLL_R_X73Y123_SLICE_X111Y123_DQ;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_A2 = CLBLL_R_X71Y124_SLICE_X106Y124_CO6;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_A3 = CLBLM_L_X72Y123_SLICE_X109Y123_AQ;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_A4 = CLBLM_L_X72Y122_SLICE_X109Y122_A5Q;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_A6 = CLBLM_L_X72Y122_SLICE_X109Y122_AQ;
  assign CLBLM_R_X67Y118_SLICE_X100Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_B1 = CLBLL_R_X73Y123_SLICE_X111Y123_DQ;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_B2 = CLBLM_L_X72Y123_SLICE_X109Y123_BQ;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_B3 = CLBLM_L_X72Y123_SLICE_X109Y123_AQ;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_B4 = 1'b1;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_B6 = CLBLM_L_X72Y123_SLICE_X109Y123_CO6;
  assign CLBLM_R_X67Y115_SLICE_X101Y115_C5 = 1'b1;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_C1 = 1'b1;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_C2 = CLBLL_R_X71Y124_SLICE_X106Y124_CO6;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_C3 = 1'b1;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_C4 = CLBLM_L_X72Y122_SLICE_X109Y122_AQ;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_C5 = 1'b1;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_C6 = CLBLM_L_X72Y122_SLICE_X109Y122_A5Q;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X72Y130_SLICE_X108Y130_D5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign RIOB33_X105Y151_IOB_X1Y152_O = 1'b1;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_D1 = 1'b1;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_D2 = 1'b1;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_D3 = 1'b1;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_D4 = 1'b1;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_D5 = 1'b1;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_D6 = 1'b1;
  assign CLBLM_R_X67Y115_SLICE_X101Y115_C6 = 1'b1;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_A1 = CLBLM_L_X60Y92_SLICE_X90Y92_BQ;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_A2 = CLBLM_L_X76Y111_SLICE_X116Y111_BQ;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_A3 = CLBLM_L_X62Y99_SLICE_X93Y99_AQ;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_A4 = CLBLM_L_X62Y99_SLICE_X93Y99_BO6;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_A5 = CLBLM_R_X63Y98_SLICE_X94Y98_BQ;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_A6 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_A1 = CLBLL_R_X73Y121_SLICE_X110Y121_CO6;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_A2 = CLBLM_L_X72Y122_SLICE_X109Y122_A5Q;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_A3 = CLBLM_L_X72Y123_SLICE_X108Y123_AQ;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_B1 = CLBLM_L_X60Y92_SLICE_X90Y92_BQ;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_B2 = CLBLM_L_X76Y111_SLICE_X116Y111_BQ;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_B3 = CLBLM_L_X62Y99_SLICE_X93Y99_AQ;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_B4 = CLBLM_R_X63Y98_SLICE_X94Y98_AQ;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_B5 = CLBLM_R_X63Y98_SLICE_X94Y98_BQ;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_B6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_AX = CLBLM_L_X72Y123_SLICE_X108Y123_BO5;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_B1 = CLBLL_R_X71Y129_SLICE_X107Y129_AO6;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_B2 = CLBLL_R_X71Y121_SLICE_X106Y121_A5Q;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_C1 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_C2 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_C3 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_C4 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_C5 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_C6 = 1'b1;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_BX = CLBLM_L_X72Y123_SLICE_X108Y123_CO5;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_C2 = CLBLL_R_X71Y129_SLICE_X107Y129_AO6;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_C3 = 1'b1;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_C4 = CLBLM_L_X72Y125_SLICE_X109Y125_CO6;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_C5 = CLBLL_R_X71Y121_SLICE_X106Y121_AQ;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_C6 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_D1 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_D2 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_D3 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_D4 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_D5 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_D6 = 1'b1;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_D1 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_D2 = 1'b1;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_D3 = 1'b1;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_D4 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_A1 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_A2 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_A3 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_A4 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_A5 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_A6 = 1'b1;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y133_SLICE_X108Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_B1 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_B2 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_B3 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_B4 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_B5 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_B6 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_C1 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_C2 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_C3 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_C4 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_C5 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_C6 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_D1 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_D2 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_D3 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_D4 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_D5 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_D6 = 1'b1;
  assign CLBLM_L_X72Y133_SLICE_X108Y133_D4 = CLBLM_L_X72Y133_SLICE_X108Y133_A5Q;
  assign CLBLM_L_X72Y133_SLICE_X108Y133_D5 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_A4 = CLBLL_R_X75Y128_SLICE_X115Y128_DO6;
  assign CLBLM_L_X72Y133_SLICE_X108Y133_D6 = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_D1 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_A5 = CLBLM_L_X74Y129_SLICE_X112Y129_A5Q;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_B3 = CLBLM_L_X74Y129_SLICE_X112Y129_A5Q;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_B4 = 1'b1;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_B5 = CLBLM_L_X74Y129_SLICE_X112Y129_AQ;
  assign RIOI3_X105Y145_OLOGIC_X1Y146_D1 = CLBLM_R_X63Y97_SLICE_X94Y97_AQ;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_A6 = 1'b1;
  assign CLBLM_L_X74Y133_SLICE_X112Y133_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_T1 = 1'b1;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_C2 = CLBLM_L_X74Y128_SLICE_X113Y128_CQ;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_C3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_C4 = CLBLL_R_X75Y128_SLICE_X115Y128_DO6;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_C5 = CLBLM_L_X74Y129_SLICE_X113Y129_AQ;
  assign CLBLM_L_X82Y130_SLICE_X128Y130_C3 = 1'b1;
  assign LIOB33_X0Y65_IOB_X0Y66_O = CLBLM_R_X65Y110_SLICE_X98Y110_A5Q;
  assign LIOB33_X0Y65_IOB_X0Y65_O = CLBLM_L_X72Y107_SLICE_X109Y107_BQ;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_D1 = 1'b1;
  assign CLBLM_R_X67Y115_SLICE_X101Y115_D1 = 1'b1;
  assign CLBLM_L_X82Y130_SLICE_X128Y130_C4 = 1'b1;
  assign CLBLM_R_X67Y115_SLICE_X101Y115_D2 = 1'b1;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_A1 = CLBLL_R_X73Y124_SLICE_X110Y124_A5Q;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_A2 = CLBLM_L_X72Y124_SLICE_X108Y124_BO6;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_A3 = CLBLM_L_X72Y124_SLICE_X109Y124_AQ;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_A4 = CLBLL_R_X73Y124_SLICE_X110Y124_AQ;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_A6 = CLBLL_R_X73Y124_SLICE_X110Y124_BQ;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_D5 = 1'b1;
  assign RIOB33_X105Y153_IOB_X1Y153_O = 1'b1;
  assign RIOB33_X105Y153_IOB_X1Y154_O = 1'b1;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_B1 = 1'b1;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_B2 = 1'b1;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_B3 = 1'b1;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_B4 = 1'b1;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_B5 = 1'b1;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_B6 = 1'b1;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_D6 = 1'b1;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_C1 = 1'b1;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_C2 = 1'b1;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_C3 = 1'b1;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_C4 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X103Y112_A1 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X103Y112_A2 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X103Y112_A3 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X103Y112_A4 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X103Y112_A5 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X103Y112_A6 = 1'b1;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_C5 = 1'b1;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_C6 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X103Y112_AX = CLBLL_R_X71Y112_SLICE_X106Y112_B5Q;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X68Y112_SLICE_X103Y112_B1 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X103Y112_B2 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X103Y112_B3 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X103Y112_B4 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X103Y112_B5 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X103Y112_B6 = 1'b1;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_D1 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X103Y112_BX = CLBLM_L_X68Y112_SLICE_X103Y112_AQ;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_D2 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X103Y112_C1 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X103Y112_C2 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X103Y112_C3 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X103Y112_C4 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X103Y112_C5 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_A1 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_A2 = CLBLM_L_X60Y99_SLICE_X90Y99_DQ;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_A3 = CLBLM_L_X60Y99_SLICE_X90Y99_BQ;
  assign CLBLM_L_X68Y112_SLICE_X103Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_A4 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_A5 = CLBLM_L_X62Y100_SLICE_X92Y100_AQ;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_A6 = CLBLM_L_X62Y101_SLICE_X92Y101_AQ;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_B1 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X103Y112_D1 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X103Y112_D2 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X103Y112_D3 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X103Y112_D4 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_B6 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X103Y112_D5 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_B2 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X103Y112_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_B3 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_B4 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_C4 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_C5 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_C6 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_C1 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X102Y112_A4 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_C2 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_C3 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X102Y112_A1 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X102Y112_A2 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X102Y112_A3 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_D1 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_D2 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_D3 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_D4 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X102Y112_B5 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X102Y112_B6 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_D5 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_D6 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X102Y112_B2 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X102Y112_C1 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X102Y112_C2 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X102Y112_C3 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X102Y112_C4 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X102Y112_C5 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X102Y112_C6 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_A1 = CLBLM_L_X62Y101_SLICE_X92Y101_AQ;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_A2 = CLBLM_L_X62Y101_SLICE_X92Y101_BO6;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_A3 = CLBLM_L_X62Y100_SLICE_X92Y100_AQ;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_A4 = CLBLM_L_X60Y99_SLICE_X90Y99_CQ;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_A5 = CLBLM_L_X60Y99_SLICE_X90Y99_BQ;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_A6 = CLBLM_L_X60Y99_SLICE_X90Y99_DQ;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_B1 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_B2 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_B4 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_B5 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_B6 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X102Y112_D1 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_B3 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X102Y112_D6 = 1'b1;
  assign CLBLM_L_X68Y112_SLICE_X102Y112_D2 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_C1 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_C2 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_C3 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_C4 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_C5 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_C6 = 1'b1;
  assign CLBLL_R_X73Y106_SLICE_X110Y106_A1 = CLBLM_L_X74Y107_SLICE_X113Y107_AQ;
  assign CLBLL_R_X73Y106_SLICE_X110Y106_A2 = CLBLL_R_X73Y107_SLICE_X111Y107_BQ;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X73Y106_SLICE_X110Y106_A3 = CLBLM_L_X62Y92_SLICE_X92Y92_AQ;
  assign CLBLL_R_X73Y106_SLICE_X110Y106_A4 = CLBLM_L_X72Y107_SLICE_X108Y107_BQ;
  assign CLBLL_R_X73Y106_SLICE_X110Y106_A5 = CLBLL_R_X71Y107_SLICE_X106Y107_C5Q;
  assign CLBLL_R_X73Y106_SLICE_X110Y106_A6 = CLBLL_R_X71Y107_SLICE_X106Y107_CQ;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_D1 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_D2 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_D3 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_D4 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_D5 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_D6 = 1'b1;
  assign CLBLL_R_X73Y106_SLICE_X110Y106_B1 = CLBLL_R_X73Y108_SLICE_X110Y108_A5Q;
  assign CLBLL_R_X73Y106_SLICE_X110Y106_B2 = CLBLM_L_X72Y107_SLICE_X108Y107_A5Q;
  assign CLBLL_R_X73Y106_SLICE_X110Y106_B3 = CLBLL_R_X71Y107_SLICE_X106Y107_C5Q;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X73Y106_SLICE_X110Y106_B5 = CLBLL_R_X73Y106_SLICE_X110Y106_AO6;
  assign CLBLL_R_X73Y106_SLICE_X110Y106_B6 = CLBLL_R_X71Y107_SLICE_X106Y107_CQ;
  assign CLBLL_R_X73Y106_SLICE_X110Y106_C1 = 1'b1;
  assign CLBLL_R_X73Y106_SLICE_X110Y106_C2 = 1'b1;
  assign CLBLL_R_X73Y106_SLICE_X110Y106_C3 = 1'b1;
  assign CLBLL_R_X73Y106_SLICE_X110Y106_C4 = 1'b1;
  assign CLBLL_R_X73Y106_SLICE_X110Y106_C5 = 1'b1;
  assign CLBLL_R_X73Y106_SLICE_X110Y106_C6 = 1'b1;
  assign RIOB33_X105Y127_IOB_X1Y128_O = CLBLM_R_X65Y110_SLICE_X99Y110_CQ;
  assign CLBLL_R_X73Y106_SLICE_X110Y106_D1 = 1'b1;
  assign CLBLL_R_X73Y106_SLICE_X110Y106_D2 = 1'b1;
  assign CLBLL_R_X73Y106_SLICE_X110Y106_D3 = 1'b1;
  assign CLBLL_R_X73Y106_SLICE_X110Y106_D4 = 1'b1;
  assign CLBLL_R_X73Y106_SLICE_X110Y106_D5 = 1'b1;
  assign CLBLL_R_X73Y106_SLICE_X110Y106_D6 = 1'b1;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_C1 = CLBLM_L_X74Y128_SLICE_X112Y128_CQ;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_C2 = CLBLM_L_X74Y129_SLICE_X112Y129_A5Q;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_C3 = CLBLM_L_X74Y128_SLICE_X112Y128_DQ;
  assign RIOB33_X105Y127_IOB_X1Y127_O = CLBLM_L_X72Y107_SLICE_X108Y107_A5Q;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_C4 = CLBLM_L_X74Y128_SLICE_X113Y128_BO6;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_C5 = CLBLL_R_X75Y128_SLICE_X114Y128_DO6;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_C6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y106_SLICE_X111Y106_A1 = 1'b1;
  assign CLBLL_R_X73Y106_SLICE_X111Y106_A2 = 1'b1;
  assign CLBLL_R_X73Y106_SLICE_X111Y106_A3 = 1'b1;
  assign CLBLL_R_X73Y106_SLICE_X111Y106_A4 = 1'b1;
  assign CLBLL_R_X73Y106_SLICE_X111Y106_A5 = 1'b1;
  assign CLBLL_R_X73Y106_SLICE_X111Y106_A6 = 1'b1;
  assign CLBLL_R_X73Y106_SLICE_X111Y106_B1 = 1'b1;
  assign CLBLL_R_X73Y106_SLICE_X111Y106_B2 = 1'b1;
  assign CLBLL_R_X73Y106_SLICE_X111Y106_B3 = 1'b1;
  assign CLBLL_R_X73Y106_SLICE_X111Y106_B4 = 1'b1;
  assign CLBLL_R_X73Y106_SLICE_X111Y106_B5 = 1'b1;
  assign CLBLL_R_X73Y106_SLICE_X111Y106_B6 = 1'b1;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_D1 = CLBLM_R_X67Y108_SLICE_X100Y108_AO6;
  assign LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y58_D1 = CLBLM_L_X72Y107_SLICE_X108Y107_BQ;
  assign CLBLL_R_X73Y106_SLICE_X111Y106_C1 = 1'b1;
  assign CLBLL_R_X73Y106_SLICE_X111Y106_C2 = 1'b1;
  assign CLBLL_R_X73Y106_SLICE_X111Y106_C3 = 1'b1;
  assign CLBLL_R_X73Y106_SLICE_X111Y106_C4 = 1'b1;
  assign CLBLL_R_X73Y106_SLICE_X111Y106_C5 = 1'b1;
  assign CLBLL_R_X73Y106_SLICE_X111Y106_C6 = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_D1 = CLBLM_L_X70Y135_SLICE_X104Y135_CO6;
  assign CLBLL_R_X73Y106_SLICE_X111Y106_D1 = 1'b1;
  assign CLBLL_R_X73Y106_SLICE_X111Y106_D2 = 1'b1;
  assign CLBLL_R_X73Y106_SLICE_X111Y106_D3 = 1'b1;
  assign CLBLL_R_X73Y106_SLICE_X111Y106_D4 = 1'b1;
  assign CLBLL_R_X73Y106_SLICE_X111Y106_D5 = 1'b1;
  assign CLBLL_R_X73Y106_SLICE_X111Y106_D6 = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_T1 = 1'b1;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_D1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_D1 = CLBLM_R_X63Y105_SLICE_X95Y105_A5Q;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_D2 = CLBLM_L_X74Y127_SLICE_X113Y127_CQ;
  assign LIOB33_X0Y67_IOB_X0Y68_O = CLBLL_R_X71Y134_SLICE_X106Y134_AQ;
  assign LIOB33_X0Y67_IOB_X0Y67_O = CLBLM_L_X72Y103_SLICE_X109Y103_AQ;
  assign LIOI3_X0Y53_OLOGIC_X0Y54_D1 = CLBLM_L_X62Y92_SLICE_X92Y92_AQ;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_D3 = CLBLM_L_X74Y128_SLICE_X112Y128_DQ;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_T1 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_C6 = 1'b1;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_D4 = CLBLL_R_X75Y128_SLICE_X115Y128_DO6;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_D5 = CLBLM_L_X74Y127_SLICE_X112Y127_AO6;
  assign LIOI3_X0Y53_OLOGIC_X0Y54_T1 = 1'b1;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_D6 = CLBLL_R_X75Y128_SLICE_X114Y128_DO6;
  assign LIOI3_X0Y53_OLOGIC_X0Y53_D1 = CLBLM_L_X62Y90_SLICE_X92Y90_AQ;
  assign LIOI3_TBYTESRC_X0Y69_OLOGIC_X0Y70_D1 = CLBLL_R_X75Y127_SLICE_X115Y127_AQ;
  assign LIOI3_X0Y53_OLOGIC_X0Y53_T1 = 1'b1;
  assign CLBLM_L_X76Y111_SLICE_X116Y111_A3 = 1'b1;
  assign RIOB33_X105Y155_IOB_X1Y155_O = 1'b1;
  assign RIOB33_X105Y155_IOB_X1Y156_O = 1'b1;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign LIOI3_TBYTESRC_X0Y69_OLOGIC_X0Y70_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y69_OLOGIC_X0Y69_D1 = CLBLM_L_X60Y92_SLICE_X90Y92_AQ;
  assign CLBLM_L_X76Y111_SLICE_X116Y111_A4 = 1'b1;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_A1 = CLBLM_L_X72Y125_SLICE_X109Y125_AQ;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_A2 = CLBLM_L_X72Y124_SLICE_X108Y124_AQ;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_A3 = CLBLL_R_X73Y124_SLICE_X110Y124_CO5;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_A4 = CLBLM_L_X74Y126_SLICE_X113Y126_CQ;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_A6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y69_OLOGIC_X0Y69_T1 = 1'b1;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_B1 = CLBLM_L_X72Y125_SLICE_X109Y125_AQ;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_B2 = CLBLM_L_X72Y125_SLICE_X109Y125_BQ;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_B3 = CLBLM_L_X72Y124_SLICE_X109Y124_AQ;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_B4 = CLBLM_L_X72Y124_SLICE_X108Y124_BO6;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_B6 = CLBLL_R_X73Y124_SLICE_X110Y124_BQ;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_C1 = 1'b1;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_C2 = CLBLL_R_X73Y128_SLICE_X111Y128_BQ;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_C3 = CLBLL_R_X75Y127_SLICE_X115Y127_CQ;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_C4 = CLBLL_R_X73Y122_SLICE_X111Y122_DQ;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_C5 = CLBLM_L_X72Y125_SLICE_X109Y125_DO6;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_C6 = CLBLM_L_X72Y126_SLICE_X108Y126_BQ;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_D1 = CLBLM_L_X72Y123_SLICE_X109Y123_BQ;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_D2 = CLBLM_L_X72Y126_SLICE_X109Y126_CQ;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_D3 = 1'b1;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_D4 = CLBLM_L_X72Y125_SLICE_X108Y125_CQ;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_D5 = 1'b1;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_D6 = CLBLL_R_X73Y125_SLICE_X111Y125_CQ;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_A1 = CLBLM_L_X64Y101_SLICE_X96Y101_A5Q;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_A2 = CLBLM_L_X64Y101_SLICE_X96Y101_BQ;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_A3 = CLBLM_L_X62Y100_SLICE_X92Y100_AQ;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_A4 = CLBLM_L_X62Y103_SLICE_X93Y103_AQ;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_A5 = CLBLM_L_X64Y101_SLICE_X96Y101_B5Q;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_A6 = 1'b1;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_A1 = 1'b1;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_A2 = CLBLL_R_X73Y125_SLICE_X110Y125_AO6;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_A3 = CLBLM_L_X72Y125_SLICE_X108Y125_AQ;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_B1 = CLBLM_L_X60Y99_SLICE_X90Y99_BQ;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_B2 = CLBLM_L_X64Y101_SLICE_X96Y101_BQ;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_B3 = CLBLM_L_X60Y99_SLICE_X90Y99_DQ;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_B4 = CLBLM_L_X64Y101_SLICE_X96Y101_B5Q;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_B5 = CLBLM_L_X62Y102_SLICE_X93Y102_DQ;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_B6 = CLBLM_L_X62Y102_SLICE_X93Y102_CQ;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_B1 = CLBLL_R_X73Y125_SLICE_X111Y125_DQ;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_B2 = CLBLM_L_X72Y125_SLICE_X108Y125_BQ;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_C1 = CLBLM_L_X62Y101_SLICE_X93Y101_AO6;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_C2 = CLBLM_L_X62Y102_SLICE_X92Y102_AQ;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_C3 = CLBLM_L_X62Y101_SLICE_X92Y101_AQ;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_C4 = CLBLM_R_X63Y101_SLICE_X94Y101_BO6;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_C5 = CLBLM_L_X62Y101_SLICE_X92Y101_AO6;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_C6 = CLBLM_L_X62Y101_SLICE_X93Y101_BO6;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_C2 = CLBLM_L_X72Y125_SLICE_X108Y125_CQ;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_C3 = CLBLM_L_X72Y125_SLICE_X108Y125_BQ;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_C4 = CLBLL_R_X73Y125_SLICE_X111Y125_DQ;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_C5 = CLBLM_L_X72Y125_SLICE_X108Y125_DO6;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_C6 = 1'b1;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_D1 = CLBLM_R_X63Y101_SLICE_X94Y101_AO6;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_D2 = CLBLM_R_X63Y101_SLICE_X94Y101_BQ;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_D3 = CLBLM_R_X63Y101_SLICE_X94Y101_BO6;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_D4 = CLBLM_L_X62Y101_SLICE_X93Y101_AO5;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_D5 = CLBLM_L_X64Y101_SLICE_X96Y101_A5Q;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_D6 = CLBLM_L_X62Y103_SLICE_X93Y103_BQ;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_D1 = CLBLM_L_X72Y124_SLICE_X109Y124_AQ;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_D2 = 1'b1;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_D3 = 1'b1;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_D4 = CLBLL_R_X73Y124_SLICE_X110Y124_BQ;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_D5 = 1'b1;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_A1 = CLBLM_L_X60Y99_SLICE_X90Y99_BQ;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_A2 = CLBLM_L_X62Y102_SLICE_X92Y102_BQ;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_A3 = CLBLM_L_X62Y102_SLICE_X92Y102_CQ;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_A4 = CLBLM_L_X64Y101_SLICE_X96Y101_B5Q;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_A5 = CLBLM_L_X60Y99_SLICE_X90Y99_DQ;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_A6 = CLBLM_L_X64Y101_SLICE_X96Y101_BQ;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_AX = CLBLM_L_X62Y100_SLICE_X92Y100_AQ;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_B1 = CLBLM_R_X63Y101_SLICE_X94Y101_AQ;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_B2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_B3 = CLBLM_L_X62Y101_SLICE_X92Y101_AQ;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_B4 = CLBLM_L_X60Y99_SLICE_X90Y99_CQ;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_B5 = CLBLM_L_X62Y100_SLICE_X92Y100_AQ;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_B6 = CLBLM_L_X60Y99_SLICE_X90Y99_DQ;
  assign CLBLL_R_X73Y107_SLICE_X110Y107_A1 = CLBLM_L_X72Y107_SLICE_X109Y107_AQ;
  assign CLBLL_R_X73Y107_SLICE_X110Y107_A2 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLL_R_X73Y107_SLICE_X110Y107_A3 = CLBLL_R_X73Y107_SLICE_X110Y107_AQ;
  assign CLBLL_R_X73Y107_SLICE_X110Y107_A4 = CLBLM_L_X72Y108_SLICE_X108Y108_BO6;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_C4 = 1'b1;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_C5 = 1'b1;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_C6 = 1'b1;
  assign CLBLL_R_X73Y107_SLICE_X110Y107_A5 = CLBLM_L_X72Y108_SLICE_X109Y108_BO6;
  assign CLBLL_R_X73Y107_SLICE_X110Y107_A6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_C1 = 1'b1;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_C2 = 1'b1;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_C3 = 1'b1;
  assign CLBLL_R_X73Y107_SLICE_X110Y107_B1 = CLBLM_L_X72Y109_SLICE_X108Y109_BO6;
  assign CLBLL_R_X73Y107_SLICE_X110Y107_B2 = CLBLL_R_X73Y107_SLICE_X110Y107_BQ;
  assign CLBLL_R_X73Y107_SLICE_X110Y107_B3 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLL_R_X73Y107_SLICE_X110Y107_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y107_SLICE_X110Y107_B5 = CLBLM_L_X72Y108_SLICE_X109Y108_BO6;
  assign CLBLL_R_X73Y107_SLICE_X110Y107_B6 = CLBLM_L_X74Y107_SLICE_X112Y107_AQ;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_D1 = 1'b1;
  assign CLBLL_R_X73Y107_SLICE_X110Y107_C1 = CLBLL_R_X73Y107_SLICE_X111Y107_AQ;
  assign CLBLL_R_X73Y107_SLICE_X110Y107_C2 = CLBLL_R_X71Y107_SLICE_X106Y107_CQ;
  assign CLBLL_R_X73Y107_SLICE_X110Y107_C3 = CLBLM_L_X72Y107_SLICE_X109Y107_A5Q;
  assign CLBLL_R_X73Y107_SLICE_X110Y107_C4 = CLBLL_R_X73Y107_SLICE_X111Y107_CQ;
  assign CLBLL_R_X73Y107_SLICE_X110Y107_C5 = CLBLM_L_X72Y107_SLICE_X108Y107_CQ;
  assign CLBLL_R_X73Y107_SLICE_X110Y107_C6 = CLBLL_R_X71Y107_SLICE_X106Y107_C5Q;
  assign CLBLL_R_X73Y107_SLICE_X110Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_D5 = 1'b1;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_D6 = 1'b1;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X73Y107_SLICE_X110Y107_D1 = CLBLM_L_X72Y106_SLICE_X108Y106_AQ;
  assign CLBLL_R_X73Y107_SLICE_X110Y107_D2 = CLBLM_L_X72Y107_SLICE_X109Y107_BQ;
  assign CLBLL_R_X73Y107_SLICE_X110Y107_D3 = CLBLM_L_X74Y107_SLICE_X112Y107_AQ;
  assign CLBLL_R_X73Y107_SLICE_X110Y107_D4 = CLBLL_R_X73Y107_SLICE_X110Y107_CO6;
  assign CLBLL_R_X73Y107_SLICE_X110Y107_D5 = CLBLL_R_X73Y107_SLICE_X111Y107_DQ;
  assign CLBLL_R_X73Y107_SLICE_X110Y107_D6 = CLBLM_L_X72Y107_SLICE_X109Y107_BO5;
  assign CLBLL_R_X73Y107_SLICE_X110Y107_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X73Y107_SLICE_X111Y107_A1 = CLBLM_L_X72Y108_SLICE_X108Y108_BO5;
  assign CLBLL_R_X73Y107_SLICE_X111Y107_A2 = CLBLL_R_X73Y107_SLICE_X111Y107_BQ;
  assign CLBLL_R_X73Y107_SLICE_X111Y107_A3 = CLBLM_L_X72Y108_SLICE_X109Y108_CO5;
  assign CLBLL_R_X73Y107_SLICE_X111Y107_A4 = CLBLL_R_X73Y107_SLICE_X111Y107_AQ;
  assign CLBLL_R_X73Y107_SLICE_X111Y107_A5 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLL_R_X73Y107_SLICE_X111Y107_A6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y107_SLICE_X111Y107_B1 = CLBLM_L_X74Y107_SLICE_X112Y107_DQ;
  assign CLBLL_R_X73Y107_SLICE_X111Y107_B2 = CLBLL_R_X73Y107_SLICE_X111Y107_BQ;
  assign CLBLL_R_X73Y107_SLICE_X111Y107_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y107_SLICE_X111Y107_B4 = CLBLM_L_X72Y108_SLICE_X108Y108_BO6;
  assign CLBLL_R_X73Y107_SLICE_X111Y107_B5 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLL_R_X73Y107_SLICE_X111Y107_B6 = CLBLM_L_X72Y108_SLICE_X109Y108_A5Q;
  assign CLBLL_R_X73Y107_SLICE_X111Y107_C1 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLL_R_X73Y107_SLICE_X111Y107_C2 = CLBLL_R_X73Y107_SLICE_X111Y107_CQ;
  assign CLBLL_R_X73Y107_SLICE_X111Y107_C3 = CLBLM_L_X74Y107_SLICE_X113Y107_AQ;
  assign CLBLL_R_X73Y107_SLICE_X111Y107_C4 = CLBLM_L_X72Y108_SLICE_X109Y108_A5Q;
  assign CLBLL_R_X73Y107_SLICE_X111Y107_C5 = CLBLM_L_X72Y108_SLICE_X108Y108_BO5;
  assign CLBLL_R_X73Y107_SLICE_X111Y107_C6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y107_SLICE_X111Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOB33_X0Y69_IOB_X0Y70_O = CLBLL_R_X75Y127_SLICE_X115Y127_AQ;
  assign LIOB33_X0Y69_IOB_X0Y69_O = CLBLM_L_X60Y92_SLICE_X90Y92_AQ;
  assign CLBLL_R_X73Y107_SLICE_X111Y107_D1 = CLBLM_L_X72Y108_SLICE_X109Y108_BO6;
  assign CLBLL_R_X73Y107_SLICE_X111Y107_D2 = CLBLL_R_X73Y107_SLICE_X111Y107_AQ;
  assign CLBLL_R_X73Y107_SLICE_X111Y107_D3 = CLBLL_R_X73Y107_SLICE_X111Y107_DQ;
  assign CLBLL_R_X73Y107_SLICE_X111Y107_D4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y107_SLICE_X111Y107_D5 = CLBLM_L_X72Y108_SLICE_X108Y108_BO5;
  assign CLBLL_R_X73Y107_SLICE_X111Y107_D6 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLL_R_X73Y107_SLICE_X111Y107_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign LIOB33_X0Y79_IOB_X0Y80_O = CLBLM_L_X60Y92_SLICE_X90Y92_BQ;
  assign RIOB33_X105Y157_IOB_X1Y158_O = 1'b1;
  assign RIOB33_X105Y157_IOB_X1Y157_O = 1'b1;
  assign CLBLM_R_X103Y75_SLICE_X162Y75_C4 = 1'b1;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_A1 = CLBLL_R_X73Y126_SLICE_X110Y126_A5Q;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_A3 = CLBLL_R_X71Y127_SLICE_X107Y127_AQ;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_A4 = CLBLL_R_X71Y126_SLICE_X106Y126_CO6;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_A5 = CLBLL_R_X73Y126_SLICE_X110Y126_BQ;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_A6 = CLBLM_L_X72Y126_SLICE_X109Y126_AQ;
  assign CLBLM_L_X72Y113_SLICE_X109Y113_D3 = 1'b1;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_B1 = CLBLL_R_X73Y126_SLICE_X110Y126_A5Q;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_B2 = CLBLM_L_X72Y126_SLICE_X109Y126_BQ;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_B3 = CLBLM_L_X72Y126_SLICE_X109Y126_AQ;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_B4 = CLBLL_R_X73Y128_SLICE_X110Y128_AQ;
  assign CLBLM_L_X72Y113_SLICE_X109Y113_D4 = 1'b1;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_B5 = CLBLL_R_X71Y126_SLICE_X106Y126_CO6;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_B6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y113_SLICE_X109Y113_D5 = 1'b1;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_C2 = CLBLM_L_X72Y126_SLICE_X109Y126_CQ;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_C3 = 1'b1;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_C4 = CLBLM_L_X72Y126_SLICE_X109Y126_BQ;
  assign CLBLM_L_X72Y113_SLICE_X109Y113_D6 = 1'b1;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_C5 = CLBLM_L_X72Y126_SLICE_X109Y126_DO6;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_C6 = CLBLL_R_X73Y128_SLICE_X110Y128_AQ;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X67Y115_SLICE_X100Y115_B4 = 1'b1;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_D1 = CLBLL_R_X71Y126_SLICE_X106Y126_CO6;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_D2 = 1'b1;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_D3 = 1'b1;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_D4 = 1'b1;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_D5 = CLBLM_L_X72Y126_SLICE_X109Y126_AQ;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_D6 = CLBLL_R_X73Y126_SLICE_X110Y126_A5Q;
  assign CLBLL_R_X71Y107_SLICE_X107Y107_D5 = CLBLL_R_X71Y107_SLICE_X106Y107_C5Q;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X103Y75_SLICE_X162Y75_C6 = 1'b1;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_A1 = CLBLM_L_X64Y102_SLICE_X96Y102_A5Q;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_A2 = CLBLM_L_X64Y102_SLICE_X96Y102_BO6;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_A3 = CLBLM_L_X62Y102_SLICE_X93Y102_AQ;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_A4 = CLBLM_L_X62Y102_SLICE_X93Y102_DQ;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_A6 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_A1 = CLBLL_R_X75Y127_SLICE_X115Y127_DQ;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_A2 = CLBLM_L_X72Y126_SLICE_X108Y126_CO6;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_A3 = CLBLM_L_X72Y126_SLICE_X108Y126_AQ;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_B1 = CLBLM_R_X63Y102_SLICE_X95Y102_AO5;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_B2 = CLBLM_L_X62Y102_SLICE_X93Y102_BQ;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_B4 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_B5 = CLBLM_R_X63Y102_SLICE_X95Y102_BQ;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_B6 = CLBLM_R_X63Y102_SLICE_X94Y102_DO6;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_B1 = CLBLM_L_X72Y126_SLICE_X108Y126_DO6;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_B2 = CLBLM_L_X72Y126_SLICE_X108Y126_BQ;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_B3 = CLBLM_L_X72Y126_SLICE_X108Y126_AQ;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_C2 = CLBLM_L_X62Y102_SLICE_X93Y102_CQ;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_C3 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_C4 = CLBLM_L_X62Y103_SLICE_X93Y103_CQ;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_C5 = CLBLM_L_X64Y102_SLICE_X96Y102_BO6;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_C6 = CLBLM_R_X63Y102_SLICE_X94Y102_DO5;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_C1 = CLBLM_L_X70Y123_SLICE_X104Y123_AQ;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_C2 = CLBLL_R_X71Y126_SLICE_X107Y126_BQ;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_C3 = CLBLL_R_X71Y126_SLICE_X107Y126_AQ;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_C4 = CLBLM_L_X70Y125_SLICE_X105Y125_AQ;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_C5 = CLBLL_R_X71Y126_SLICE_X106Y126_AQ;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_C6 = CLBLM_L_X70Y124_SLICE_X105Y124_BO6;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_D1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_D2 = CLBLM_L_X62Y102_SLICE_X93Y102_CQ;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_D3 = CLBLM_L_X62Y102_SLICE_X93Y102_DQ;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_D4 = CLBLM_R_X63Y103_SLICE_X94Y103_AO5;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_D5 = CLBLM_L_X64Y102_SLICE_X96Y102_BO6;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_D6 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_D1 = CLBLM_L_X72Y127_SLICE_X108Y127_AQ;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_D2 = CLBLM_L_X72Y127_SLICE_X108Y127_A5Q;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_D3 = 1'b1;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_D4 = CLBLM_L_X72Y126_SLICE_X108Y126_CO6;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_A1 = CLBLM_R_X63Y102_SLICE_X94Y102_DO6;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_A2 = CLBLM_R_X63Y103_SLICE_X94Y103_AO6;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_A3 = CLBLM_L_X62Y102_SLICE_X92Y102_AQ;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_A4 = CLBLM_L_X62Y102_SLICE_X93Y102_BQ;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_A6 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_B1 = CLBLM_R_X63Y102_SLICE_X94Y102_DO6;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_B2 = CLBLM_L_X62Y102_SLICE_X92Y102_BQ;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_B3 = CLBLM_L_X62Y102_SLICE_X92Y102_AQ;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_B4 = CLBLM_R_X63Y102_SLICE_X94Y102_DO5;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y108_SLICE_X110Y108_A1 = CLBLM_L_X72Y107_SLICE_X109Y107_DO6;
  assign CLBLL_R_X73Y108_SLICE_X110Y108_A2 = CLBLL_R_X73Y108_SLICE_X110Y108_A5Q;
  assign CLBLL_R_X73Y108_SLICE_X110Y108_A3 = CLBLL_R_X73Y113_SLICE_X110Y113_AQ;
  assign CLBLL_R_X73Y108_SLICE_X110Y108_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y108_SLICE_X110Y108_A5 = CLBLM_L_X72Y107_SLICE_X108Y107_CQ;
  assign CLBLL_R_X73Y108_SLICE_X110Y108_A6 = 1'b1;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_B6 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_C4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_C1 = CLBLM_L_X62Y102_SLICE_X92Y102_BQ;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_C6 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLL_R_X73Y108_SLICE_X110Y108_B1 = CLBLM_L_X72Y109_SLICE_X108Y109_BO6;
  assign CLBLL_R_X73Y108_SLICE_X110Y108_B2 = CLBLL_R_X73Y108_SLICE_X110Y108_BQ;
  assign CLBLL_R_X73Y108_SLICE_X110Y108_B3 = CLBLM_L_X72Y108_SLICE_X109Y108_BO5;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X73Y108_SLICE_X110Y108_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y108_SLICE_X110Y108_B5 = CLBLL_R_X73Y107_SLICE_X110Y107_BQ;
  assign CLBLL_R_X73Y108_SLICE_X110Y108_B6 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLL_R_X73Y108_SLICE_X110Y108_C1 = 1'b1;
  assign CLBLL_R_X73Y108_SLICE_X110Y108_C2 = 1'b1;
  assign CLBLL_R_X73Y108_SLICE_X110Y108_C3 = 1'b1;
  assign CLBLL_R_X73Y108_SLICE_X110Y108_C4 = 1'b1;
  assign CLBLL_R_X73Y108_SLICE_X110Y108_C5 = 1'b1;
  assign CLBLL_R_X73Y108_SLICE_X110Y108_C6 = 1'b1;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_D1 = CLBLM_L_X62Y100_SLICE_X92Y100_AQ;
  assign CLBLL_R_X73Y108_SLICE_X110Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_D2 = CLBLM_R_X63Y102_SLICE_X94Y102_BQ;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_D3 = CLBLM_L_X64Y101_SLICE_X96Y101_BQ;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_D4 = CLBLM_L_X64Y101_SLICE_X96Y101_B5Q;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_D5 = CLBLM_L_X62Y103_SLICE_X92Y103_A5Q;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_D6 = CLBLM_L_X62Y102_SLICE_X93Y102_BQ;
  assign CLBLL_R_X73Y108_SLICE_X110Y108_D1 = 1'b1;
  assign CLBLL_R_X73Y108_SLICE_X110Y108_D2 = 1'b1;
  assign CLBLL_R_X73Y108_SLICE_X110Y108_D3 = 1'b1;
  assign CLBLL_R_X73Y108_SLICE_X110Y108_D4 = 1'b1;
  assign CLBLL_R_X73Y108_SLICE_X110Y108_D5 = 1'b1;
  assign CLBLL_R_X73Y108_SLICE_X110Y108_D6 = 1'b1;
  assign CLBLL_R_X73Y108_SLICE_X110Y108_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_D5 = 1'b1;
  assign CLBLM_L_X76Y111_SLICE_X116Y111_C1 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X108Y113_BX = CLBLM_L_X70Y113_SLICE_X104Y113_CQ;
  assign CLBLL_R_X73Y108_SLICE_X111Y108_A1 = 1'b1;
  assign CLBLL_R_X73Y108_SLICE_X111Y108_A2 = 1'b1;
  assign CLBLL_R_X73Y108_SLICE_X111Y108_A3 = 1'b1;
  assign CLBLL_R_X73Y108_SLICE_X111Y108_A4 = 1'b1;
  assign CLBLL_R_X73Y108_SLICE_X111Y108_A5 = 1'b1;
  assign CLBLL_R_X73Y108_SLICE_X111Y108_A6 = 1'b1;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_D6 = 1'b1;
  assign CLBLM_L_X76Y111_SLICE_X116Y111_C2 = 1'b1;
  assign LIOB33_X0Y71_IOB_X0Y71_O = CLBLM_L_X60Y94_SLICE_X90Y94_AQ;
  assign CLBLL_R_X73Y108_SLICE_X111Y108_B1 = 1'b1;
  assign CLBLL_R_X73Y108_SLICE_X111Y108_B2 = 1'b1;
  assign CLBLL_R_X73Y108_SLICE_X111Y108_B3 = 1'b1;
  assign CLBLL_R_X73Y108_SLICE_X111Y108_B4 = 1'b1;
  assign CLBLL_R_X73Y108_SLICE_X111Y108_B5 = 1'b1;
  assign CLBLL_R_X73Y108_SLICE_X111Y108_B6 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X108Y113_C5 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X108Y113_C6 = 1'b1;
  assign CLBLL_R_X73Y108_SLICE_X111Y108_C1 = 1'b1;
  assign CLBLL_R_X73Y108_SLICE_X111Y108_C2 = 1'b1;
  assign CLBLL_R_X73Y108_SLICE_X111Y108_C3 = 1'b1;
  assign CLBLL_R_X73Y108_SLICE_X111Y108_C4 = 1'b1;
  assign CLBLL_R_X73Y108_SLICE_X111Y108_C5 = 1'b1;
  assign CLBLL_R_X73Y108_SLICE_X111Y108_C6 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_A1 = CLBLL_R_X75Y123_SLICE_X115Y123_DO6;
  assign CLBLM_L_X78Y130_SLICE_X121Y130_A2 = 1'b1;
  assign CLBLM_L_X76Y111_SLICE_X116Y111_C3 = 1'b1;
  assign CLBLL_R_X73Y108_SLICE_X111Y108_D1 = 1'b1;
  assign CLBLL_R_X73Y108_SLICE_X111Y108_D2 = 1'b1;
  assign CLBLL_R_X73Y108_SLICE_X111Y108_D3 = 1'b1;
  assign CLBLL_R_X73Y108_SLICE_X111Y108_D4 = 1'b1;
  assign CLBLL_R_X73Y108_SLICE_X111Y108_D5 = 1'b1;
  assign CLBLL_R_X73Y108_SLICE_X111Y108_D6 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X108Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X78Y130_SLICE_X121Y130_A3 = 1'b1;
  assign RIOB33_X105Y159_IOB_X1Y159_O = 1'b1;
  assign RIOB33_X105Y159_IOB_X1Y160_O = CLBLM_L_X74Y120_SLICE_X112Y120_AO6;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_A2 = CLBLL_R_X75Y124_SLICE_X114Y124_BQ;
  assign CLBLM_L_X76Y111_SLICE_X116Y111_C4 = 1'b1;
  assign CLBLM_L_X78Y130_SLICE_X121Y130_A4 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_A3 = CLBLM_L_X76Y125_SLICE_X117Y125_AQ;
  assign CLBLM_L_X76Y111_SLICE_X116Y111_C5 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X108Y113_D4 = 1'b1;
  assign CLBLM_L_X78Y130_SLICE_X121Y130_A5 = 1'b1;
  assign CLBLM_L_X72Y113_SLICE_X108Y113_D5 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_A4 = CLBLL_R_X73Y125_SLICE_X111Y125_AQ;
  assign CLBLM_L_X76Y111_SLICE_X116Y111_C6 = 1'b1;
  assign CLBLM_L_X78Y130_SLICE_X121Y130_A6 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_A5 = CLBLL_R_X75Y124_SLICE_X114Y124_AQ;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_A1 = CLBLL_R_X73Y127_SLICE_X111Y127_CQ;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_A2 = CLBLL_R_X73Y126_SLICE_X110Y126_A5Q;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_A3 = CLBLM_L_X72Y127_SLICE_X109Y127_BO6;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_A4 = CLBLL_R_X73Y127_SLICE_X110Y127_AQ;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_A5 = CLBLM_L_X72Y126_SLICE_X109Y126_AQ;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_A6 = CLBLM_L_X72Y127_SLICE_X109Y127_CO6;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_AX = CLBLL_R_X75Y127_SLICE_X114Y127_AQ;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_B1 = CLBLL_R_X73Y127_SLICE_X110Y127_DQ;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_B2 = CLBLL_R_X73Y126_SLICE_X110Y126_A5Q;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_B3 = CLBLM_L_X72Y126_SLICE_X109Y126_AQ;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_B4 = CLBLL_R_X73Y127_SLICE_X111Y127_AQ;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_B5 = 1'b1;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_B6 = CLBLL_R_X71Y127_SLICE_X107Y127_AQ;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_A6 = CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_D1 = CLBLM_L_X72Y122_SLICE_X108Y122_AO6;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_BX = CLBLM_L_X72Y128_SLICE_X108Y128_A5Q;
  assign CLBLM_R_X103Y75_SLICE_X163Y75_A6 = 1'b1;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_C1 = CLBLM_L_X72Y126_SLICE_X109Y126_AQ;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_C2 = CLBLL_R_X73Y126_SLICE_X110Y126_A5Q;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_C3 = 1'b1;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_C4 = CLBLL_R_X71Y127_SLICE_X107Y127_AQ;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_C5 = CLBLL_R_X73Y127_SLICE_X110Y127_BQ;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_C6 = CLBLL_R_X75Y127_SLICE_X114Y127_BQ;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_CE = CLBLM_L_X76Y109_SLICE_X116Y109_AO6;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_T1 = 1'b1;
  assign CLBLM_R_X103Y75_SLICE_X163Y75_AX = CLBLM_R_X103Y76_SLICE_X162Y76_AQ;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_D1 = 1'b1;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_D2 = 1'b1;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_D3 = 1'b1;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_D4 = 1'b1;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_D5 = 1'b1;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_D6 = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_D1 = CLBLM_L_X70Y134_SLICE_X104Y134_CO5;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X103Y75_SLICE_X163Y75_B1 = 1'b1;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_A1 = CLBLM_L_X62Y103_SLICE_X93Y103_AQ;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_A2 = CLBLM_L_X62Y103_SLICE_X93Y103_BQ;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_A3 = CLBLM_L_X64Y102_SLICE_X96Y102_BO6;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_A4 = CLBLM_R_X63Y102_SLICE_X95Y102_AO5;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_A6 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_A2 = CLBLM_L_X72Y126_SLICE_X108Y126_CO6;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_A3 = CLBLM_L_X72Y127_SLICE_X108Y127_AQ;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_B1 = CLBLM_L_X64Y102_SLICE_X96Y102_A5Q;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_B2 = CLBLM_L_X62Y103_SLICE_X93Y103_BQ;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_B3 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_B4 = CLBLM_L_X62Y103_SLICE_X93Y103_DQ;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_B6 = CLBLM_R_X63Y103_SLICE_X95Y103_BO6;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_AX = CLBLM_L_X72Y127_SLICE_X108Y127_BO5;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_B1 = CLBLM_L_X72Y128_SLICE_X108Y128_A5Q;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_B2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_C1 = CLBLM_L_X64Y102_SLICE_X96Y102_BO6;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_C2 = CLBLM_L_X62Y103_SLICE_X93Y103_CQ;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_C3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_C4 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_C5 = CLBLM_L_X62Y103_SLICE_X93Y103_AQ;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_C6 = CLBLM_R_X63Y103_SLICE_X94Y103_AO6;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_C1 = 1'b1;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_C2 = CLBLM_L_X72Y127_SLICE_X108Y127_CQ;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_C3 = CLBLM_L_X72Y126_SLICE_X108Y126_CO6;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_C4 = CLBLM_L_X72Y127_SLICE_X108Y127_A5Q;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_C5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_C6 = CLBLM_L_X74Y127_SLICE_X112Y127_BO6;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_D1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_D2 = CLBLM_R_X63Y103_SLICE_X95Y103_BO6;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_D3 = CLBLM_L_X62Y103_SLICE_X93Y103_DQ;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_D4 = CLBLM_R_X63Y103_SLICE_X94Y103_AO5;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_D5 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_D6 = CLBLM_L_X62Y103_SLICE_X92Y103_BQ;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_D1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_D2 = CLBLM_L_X72Y127_SLICE_X108Y127_AQ;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_D3 = CLBLM_L_X72Y127_SLICE_X108Y127_DQ;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_D4 = CLBLM_L_X72Y127_SLICE_X108Y127_A5Q;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_A1 = CLBLM_R_X63Y103_SLICE_X95Y103_AQ;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_A2 = CLBLM_R_X63Y103_SLICE_X94Y103_AO6;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_A3 = CLBLM_L_X62Y103_SLICE_X92Y103_AQ;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_A4 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_A6 = CLBLM_R_X63Y103_SLICE_X95Y103_BO6;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X103Y75_SLICE_X163Y75_C1 = 1'b1;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_AX = CLBLM_R_X63Y101_SLICE_X94Y101_AQ;
  assign CLBLM_R_X103Y75_SLICE_X163Y75_C2 = 1'b1;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_B1 = CLBLM_L_X62Y103_SLICE_X92Y103_AQ;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_B2 = CLBLM_L_X62Y103_SLICE_X92Y103_BQ;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_B3 = CLBLM_R_X63Y102_SLICE_X94Y102_DO5;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_B4 = CLBLM_R_X63Y103_SLICE_X95Y103_BO6;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_B6 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLL_R_X73Y109_SLICE_X110Y109_A1 = CLBLM_L_X72Y109_SLICE_X109Y109_A5Q;
  assign CLBLL_R_X73Y109_SLICE_X110Y109_A2 = CLBLM_L_X72Y109_SLICE_X108Y109_AQ;
  assign CLBLL_R_X73Y109_SLICE_X110Y109_A3 = CLBLM_L_X72Y116_SLICE_X108Y116_AQ;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_BX = CLBLM_L_X62Y103_SLICE_X92Y103_A5Q;
  assign CLBLL_R_X73Y109_SLICE_X110Y109_A4 = CLBLM_L_X72Y109_SLICE_X109Y109_C5Q;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_C1 = CLBLM_L_X64Y101_SLICE_X96Y101_B5Q;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_C2 = CLBLM_L_X62Y103_SLICE_X92Y103_AQ;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_C3 = CLBLM_L_X64Y101_SLICE_X96Y101_A5Q;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_C4 = CLBLM_L_X62Y103_SLICE_X92Y103_A5Q;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_C5 = 1'b1;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_C6 = CLBLM_L_X64Y101_SLICE_X96Y101_BQ;
  assign CLBLL_R_X73Y109_SLICE_X110Y109_B1 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X110Y109_B2 = 1'b1;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X73Y109_SLICE_X110Y109_B3 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X110Y109_B4 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X110Y109_B5 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X110Y109_B6 = 1'b1;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_D1 = 1'b1;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_D2 = 1'b1;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_D3 = 1'b1;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_D4 = 1'b1;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_D5 = 1'b1;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_D6 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X110Y109_C5 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X110Y109_C6 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X110Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X73Y109_SLICE_X110Y109_D1 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X110Y109_D2 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X110Y109_D3 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X110Y109_D4 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X110Y109_D5 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X110Y109_D6 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X110Y109_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y134_SLICE_X109Y134_C6 = 1'b1;
  assign LIOB33_X0Y73_IOB_X0Y74_O = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign LIOB33_X0Y73_IOB_X0Y73_O = CLBLM_L_X62Y105_SLICE_X93Y105_A5Q;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_B1 = 1'b1;
  assign CLBLM_L_X78Y130_SLICE_X121Y130_B3 = 1'b1;
  assign CLBLM_R_X103Y75_SLICE_X163Y75_D1 = 1'b1;
  assign CLBLM_R_X103Y75_SLICE_X163Y75_D2 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X111Y109_A1 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X111Y109_A2 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X111Y109_A3 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X111Y109_A4 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X111Y109_A5 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X111Y109_A6 = 1'b1;
  assign CLBLM_R_X103Y75_SLICE_X163Y75_D3 = 1'b1;
  assign LIOI3_X0Y51_OLOGIC_X0Y52_T1 = 1'b1;
  assign CLBLM_R_X103Y75_SLICE_X163Y75_D4 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X111Y109_B1 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X111Y109_B2 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X111Y109_B3 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X111Y109_B4 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X111Y109_B5 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X111Y109_B6 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_B2 = CLBLM_L_X74Y127_SLICE_X112Y127_AQ;
  assign CLBLM_L_X78Y130_SLICE_X121Y130_B4 = 1'b1;
  assign CLBLM_R_X103Y75_SLICE_X163Y75_D5 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X111Y109_C1 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X111Y109_C2 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X111Y109_C3 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X111Y109_C4 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X111Y109_C5 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X111Y109_C6 = 1'b1;
  assign CLBLM_R_X103Y75_SLICE_X163Y75_D6 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X111Y109_D1 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X111Y109_D2 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X111Y109_D3 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X111Y109_D4 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X111Y109_D5 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X111Y109_D6 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_B3 = CLBLM_L_X74Y125_SLICE_X112Y125_AQ;
  assign CLBLM_L_X78Y130_SLICE_X121Y130_B5 = 1'b1;
  assign CLBLM_R_X103Y75_SLICE_X163Y75_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y134_SLICE_X109Y134_D6 = 1'b1;
  assign CLBLM_R_X103Y75_SLICE_X162Y75_A1 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_B4 = CLBLL_R_X73Y123_SLICE_X110Y123_CQ;
  assign CLBLM_R_X103Y75_SLICE_X162Y75_A2 = 1'b1;
  assign CLBLM_R_X103Y75_SLICE_X162Y75_A3 = CLBLM_R_X103Y75_SLICE_X162Y75_AQ;
  assign CLBLM_L_X76Y111_SLICE_X116Y111_D1 = 1'b1;
  assign CLBLM_R_X103Y75_SLICE_X162Y75_A4 = CLBLM_R_X103Y75_SLICE_X163Y75_BQ;
  assign CLBLM_R_X103Y75_SLICE_X162Y75_A5 = CLBLM_R_X103Y76_SLICE_X162Y76_AQ;
  assign CLBLM_R_X103Y75_SLICE_X162Y75_A6 = CLBLM_R_X103Y75_SLICE_X162Y75_CQ;
  assign CLBLM_L_X76Y111_SLICE_X116Y111_D2 = 1'b1;
  assign CLBLM_L_X72Y134_SLICE_X108Y134_A4 = CLBLL_R_X73Y132_SLICE_X110Y132_AO6;
  assign CLBLM_R_X103Y75_SLICE_X162Y75_AX = CLBLM_R_X103Y75_SLICE_X163Y75_AQ;
  assign CLBLL_R_X75Y121_SLICE_X114Y121_A1 = CLBLM_L_X76Y123_SLICE_X116Y123_BQ;
  assign CLBLL_R_X75Y121_SLICE_X114Y121_A2 = CLBLL_R_X75Y121_SLICE_X114Y121_BQ;
  assign CLBLL_R_X75Y121_SLICE_X114Y121_A3 = CLBLL_R_X75Y123_SLICE_X115Y123_AQ;
  assign CLBLL_R_X75Y121_SLICE_X114Y121_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y121_SLICE_X114Y121_A5 = CLBLM_L_X70Y105_SLICE_X105Y105_AQ;
  assign CLBLL_R_X75Y121_SLICE_X114Y121_A6 = 1'b1;
  assign CLBLM_R_X103Y75_SLICE_X162Y75_B2 = 1'b1;
  assign CLBLM_L_X76Y111_SLICE_X116Y111_D3 = 1'b1;
  assign CLBLL_R_X75Y121_SLICE_X114Y121_B1 = CLBLM_L_X74Y123_SLICE_X113Y123_CO5;
  assign CLBLL_R_X75Y121_SLICE_X114Y121_B2 = CLBLL_R_X75Y121_SLICE_X114Y121_BQ;
  assign CLBLL_R_X75Y121_SLICE_X114Y121_B3 = CLBLL_R_X75Y123_SLICE_X115Y123_AQ;
  assign CLBLL_R_X75Y121_SLICE_X114Y121_B4 = CLBLL_R_X75Y122_SLICE_X114Y122_AQ;
  assign CLBLL_R_X75Y121_SLICE_X114Y121_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y121_SLICE_X114Y121_B6 = CLBLL_R_X75Y121_SLICE_X114Y121_CO6;
  assign CLBLM_R_X103Y75_SLICE_X162Y75_B3 = 1'b1;
  assign CLBLM_R_X103Y75_SLICE_X162Y75_B4 = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_D1 = CLBLM_R_X65Y106_SLICE_X99Y106_DQ;
  assign CLBLL_R_X75Y121_SLICE_X114Y121_C1 = CLBLL_R_X75Y123_SLICE_X115Y123_AQ;
  assign CLBLL_R_X75Y121_SLICE_X114Y121_C2 = CLBLM_L_X76Y123_SLICE_X116Y123_BQ;
  assign CLBLL_R_X75Y121_SLICE_X114Y121_C3 = CLBLM_L_X74Y123_SLICE_X113Y123_DQ;
  assign CLBLL_R_X75Y121_SLICE_X114Y121_C4 = 1'b1;
  assign CLBLL_R_X75Y121_SLICE_X114Y121_C5 = CLBLL_R_X75Y122_SLICE_X114Y122_CQ;
  assign CLBLL_R_X75Y121_SLICE_X114Y121_C6 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_A1 = CLBLM_L_X74Y134_SLICE_X112Y134_DQ;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_A2 = CLBLM_L_X72Y123_SLICE_X108Y123_BQ;
  assign CLBLL_R_X75Y121_SLICE_X114Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_A3 = CLBLM_L_X72Y128_SLICE_X109Y128_AQ;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_A4 = CLBLL_R_X77Y128_SLICE_X119Y128_AQ;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_A6 = 1'b1;
  assign CLBLL_R_X75Y121_SLICE_X114Y121_D1 = 1'b1;
  assign CLBLL_R_X75Y121_SLICE_X114Y121_D2 = 1'b1;
  assign CLBLL_R_X75Y121_SLICE_X114Y121_D3 = 1'b1;
  assign CLBLL_R_X75Y121_SLICE_X114Y121_D4 = 1'b1;
  assign CLBLL_R_X75Y121_SLICE_X114Y121_D5 = 1'b1;
  assign CLBLL_R_X75Y121_SLICE_X114Y121_D6 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_B1 = 1'b1;
  assign CLBLL_R_X75Y121_SLICE_X114Y121_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_B3 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_B4 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_B5 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_B6 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_C1 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_C2 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_C3 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_C4 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_C5 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_C6 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_D1 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_D2 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_D3 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_D4 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_D5 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_D6 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X82Y130_SLICE_X129Y130_B1 = 1'b1;
  assign CLBLL_R_X75Y121_SLICE_X115Y121_A1 = 1'b1;
  assign CLBLL_R_X75Y121_SLICE_X115Y121_A2 = 1'b1;
  assign CLBLL_R_X75Y121_SLICE_X115Y121_A3 = 1'b1;
  assign CLBLL_R_X75Y121_SLICE_X115Y121_A4 = 1'b1;
  assign CLBLL_R_X75Y121_SLICE_X115Y121_A5 = 1'b1;
  assign CLBLL_R_X75Y121_SLICE_X115Y121_A6 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_A1 = CLBLM_L_X74Y128_SLICE_X112Y128_CQ;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_A2 = CLBLM_L_X74Y127_SLICE_X112Y127_AO6;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_C1 = 1'b1;
  assign CLBLL_R_X75Y121_SLICE_X115Y121_B1 = 1'b1;
  assign CLBLL_R_X75Y121_SLICE_X115Y121_B2 = 1'b1;
  assign CLBLL_R_X75Y121_SLICE_X115Y121_B3 = 1'b1;
  assign CLBLL_R_X75Y121_SLICE_X115Y121_B4 = 1'b1;
  assign CLBLL_R_X75Y121_SLICE_X115Y121_B5 = 1'b1;
  assign CLBLL_R_X75Y121_SLICE_X115Y121_B6 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_A6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_AX = CLBLM_L_X72Y128_SLICE_X108Y128_BO6;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_B1 = 1'b1;
  assign CLBLL_R_X75Y121_SLICE_X115Y121_C1 = 1'b1;
  assign CLBLL_R_X75Y121_SLICE_X115Y121_C2 = 1'b1;
  assign CLBLL_R_X75Y121_SLICE_X115Y121_C3 = 1'b1;
  assign CLBLL_R_X75Y121_SLICE_X115Y121_C4 = 1'b1;
  assign CLBLL_R_X75Y121_SLICE_X115Y121_C5 = 1'b1;
  assign CLBLL_R_X75Y121_SLICE_X115Y121_C6 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_C1 = CLBLM_L_X72Y127_SLICE_X108Y127_AQ;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_C2 = CLBLM_L_X72Y128_SLICE_X108Y128_CQ;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_C3 = CLBLM_L_X72Y126_SLICE_X108Y126_CO6;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_C4 = CLBLM_L_X72Y128_SLICE_X108Y128_A5Q;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_C5 = CLBLM_L_X72Y127_SLICE_X108Y127_CQ;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_C6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X75Y121_SLICE_X115Y121_D1 = 1'b1;
  assign CLBLL_R_X75Y121_SLICE_X115Y121_D2 = 1'b1;
  assign CLBLL_R_X75Y121_SLICE_X115Y121_D3 = 1'b1;
  assign CLBLL_R_X75Y121_SLICE_X115Y121_D4 = 1'b1;
  assign CLBLL_R_X75Y121_SLICE_X115Y121_D5 = 1'b1;
  assign CLBLL_R_X75Y121_SLICE_X115Y121_D6 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_D1 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_D2 = CLBLM_L_X72Y128_SLICE_X108Y128_CQ;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_D3 = CLBLM_L_X74Y128_SLICE_X113Y128_CQ;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_D4 = CLBLM_L_X72Y128_SLICE_X108Y128_DQ;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_D5 = CLBLM_L_X72Y128_SLICE_X108Y128_BO5;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_D6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X67Y115_SLICE_X100Y115_D5 = 1'b1;
  assign CLBLM_L_X82Y130_SLICE_X129Y130_C3 = 1'b1;
  assign CLBLM_L_X82Y130_SLICE_X129Y130_C5 = 1'b1;
  assign CLBLM_L_X82Y130_SLICE_X129Y130_C6 = 1'b1;
  assign CLBLM_R_X67Y115_SLICE_X100Y115_D6 = 1'b1;
  assign LIOB33_X0Y75_IOB_X0Y75_O = CLBLM_L_X60Y101_SLICE_X90Y101_BQ;
  assign LIOB33_X0Y75_IOB_X0Y76_O = CLBLM_L_X60Y99_SLICE_X90Y99_AQ;
  assign CLBLM_R_X103Y75_SLICE_X162Y75_D6 = 1'b1;
  assign LIOB33_X0Y113_IOB_X0Y114_O = CLBLL_R_X71Y124_SLICE_X106Y124_AQ;
  assign RIOB33_X105Y163_IOB_X1Y164_O = CLBLL_R_X77Y124_SLICE_X118Y124_AO6;
  assign RIOB33_X105Y163_IOB_X1Y163_O = 1'b0;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_B3 = CLBLL_R_X77Y129_SLICE_X119Y129_BQ;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_B5 = CLBLL_R_X73Y132_SLICE_X111Y132_AO6;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_B6 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_C3 = CLBLM_L_X76Y125_SLICE_X117Y125_BQ;
  assign CLBLM_R_X67Y115_SLICE_X100Y115_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X75Y122_SLICE_X114Y122_A1 = CLBLM_L_X74Y123_SLICE_X113Y123_CO5;
  assign CLBLL_R_X75Y122_SLICE_X114Y122_A2 = CLBLL_R_X75Y122_SLICE_X114Y122_DO6;
  assign CLBLL_R_X75Y122_SLICE_X114Y122_A3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y122_SLICE_X114Y122_A4 = CLBLM_L_X76Y123_SLICE_X116Y123_BQ;
  assign CLBLL_R_X75Y122_SLICE_X114Y122_A5 = CLBLL_R_X75Y121_SLICE_X114Y121_BQ;
  assign CLBLL_R_X75Y122_SLICE_X114Y122_A6 = CLBLL_R_X75Y123_SLICE_X115Y123_AQ;
  assign CLBLL_R_X75Y122_SLICE_X114Y122_B1 = CLBLL_R_X75Y123_SLICE_X114Y123_CO6;
  assign CLBLL_R_X75Y122_SLICE_X114Y122_B2 = CLBLL_R_X75Y122_SLICE_X114Y122_BQ;
  assign CLBLL_R_X75Y122_SLICE_X114Y122_B3 = CLBLL_R_X75Y121_SLICE_X114Y121_AO5;
  assign CLBLL_R_X75Y122_SLICE_X114Y122_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y122_SLICE_X114Y122_B5 = CLBLL_R_X75Y122_SLICE_X114Y122_CQ;
  assign CLBLL_R_X75Y122_SLICE_X114Y122_B6 = CLBLM_L_X74Y122_SLICE_X113Y122_AQ;
  assign CLBLL_R_X75Y122_SLICE_X114Y122_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y122_SLICE_X114Y122_C2 = CLBLL_R_X75Y122_SLICE_X114Y122_CQ;
  assign CLBLL_R_X75Y122_SLICE_X114Y122_C3 = CLBLM_L_X74Y123_SLICE_X113Y123_DQ;
  assign CLBLL_R_X75Y122_SLICE_X114Y122_C4 = CLBLL_R_X75Y121_SLICE_X114Y121_AO5;
  assign CLBLL_R_X75Y122_SLICE_X114Y122_C5 = CLBLL_R_X75Y123_SLICE_X114Y123_AO5;
  assign CLBLL_R_X75Y122_SLICE_X114Y122_C6 = CLBLM_L_X74Y122_SLICE_X113Y122_AQ;
  assign CLBLL_R_X75Y122_SLICE_X114Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_A1 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_A2 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_A3 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_A4 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_A5 = 1'b1;
  assign CLBLL_R_X75Y122_SLICE_X114Y122_D1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y122_SLICE_X114Y122_D2 = CLBLL_R_X75Y122_SLICE_X114Y122_AQ;
  assign CLBLL_R_X75Y122_SLICE_X114Y122_D3 = CLBLL_R_X75Y122_SLICE_X114Y122_BQ;
  assign CLBLL_R_X75Y122_SLICE_X114Y122_D4 = CLBLL_R_X75Y123_SLICE_X115Y123_AQ;
  assign CLBLL_R_X75Y122_SLICE_X114Y122_D5 = CLBLL_R_X75Y123_SLICE_X114Y123_AO5;
  assign CLBLL_R_X75Y122_SLICE_X114Y122_D6 = CLBLM_L_X74Y122_SLICE_X113Y122_AQ;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_B1 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_B2 = 1'b1;
  assign CLBLL_R_X75Y122_SLICE_X114Y122_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_B3 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_B4 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_B5 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_B6 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_C1 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_C2 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_C3 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_C4 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_C5 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_C6 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_D6 = 1'b1;
  assign CLBLM_L_X82Y130_SLICE_X128Y130_C1 = 1'b1;
  assign CLBLM_L_X82Y130_SLICE_X128Y130_C2 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_D1 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_D2 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_D3 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_D4 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_D5 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_D6 = 1'b1;
  assign CLBLL_R_X75Y122_SLICE_X115Y122_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y122_SLICE_X115Y122_A2 = CLBLL_R_X75Y122_SLICE_X115Y122_BQ;
  assign CLBLL_R_X75Y122_SLICE_X115Y122_A3 = CLBLM_L_X74Y121_SLICE_X113Y121_AQ;
  assign CLBLL_R_X75Y122_SLICE_X115Y122_A4 = CLBLL_R_X75Y123_SLICE_X114Y123_AO6;
  assign CLBLL_R_X75Y122_SLICE_X115Y122_A5 = CLBLL_R_X75Y122_SLICE_X115Y122_A5Q;
  assign CLBLL_R_X75Y122_SLICE_X115Y122_A6 = 1'b1;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_A1 = CLBLM_L_X64Y106_SLICE_X96Y106_DO6;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_A2 = CLBLM_L_X64Y105_SLICE_X96Y105_BO5;
  assign CLBLL_R_X75Y122_SLICE_X115Y122_B1 = CLBLL_R_X79Y127_SLICE_X122Y127_BQ;
  assign CLBLL_R_X75Y122_SLICE_X115Y122_B2 = CLBLL_R_X75Y122_SLICE_X115Y122_BQ;
  assign CLBLL_R_X75Y122_SLICE_X115Y122_B3 = CLBLL_R_X75Y123_SLICE_X114Y123_AO6;
  assign CLBLL_R_X75Y122_SLICE_X115Y122_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y122_SLICE_X115Y122_B5 = CLBLM_L_X76Y122_SLICE_X116Y122_AQ;
  assign CLBLL_R_X75Y122_SLICE_X115Y122_B6 = 1'b1;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_A3 = CLBLM_L_X62Y105_SLICE_X93Y105_AQ;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_A4 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y122_SLICE_X115Y122_C1 = 1'b1;
  assign CLBLL_R_X75Y122_SLICE_X115Y122_C2 = 1'b1;
  assign CLBLL_R_X75Y122_SLICE_X115Y122_C3 = 1'b1;
  assign CLBLL_R_X75Y122_SLICE_X115Y122_C4 = 1'b1;
  assign CLBLL_R_X75Y122_SLICE_X115Y122_C5 = 1'b1;
  assign CLBLL_R_X75Y122_SLICE_X115Y122_C6 = 1'b1;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_B1 = CLBLM_L_X64Y106_SLICE_X96Y106_DO6;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_B2 = CLBLM_L_X62Y105_SLICE_X93Y105_BQ;
  assign CLBLL_R_X75Y122_SLICE_X115Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_B5 = CLBLM_L_X62Y107_SLICE_X93Y107_AQ;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_B6 = CLBLM_L_X64Y105_SLICE_X96Y105_AO6;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_C1 = CLBLM_L_X64Y106_SLICE_X96Y106_DO5;
  assign CLBLL_R_X75Y122_SLICE_X115Y122_D1 = 1'b1;
  assign CLBLL_R_X75Y122_SLICE_X115Y122_D2 = 1'b1;
  assign CLBLL_R_X75Y122_SLICE_X115Y122_D3 = 1'b1;
  assign CLBLL_R_X75Y122_SLICE_X115Y122_D4 = 1'b1;
  assign CLBLL_R_X75Y122_SLICE_X115Y122_D5 = 1'b1;
  assign CLBLL_R_X75Y122_SLICE_X115Y122_D6 = 1'b1;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_C6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X75Y122_SLICE_X115Y122_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_D3 = CLBLM_L_X62Y106_SLICE_X92Y106_BQ;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_D1 = CLBLM_R_X63Y105_SLICE_X95Y105_BQ;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_D2 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_D4 = CLBLM_R_X63Y105_SLICE_X95Y105_A5Q;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_D5 = CLBLM_L_X62Y105_SLICE_X93Y105_AQ;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_D6 = CLBLM_L_X62Y107_SLICE_X93Y107_BQ;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_D1 = 1'b1;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_A1 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X110Y111_A1 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X110Y111_A2 = CLBLL_R_X73Y104_SLICE_X110Y104_AQ;
  assign CLBLL_R_X73Y111_SLICE_X110Y111_A3 = CLBLL_R_X73Y111_SLICE_X110Y111_AQ;
  assign CLBLL_R_X73Y111_SLICE_X110Y111_A4 = CLBLM_L_X72Y118_SLICE_X109Y118_A5Q;
  assign CLBLL_R_X73Y111_SLICE_X110Y111_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y111_SLICE_X110Y111_A6 = CLBLL_R_X73Y111_SLICE_X110Y111_A5Q;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_A2 = 1'b1;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_A3 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X110Y111_AX = CLBLM_L_X72Y118_SLICE_X109Y118_A5Q;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_A4 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X110Y111_B1 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X110Y111_B2 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X110Y111_B3 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X110Y111_B4 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X110Y111_B5 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X110Y111_B6 = 1'b1;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_B2 = 1'b1;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_B3 = 1'b1;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_B4 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X110Y111_C1 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X110Y111_C2 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X110Y111_C3 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X110Y111_C4 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X110Y111_C5 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X110Y111_C6 = 1'b1;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_C1 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X110Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_C2 = 1'b1;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_C3 = 1'b1;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_C4 = 1'b1;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_C5 = 1'b1;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_C6 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X110Y111_D1 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X110Y111_D2 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X110Y111_D3 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X110Y111_D4 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X110Y111_D5 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X110Y111_D6 = 1'b1;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_D4 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X110Y111_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_D1 = 1'b1;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_D2 = 1'b1;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_D3 = 1'b1;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_D5 = 1'b1;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_D6 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_B6 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X124Y132_B1 = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_T1 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X124Y132_B2 = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_D1 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X124Y132_B3 = 1'b1;
  assign CLBLM_L_X82Y130_SLICE_X128Y130_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign LIOI3_X0Y59_OLOGIC_X0Y60_D1 = CLBLM_L_X72Y106_SLICE_X108Y106_A5Q;
  assign CLBLM_L_X80Y132_SLICE_X124Y132_B4 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X111Y111_A1 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X111Y111_A2 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X111Y111_A3 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X111Y111_A4 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X111Y111_A5 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X111Y111_A6 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X124Y132_B5 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X124Y132_B6 = 1'b1;
  assign LIOI3_X0Y59_OLOGIC_X0Y60_T1 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X111Y111_B1 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X111Y111_B2 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X111Y111_B3 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X111Y111_B4 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X111Y111_B5 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X111Y111_B6 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_C3 = 1'b1;
  assign RIOI3_X105Y103_OLOGIC_X1Y104_D1 = CLBLM_L_X72Y106_SLICE_X108Y106_AQ;
  assign CLBLL_R_X73Y111_SLICE_X111Y111_C1 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X111Y111_C2 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X111Y111_C3 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X111Y111_C4 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X111Y111_C5 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X111Y111_C6 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_C5 = 1'b1;
  assign LIOI3_X0Y59_OLOGIC_X0Y59_D1 = CLBLM_L_X60Y101_SLICE_X90Y101_AQ;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_C6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y94_D1 = CLBLM_L_X62Y106_SLICE_X92Y106_AQ;
  assign RIOI3_X105Y103_OLOGIC_X1Y104_T1 = 1'b1;
  assign LIOI3_X0Y59_OLOGIC_X0Y59_T1 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X111Y111_D1 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X111Y111_D2 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X111Y111_D3 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X111Y111_D4 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X111Y111_D5 = 1'b1;
  assign CLBLL_R_X73Y111_SLICE_X111Y111_D6 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X124Y132_C1 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X124Y132_C2 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y94_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_D1 = CLBLM_L_X68Y105_SLICE_X102Y105_AQ;
  assign CLBLM_L_X80Y132_SLICE_X124Y132_C3 = 1'b1;
  assign RIOI3_X105Y103_OLOGIC_X1Y103_T1 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X80Y132_SLICE_X124Y132_C4 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y93_D1 = CLBLM_L_X62Y95_SLICE_X92Y95_BQ;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_T1 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X124Y132_C5 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X124Y132_C6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y93_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_D1 = CLBLM_L_X64Y97_SLICE_X97Y97_AQ;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_D6 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_T1 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X124Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_D4 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_D5 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_D6 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_A1 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_D5 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_A1 = CLBLM_L_X74Y123_SLICE_X113Y123_A5Q;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_A2 = CLBLL_R_X75Y123_SLICE_X114Y123_BQ;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_A3 = CLBLL_R_X75Y113_SLICE_X114Y113_AQ;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_A4 = CLBLM_L_X76Y123_SLICE_X117Y123_AQ;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_A5 = CLBLM_L_X74Y123_SLICE_X113Y123_BQ;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_A6 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X124Y132_D1 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_A3 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_B1 = CLBLM_L_X74Y123_SLICE_X113Y123_CO5;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_B2 = CLBLL_R_X75Y123_SLICE_X114Y123_BQ;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_B3 = CLBLM_L_X76Y123_SLICE_X116Y123_BQ;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_B4 = CLBLL_R_X75Y121_SLICE_X114Y121_BQ;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_B5 = CLBLL_R_X75Y123_SLICE_X115Y123_AQ;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_B6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X80Y132_SLICE_X124Y132_D2 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X124Y132_D3 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X124Y132_D4 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_C1 = CLBLL_R_X75Y113_SLICE_X114Y113_AQ;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_C2 = CLBLM_L_X76Y123_SLICE_X117Y123_AQ;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_C3 = CLBLM_L_X74Y123_SLICE_X113Y123_BQ;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_A6 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_C4 = CLBLL_R_X75Y123_SLICE_X114Y123_BQ;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_C5 = CLBLM_L_X74Y123_SLICE_X113Y123_A5Q;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_C6 = CLBLM_L_X74Y123_SLICE_X113Y123_DQ;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_D6 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X80Y132_SLICE_X124Y132_D5 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X124Y132_D6 = 1'b1;
  assign CLBLM_L_X72Y130_SLICE_X109Y130_A1 = CLBLM_L_X72Y130_SLICE_X108Y130_DQ;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_D1 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_D2 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_D3 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_D4 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_D5 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_D6 = 1'b1;
  assign CLBLM_L_X72Y130_SLICE_X109Y130_A2 = CLBLM_L_X72Y133_SLICE_X109Y133_DO6;
  assign CLBLM_L_X72Y130_SLICE_X109Y130_A3 = CLBLM_L_X72Y130_SLICE_X109Y130_AQ;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y130_SLICE_X109Y130_A4 = CLBLM_L_X72Y131_SLICE_X108Y131_A5Q;
  assign CLBLM_L_X72Y130_SLICE_X109Y130_A5 = CLBLM_L_X72Y131_SLICE_X108Y131_AQ;
  assign CLBLM_L_X72Y130_SLICE_X109Y130_A6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y130_SLICE_X109Y130_B1 = CLBLM_L_X72Y130_SLICE_X108Y130_DQ;
  assign CLBLM_L_X72Y130_SLICE_X109Y130_B2 = CLBLM_L_X72Y130_SLICE_X109Y130_BQ;
  assign CLBLM_L_X72Y130_SLICE_X109Y130_B3 = CLBLM_L_X72Y130_SLICE_X109Y130_AQ;
  assign CLBLM_L_X72Y130_SLICE_X109Y130_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y130_SLICE_X109Y130_B5 = 1'b1;
  assign CLBLM_L_X72Y130_SLICE_X109Y130_B6 = CLBLM_L_X72Y131_SLICE_X109Y131_AO5;
  assign CLBLM_L_X72Y130_SLICE_X109Y130_C1 = CLBLM_L_X72Y131_SLICE_X108Y131_AQ;
  assign CLBLM_L_X72Y130_SLICE_X109Y130_C2 = CLBLM_L_X72Y133_SLICE_X109Y133_DO6;
  assign CLBLM_L_X72Y130_SLICE_X109Y130_C3 = CLBLM_L_X72Y131_SLICE_X108Y131_A5Q;
  assign CLBLM_L_X72Y130_SLICE_X109Y130_C4 = CLBLM_L_X72Y130_SLICE_X109Y130_BQ;
  assign CLBLM_L_X72Y130_SLICE_X109Y130_C5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y130_SLICE_X109Y130_C6 = CLBLM_L_X72Y130_SLICE_X109Y130_CQ;
  assign CLBLM_L_X72Y130_SLICE_X109Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X80Y132_SLICE_X124Y132_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y130_SLICE_X109Y130_D1 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_A1 = CLBLM_L_X76Y123_SLICE_X117Y123_AQ;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_A2 = CLBLM_L_X74Y109_SLICE_X113Y109_AQ;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_A3 = CLBLM_L_X74Y123_SLICE_X113Y123_BQ;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_A4 = CLBLM_L_X74Y123_SLICE_X113Y123_A5Q;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_A6 = 1'b1;
  assign CLBLM_L_X72Y130_SLICE_X109Y130_D2 = 1'b1;
  assign CLBLM_L_X72Y130_SLICE_X109Y130_D3 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_AX = CLBLL_R_X75Y124_SLICE_X115Y124_B5Q;
  assign CLBLM_L_X72Y130_SLICE_X109Y130_D4 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_B1 = CLBLM_L_X76Y123_SLICE_X116Y123_A5Q;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_B2 = CLBLM_L_X76Y125_SLICE_X117Y125_AQ;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_B3 = CLBLL_R_X75Y124_SLICE_X114Y124_AQ;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_B4 = CLBLL_R_X75Y124_SLICE_X114Y124_BQ;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_B5 = CLBLL_R_X77Y123_SLICE_X119Y123_AQ;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_B6 = CLBLM_L_X78Y124_SLICE_X120Y124_CQ;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_A1 = CLBLM_R_X63Y105_SLICE_X95Y105_A5Q;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_A2 = CLBLM_R_X63Y105_SLICE_X94Y105_CQ;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_A3 = CLBLM_R_X63Y105_SLICE_X94Y105_C5Q;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_C1 = CLBLL_R_X77Y123_SLICE_X119Y123_AQ;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_C2 = CLBLM_L_X76Y122_SLICE_X116Y122_A5Q;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_C3 = CLBLM_L_X78Y124_SLICE_X120Y124_CQ;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_C4 = CLBLM_L_X76Y122_SLICE_X116Y122_AQ;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_C5 = CLBLM_L_X76Y123_SLICE_X116Y123_A5Q;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_C6 = CLBLM_L_X76Y122_SLICE_X116Y122_BQ;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_CE = CLBLM_L_X76Y123_SLICE_X116Y123_DO6;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_AX = CLBLM_L_X60Y101_SLICE_X90Y101_BQ;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_B1 = CLBLM_L_X64Y105_SLICE_X96Y105_BO5;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_B2 = CLBLM_L_X62Y106_SLICE_X93Y106_BQ;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_B3 = CLBLM_L_X64Y106_SLICE_X97Y106_C5Q;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_B5 = CLBLM_L_X62Y105_SLICE_X93Y105_CQ;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_D1 = CLBLL_R_X77Y123_SLICE_X119Y123_AQ;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_D2 = CLBLM_L_X78Y124_SLICE_X120Y124_CQ;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_D3 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_D4 = CLBLM_L_X76Y123_SLICE_X116Y123_A5Q;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_D5 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_D6 = 1'b1;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_C1 = CLBLM_L_X64Y106_SLICE_X96Y106_AQ;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_C2 = CLBLM_L_X62Y106_SLICE_X93Y106_CQ;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_C6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_D1 = CLBLM_L_X64Y105_SLICE_X97Y105_DO6;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_D2 = CLBLM_R_X63Y106_SLICE_X94Y106_DO6;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_D3 = CLBLM_L_X62Y107_SLICE_X93Y107_DO6;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_D4 = CLBLM_L_X62Y106_SLICE_X93Y106_AO5;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_D5 = CLBLM_R_X63Y107_SLICE_X94Y107_CO6;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_D6 = CLBLM_L_X62Y106_SLICE_X92Y106_CO6;
  assign CLBLM_L_X72Y130_SLICE_X108Y130_D1 = CLBLL_R_X71Y130_SLICE_X106Y130_BQ;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y130_SLICE_X108Y130_D2 = CLBLM_L_X72Y130_SLICE_X108Y130_CQ;
  assign CLBLM_L_X72Y130_SLICE_X108Y130_D3 = CLBLM_L_X72Y130_SLICE_X108Y130_DQ;
  assign CLBLM_L_X72Y130_SLICE_X108Y130_D4 = CLBLL_R_X71Y125_SLICE_X107Y125_BO6;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_A1 = CLBLM_R_X63Y105_SLICE_X94Y105_CQ;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_A2 = CLBLM_L_X64Y106_SLICE_X96Y106_AQ;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_A3 = CLBLM_L_X62Y106_SLICE_X92Y106_AQ;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_A4 = CLBLM_L_X62Y106_SLICE_X93Y106_AQ;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_A5 = CLBLM_R_X63Y105_SLICE_X94Y105_C5Q;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_A6 = CLBLM_L_X62Y106_SLICE_X93Y106_CQ;
  assign CLBLM_L_X72Y130_SLICE_X108Y130_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X67Y96_SLICE_X101Y96_A1 = CLBLM_R_X67Y96_SLICE_X101Y96_CQ;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_AX = CLBLM_L_X62Y106_SLICE_X93Y106_AQ;
  assign CLBLM_R_X67Y96_SLICE_X101Y96_A2 = CLBLM_R_X67Y98_SLICE_X101Y98_BO6;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_B1 = CLBLM_L_X64Y106_SLICE_X96Y106_CQ;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_B2 = CLBLM_L_X62Y107_SLICE_X93Y107_BQ;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_B3 = CLBLM_L_X62Y106_SLICE_X92Y106_AQ;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_B4 = CLBLM_R_X63Y105_SLICE_X94Y105_CQ;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_B5 = CLBLM_R_X63Y105_SLICE_X94Y105_C5Q;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_B6 = CLBLM_R_X63Y107_SLICE_X95Y107_BQ;
  assign CLBLM_R_X67Y96_SLICE_X101Y96_A3 = CLBLM_R_X67Y96_SLICE_X101Y96_AQ;
  assign CLBLM_R_X67Y96_SLICE_X101Y96_A4 = CLBLM_R_X67Y98_SLICE_X100Y98_B5Q;
  assign CLBLM_R_X67Y96_SLICE_X101Y96_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_BX = CLBLM_L_X62Y106_SLICE_X92Y106_AQ;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_C1 = CLBLM_L_X62Y106_SLICE_X92Y106_AO6;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_C2 = CLBLM_R_X63Y106_SLICE_X94Y106_CO6;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_C3 = CLBLM_R_X63Y106_SLICE_X95Y106_DO6;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_C4 = CLBLM_L_X62Y107_SLICE_X92Y107_AO6;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_C5 = CLBLM_L_X62Y106_SLICE_X92Y106_DO6;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_C6 = CLBLM_L_X62Y106_SLICE_X92Y106_BO6;
  assign CLBLM_R_X67Y96_SLICE_X101Y96_B4 = CLBLM_R_X67Y98_SLICE_X100Y98_B5Q;
  assign CLBLM_R_X67Y96_SLICE_X101Y96_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y96_SLICE_X101Y96_B6 = CLBLM_R_X67Y98_SLICE_X101Y98_CO6;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X67Y96_SLICE_X101Y96_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y96_SLICE_X101Y96_C2 = CLBLM_R_X67Y96_SLICE_X101Y96_CQ;
  assign CLBLM_R_X67Y96_SLICE_X101Y96_C3 = CLBLM_R_X67Y98_SLICE_X100Y98_CO5;
  assign CLBLM_R_X67Y96_SLICE_X101Y96_C4 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_D1 = CLBLM_R_X63Y105_SLICE_X94Y105_C5Q;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_D2 = CLBLM_L_X64Y106_SLICE_X96Y106_A5Q;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_D3 = CLBLM_R_X63Y105_SLICE_X95Y105_A5Q;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_D4 = CLBLM_L_X62Y105_SLICE_X93Y105_CQ;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_D5 = 1'b1;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_D6 = CLBLM_R_X63Y105_SLICE_X94Y105_CQ;
  assign CLBLM_R_X67Y96_SLICE_X101Y96_D1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y96_SLICE_X101Y96_D2 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X67Y96_SLICE_X101Y96_D3 = CLBLM_R_X67Y96_SLICE_X101Y96_DQ;
  assign CLBLM_R_X67Y96_SLICE_X101Y96_D4 = CLBLM_R_X67Y98_SLICE_X101Y98_CO6;
  assign CLBLM_R_X67Y96_SLICE_X101Y96_D5 = CLBLM_R_X67Y98_SLICE_X100Y98_CO5;
  assign CLBLM_R_X67Y96_SLICE_X101Y96_D6 = CLBLM_R_X67Y97_SLICE_X101Y97_DQ;
  assign CLBLM_R_X67Y96_SLICE_X100Y96_A1 = 1'b1;
  assign CLBLM_R_X67Y96_SLICE_X100Y96_A2 = 1'b1;
  assign CLBLM_R_X67Y96_SLICE_X100Y96_A3 = 1'b1;
  assign CLBLM_R_X67Y96_SLICE_X100Y96_A4 = 1'b1;
  assign CLBLM_R_X67Y96_SLICE_X100Y96_A5 = 1'b1;
  assign CLBLM_R_X67Y96_SLICE_X100Y96_A6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_D1 = CLBLL_R_X73Y103_SLICE_X111Y103_A5Q;
  assign CLBLM_R_X67Y96_SLICE_X100Y96_B1 = 1'b1;
  assign CLBLM_R_X67Y96_SLICE_X100Y96_B2 = 1'b1;
  assign CLBLM_R_X67Y96_SLICE_X100Y96_B3 = 1'b1;
  assign CLBLM_R_X67Y96_SLICE_X100Y96_B4 = 1'b1;
  assign CLBLM_R_X67Y96_SLICE_X100Y96_B5 = 1'b1;
  assign CLBLM_R_X67Y96_SLICE_X100Y96_B6 = 1'b1;
  assign CLBLM_R_X67Y96_SLICE_X100Y96_C1 = 1'b1;
  assign CLBLM_R_X67Y96_SLICE_X100Y96_C2 = 1'b1;
  assign CLBLM_R_X67Y96_SLICE_X100Y96_C3 = 1'b1;
  assign CLBLM_R_X67Y96_SLICE_X100Y96_C4 = 1'b1;
  assign CLBLM_R_X67Y96_SLICE_X100Y96_C5 = 1'b1;
  assign CLBLM_R_X67Y96_SLICE_X100Y96_C6 = 1'b1;
  assign CLBLM_R_X67Y96_SLICE_X100Y96_D1 = 1'b1;
  assign CLBLM_R_X67Y96_SLICE_X100Y96_D2 = 1'b1;
  assign CLBLM_R_X67Y96_SLICE_X100Y96_D3 = 1'b1;
  assign CLBLM_R_X67Y96_SLICE_X100Y96_D4 = 1'b1;
  assign CLBLM_R_X67Y96_SLICE_X100Y96_D5 = 1'b1;
  assign CLBLM_R_X67Y96_SLICE_X100Y96_D6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_T1 = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_T1 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_B5 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_B6 = 1'b1;
  assign LIOI3_SING_X0Y50_OLOGIC_X0Y50_D1 = CLBLM_L_X60Y97_SLICE_X90Y97_DQ;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_A2 = CLBLM_L_X76Y125_SLICE_X117Y125_AQ;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_A3 = CLBLL_R_X75Y124_SLICE_X114Y124_AQ;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_A4 = CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_A5 = CLBLL_R_X75Y124_SLICE_X114Y124_BQ;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_A6 = CLBLL_R_X75Y123_SLICE_X115Y123_DO6;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y63_D1 = CLBLL_R_X73Y102_SLICE_X111Y102_A5Q;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_B2 = CLBLL_R_X75Y124_SLICE_X114Y124_BQ;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_B3 = 1'b1;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_B4 = CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_B5 = CLBLM_L_X76Y125_SLICE_X117Y125_AQ;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_B6 = CLBLL_R_X75Y123_SLICE_X115Y123_DO6;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_C1 = CLBLL_R_X75Y124_SLICE_X114Y124_C5Q;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_C2 = CLBLL_R_X75Y124_SLICE_X114Y124_D5Q;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_C3 = CLBLL_R_X75Y124_SLICE_X114Y124_DQ;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_C4 = CLBLM_L_X76Y118_SLICE_X117Y118_CQ;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_C5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_C6 = 1'b1;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_D1 = CLBLM_L_X74Y123_SLICE_X112Y123_BQ;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_D2 = CLBLL_R_X75Y124_SLICE_X114Y124_D5Q;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_D3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_D4 = CLBLM_L_X76Y123_SLICE_X117Y123_CQ;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_D5 = CLBLL_R_X75Y121_SLICE_X114Y121_AQ;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_D6 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_A1 = CLBLM_L_X72Y131_SLICE_X108Y131_A5Q;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_A2 = 1'b1;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_A3 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_A4 = CLBLM_L_X72Y133_SLICE_X109Y133_DO6;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_A5 = CLBLM_L_X72Y131_SLICE_X108Y131_AQ;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_A6 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_B1 = CLBLM_L_X72Y134_SLICE_X109Y134_AO5;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_B2 = CLBLM_L_X72Y131_SLICE_X109Y131_BQ;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_B3 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_B5 = CLBLM_L_X72Y131_SLICE_X109Y131_DQ;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_B6 = CLBLM_L_X72Y131_SLICE_X109Y131_AO5;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_C1 = CLBLM_L_X72Y131_SLICE_X108Y131_AQ;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_C2 = CLBLM_L_X72Y131_SLICE_X109Y131_CQ;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_C3 = CLBLM_L_X72Y134_SLICE_X109Y134_BO5;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_C4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_C5 = CLBLM_L_X72Y131_SLICE_X108Y131_A5Q;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_C6 = CLBLM_L_X72Y133_SLICE_X109Y133_DO6;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y63_T1 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_A1 = CLBLL_R_X75Y124_SLICE_X115Y124_B5Q;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_A2 = CLBLM_L_X74Y123_SLICE_X113Y123_CO5;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_A3 = CLBLL_R_X75Y124_SLICE_X115Y124_AQ;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_A5 = CLBLL_R_X75Y122_SLICE_X114Y122_AQ;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_A6 = CLBLM_L_X76Y124_SLICE_X116Y124_AQ;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_D1 = CLBLM_L_X72Y131_SLICE_X108Y131_AQ;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_D2 = CLBLM_L_X72Y131_SLICE_X109Y131_CQ;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_B1 = CLBLM_L_X76Y124_SLICE_X116Y124_CO6;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_B2 = CLBLL_R_X75Y124_SLICE_X114Y124_CQ;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_B3 = CLBLL_R_X75Y124_SLICE_X115Y124_B5Q;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_B4 = CLBLL_R_X75Y123_SLICE_X115Y123_AO5;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_B6 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_D4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_A1 = CLBLM_L_X62Y107_SLICE_X93Y107_AQ;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_A2 = CLBLM_R_X63Y106_SLICE_X95Y106_BQ;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_C1 = CLBLM_L_X74Y123_SLICE_X113Y123_CO5;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_C2 = CLBLL_R_X75Y124_SLICE_X115Y124_CQ;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_C3 = CLBLM_L_X76Y124_SLICE_X116Y124_A5Q;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_C4 = 1'b1;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_C5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_C6 = CLBLL_R_X79Y127_SLICE_X122Y127_CQ;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_A3 = CLBLM_L_X64Y106_SLICE_X96Y106_BO5;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_A4 = CLBLM_L_X64Y105_SLICE_X96Y105_AO6;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_A6 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_AX = CLBLL_R_X75Y107_SLICE_X114Y107_AQ;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_B1 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_B2 = CLBLM_L_X62Y107_SLICE_X92Y107_BO6;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_D1 = CLBLM_L_X74Y123_SLICE_X113Y123_CO5;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_D2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_D3 = CLBLL_R_X75Y124_SLICE_X115Y124_DQ;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_D4 = 1'b1;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_D5 = CLBLL_R_X79Y127_SLICE_X122Y127_BQ;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_D6 = CLBLM_L_X76Y124_SLICE_X116Y124_CQ;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_B6 = CLBLM_L_X62Y107_SLICE_X93Y107_BQ;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_C1 = CLBLM_R_X63Y105_SLICE_X95Y105_A5Q;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_C2 = CLBLL_R_X75Y107_SLICE_X114Y107_AQ;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_C3 = CLBLM_L_X62Y107_SLICE_X93Y107_BQ;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_C4 = CLBLM_L_X62Y107_SLICE_X93Y107_A5Q;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_C5 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_C6 = 1'b1;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_D1 = CLBLM_L_X62Y107_SLICE_X93Y107_CO5;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_D2 = CLBLM_R_X63Y105_SLICE_X94Y105_CQ;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_D3 = CLBLM_R_X63Y105_SLICE_X94Y105_C5Q;
  assign CLBLL_R_X73Y113_SLICE_X110Y113_A1 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X110Y113_A2 = CLBLL_R_X73Y108_SLICE_X110Y108_AQ;
  assign CLBLL_R_X73Y113_SLICE_X110Y113_A3 = CLBLL_R_X73Y113_SLICE_X110Y113_AQ;
  assign CLBLL_R_X73Y113_SLICE_X110Y113_A4 = CLBLL_R_X71Y117_SLICE_X106Y117_A5Q;
  assign CLBLL_R_X73Y113_SLICE_X110Y113_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y113_SLICE_X110Y113_A6 = CLBLL_R_X73Y113_SLICE_X110Y113_A5Q;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_D4 = CLBLM_L_X62Y105_SLICE_X93Y105_DO6;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_D5 = CLBLM_L_X62Y107_SLICE_X93Y107_AQ;
  assign CLBLL_R_X73Y113_SLICE_X110Y113_AX = CLBLL_R_X71Y117_SLICE_X106Y117_A5Q;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_D6 = CLBLL_R_X75Y107_SLICE_X114Y107_AQ;
  assign CLBLL_R_X73Y113_SLICE_X110Y113_B1 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X110Y113_B2 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X110Y113_B3 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X110Y113_B4 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X110Y113_B5 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X110Y113_B6 = 1'b1;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_A1 = CLBLM_R_X63Y105_SLICE_X94Y105_C5Q;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_A2 = CLBLM_R_X63Y107_SLICE_X94Y107_AQ;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_A3 = CLBLM_L_X62Y106_SLICE_X92Y106_BQ;
  assign CLBLL_R_X73Y113_SLICE_X110Y113_C1 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X110Y113_C2 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X110Y113_C3 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X110Y113_C4 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X110Y113_C5 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X110Y113_C6 = 1'b1;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_B1 = CLBLM_L_X62Y106_SLICE_X93Y106_AQ;
  assign CLBLL_R_X73Y113_SLICE_X110Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_B2 = CLBLM_L_X60Y101_SLICE_X90Y101_BQ;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_B4 = CLBLM_L_X62Y107_SLICE_X93Y107_BQ;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_B5 = CLBLM_L_X62Y107_SLICE_X93Y107_A5Q;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_B6 = CLBLL_R_X75Y107_SLICE_X114Y107_AQ;
  assign CLBLL_R_X73Y113_SLICE_X110Y113_D1 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X110Y113_D2 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X110Y113_D3 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X110Y113_D4 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X110Y113_D5 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X110Y113_D6 = 1'b1;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_C2 = 1'b1;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_C3 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X110Y113_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_C6 = 1'b1;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_D1 = 1'b1;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_D2 = 1'b1;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_D3 = 1'b1;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_D4 = 1'b1;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_D5 = 1'b1;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_D6 = 1'b1;
  assign CLBLM_R_X67Y97_SLICE_X101Y97_D1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y97_SLICE_X101Y97_D2 = CLBLM_R_X67Y97_SLICE_X101Y97_CQ;
  assign CLBLM_R_X67Y97_SLICE_X101Y97_D3 = CLBLM_R_X67Y97_SLICE_X101Y97_DQ;
  assign CLBLM_R_X67Y97_SLICE_X101Y97_D4 = CLBLM_R_X67Y98_SLICE_X100Y98_CO6;
  assign CLBLM_R_X67Y97_SLICE_X101Y97_D5 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X67Y97_SLICE_X101Y97_D6 = CLBLM_R_X67Y98_SLICE_X101Y98_CO6;
  assign CLBLM_R_X67Y97_SLICE_X101Y97_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X67Y97_SLICE_X100Y97_A1 = CLBLM_R_X67Y98_SLICE_X101Y98_DQ;
  assign CLBLM_R_X67Y97_SLICE_X100Y97_A2 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X67Y97_SLICE_X100Y97_A3 = CLBLM_R_X67Y97_SLICE_X100Y97_AQ;
  assign CLBLM_R_X67Y97_SLICE_X100Y97_A4 = CLBLM_R_X67Y98_SLICE_X101Y98_CO5;
  assign CLBLM_R_X67Y97_SLICE_X100Y97_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y97_SLICE_X100Y97_A6 = CLBLM_R_X67Y98_SLICE_X100Y98_CO6;
  assign CLBLL_R_X73Y113_SLICE_X111Y113_A1 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X111Y113_A2 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X111Y113_A3 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X111Y113_A4 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X111Y113_A5 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X111Y113_A6 = 1'b1;
  assign CLBLM_R_X67Y97_SLICE_X100Y97_B1 = 1'b1;
  assign CLBLM_R_X67Y97_SLICE_X100Y97_B2 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X111Y113_B1 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X111Y113_B2 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X111Y113_B3 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X111Y113_B4 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X111Y113_B5 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X111Y113_B6 = 1'b1;
  assign CLBLM_R_X67Y97_SLICE_X100Y97_B4 = 1'b1;
  assign CLBLM_R_X67Y97_SLICE_X100Y97_B5 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X111Y113_C1 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X111Y113_C2 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X111Y113_C3 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X111Y113_C4 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X111Y113_C5 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X111Y113_C6 = 1'b1;
  assign CLBLM_R_X67Y97_SLICE_X100Y97_C3 = 1'b1;
  assign CLBLM_R_X67Y97_SLICE_X100Y97_C4 = 1'b1;
  assign CLBLM_R_X67Y97_SLICE_X100Y97_C5 = 1'b1;
  assign CLBLM_R_X67Y97_SLICE_X100Y97_C6 = 1'b1;
  assign CLBLM_R_X67Y97_SLICE_X100Y97_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X67Y97_SLICE_X100Y97_D1 = 1'b1;
  assign CLBLM_R_X67Y97_SLICE_X100Y97_D2 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X111Y113_D1 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X111Y113_D2 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X111Y113_D3 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X111Y113_D4 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X111Y113_D5 = 1'b1;
  assign CLBLL_R_X73Y113_SLICE_X111Y113_D6 = 1'b1;
  assign CLBLM_R_X67Y97_SLICE_X100Y97_D3 = 1'b1;
  assign CLBLM_R_X67Y97_SLICE_X100Y97_D4 = 1'b1;
  assign CLBLM_R_X67Y97_SLICE_X100Y97_D5 = 1'b1;
  assign CLBLM_R_X67Y97_SLICE_X100Y97_D6 = 1'b1;
  assign CLBLM_R_X67Y97_SLICE_X100Y97_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_D1 = CLBLL_R_X73Y134_SLICE_X110Y134_AO5;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_T1 = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_D1 = CLBLM_L_X70Y125_SLICE_X104Y125_DO6;
  assign LIOI3_X0Y61_OLOGIC_X0Y62_D1 = CLBLM_R_X65Y110_SLICE_X99Y110_B5Q;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_T1 = 1'b1;
  assign LIOI3_X0Y61_OLOGIC_X0Y62_T1 = 1'b1;
  assign RIOI3_X105Y105_OLOGIC_X1Y106_D1 = CLBLL_R_X75Y103_SLICE_X115Y103_AQ;
  assign LIOI3_X0Y61_OLOGIC_X0Y61_D1 = CLBLM_R_X65Y109_SLICE_X98Y109_A5Q;
  assign RIOI3_X105Y105_OLOGIC_X1Y106_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1 = CLBLM_L_X70Y110_SLICE_X104Y110_CQ;
  assign LIOI3_X0Y61_OLOGIC_X0Y61_T1 = 1'b1;
  assign CLBLM_L_X72Y132_SLICE_X109Y132_A1 = CLBLM_L_X74Y134_SLICE_X113Y134_CQ;
  assign CLBLM_L_X72Y132_SLICE_X109Y132_A2 = CLBLM_L_X60Y92_SLICE_X90Y92_AQ;
  assign CLBLM_L_X72Y132_SLICE_X109Y132_A3 = CLBLL_R_X73Y133_SLICE_X110Y133_A5Q;
  assign CLBLM_L_X72Y132_SLICE_X109Y132_A4 = CLBLM_L_X74Y134_SLICE_X113Y134_A5Q;
  assign CLBLM_L_X72Y132_SLICE_X109Y132_A5 = CLBLM_L_X70Y136_SLICE_X105Y136_CO6;
  assign CLBLM_L_X72Y132_SLICE_X109Y132_A6 = CLBLL_R_X73Y132_SLICE_X111Y132_BO6;
  assign LIOB33_X0Y83_IOB_X0Y83_O = CLBLM_L_X70Y99_SLICE_X104Y99_AQ;
  assign LIOB33_X0Y83_IOB_X0Y84_O = CLBLM_L_X60Y99_SLICE_X90Y99_CQ;
  assign CLBLM_L_X72Y132_SLICE_X109Y132_AX = CLBLM_L_X72Y133_SLICE_X108Y133_AQ;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1 = 1'b1;
  assign CLBLM_L_X72Y132_SLICE_X109Y132_B1 = CLBLM_L_X72Y132_SLICE_X109Y132_DO6;
  assign CLBLM_L_X72Y132_SLICE_X109Y132_B2 = CLBLM_L_X72Y132_SLICE_X109Y132_CO6;
  assign CLBLM_L_X72Y132_SLICE_X109Y132_B3 = CLBLL_R_X71Y131_SLICE_X106Y131_AQ;
  assign CLBLM_L_X72Y132_SLICE_X109Y132_B4 = CLBLM_L_X72Y132_SLICE_X108Y132_BQ;
  assign CLBLM_L_X72Y132_SLICE_X109Y132_B5 = CLBLM_L_X72Y134_SLICE_X108Y134_AQ;
  assign CLBLM_L_X72Y132_SLICE_X109Y132_B6 = CLBLL_R_X71Y131_SLICE_X107Y131_A5Q;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1 = RIOB33_X105Y55_IOB_X1Y55_I;
  assign CLBLM_L_X72Y132_SLICE_X109Y132_C1 = CLBLM_L_X72Y132_SLICE_X108Y132_CQ;
  assign CLBLM_L_X72Y132_SLICE_X109Y132_C2 = CLBLM_L_X72Y133_SLICE_X108Y133_CQ;
  assign CLBLM_L_X72Y132_SLICE_X109Y132_C3 = 1'b1;
  assign CLBLM_L_X72Y132_SLICE_X109Y132_C4 = CLBLL_R_X71Y131_SLICE_X107Y131_A5Q;
  assign CLBLM_L_X72Y132_SLICE_X109Y132_C5 = CLBLL_R_X71Y131_SLICE_X106Y131_AQ;
  assign CLBLM_L_X72Y132_SLICE_X109Y132_C6 = CLBLL_R_X71Y132_SLICE_X106Y132_AQ;
  assign CLBLM_L_X72Y132_SLICE_X109Y132_CE = CLBLM_L_X76Y109_SLICE_X116Y109_AO6;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_T1 = 1'b1;
  assign CLBLM_L_X72Y132_SLICE_X109Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_D1 = CLBLM_L_X62Y99_SLICE_X93Y99_AQ;
  assign CLBLM_L_X72Y132_SLICE_X109Y132_D1 = CLBLM_L_X72Y132_SLICE_X108Y132_AQ;
  assign CLBLM_L_X72Y132_SLICE_X109Y132_D2 = CLBLL_R_X71Y131_SLICE_X107Y131_A5Q;
  assign CLBLM_L_X72Y132_SLICE_X109Y132_D3 = 1'b1;
  assign CLBLM_L_X72Y132_SLICE_X109Y132_D4 = CLBLL_R_X71Y131_SLICE_X106Y131_AQ;
  assign CLBLM_L_X72Y132_SLICE_X109Y132_D5 = CLBLM_L_X72Y132_SLICE_X108Y132_DQ;
  assign CLBLM_L_X72Y132_SLICE_X109Y132_D6 = CLBLL_R_X71Y132_SLICE_X106Y132_AQ;
  assign RIOB33_X105Y171_IOB_X1Y171_O = 1'b1;
  assign RIOB33_X105Y171_IOB_X1Y172_O = 1'b1;
  assign CLBLM_L_X72Y132_SLICE_X109Y132_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X103Y76_SLICE_X163Y76_AX = CLBLM_R_X103Y75_SLICE_X163Y75_BQ;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_T1 = 1'b1;
  assign CLBLM_L_X72Y132_SLICE_X108Y132_A1 = CLBLL_R_X71Y132_SLICE_X107Y132_AQ;
  assign CLBLM_L_X72Y132_SLICE_X108Y132_A2 = CLBLM_L_X72Y134_SLICE_X108Y134_AQ;
  assign CLBLM_L_X72Y132_SLICE_X108Y132_A3 = CLBLM_L_X72Y132_SLICE_X108Y132_AQ;
  assign CLBLM_L_X72Y132_SLICE_X108Y132_A4 = CLBLM_L_X72Y133_SLICE_X108Y133_BO6;
  assign CLBLM_L_X72Y132_SLICE_X108Y132_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y132_SLICE_X108Y132_A6 = CLBLL_R_X73Y132_SLICE_X110Y132_AO6;
  assign CLBLM_R_X103Y76_SLICE_X163Y76_B1 = 1'b1;
  assign CLBLM_L_X72Y132_SLICE_X108Y132_B1 = CLBLL_R_X73Y132_SLICE_X110Y132_AO6;
  assign CLBLM_L_X72Y132_SLICE_X108Y132_B2 = CLBLM_L_X72Y132_SLICE_X108Y132_BQ;
  assign CLBLM_L_X72Y132_SLICE_X108Y132_B3 = CLBLM_L_X72Y132_SLICE_X108Y132_CQ;
  assign CLBLM_L_X72Y132_SLICE_X108Y132_B4 = CLBLM_L_X72Y133_SLICE_X108Y133_BO6;
  assign CLBLM_L_X72Y132_SLICE_X108Y132_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y132_SLICE_X108Y132_B6 = CLBLM_L_X72Y133_SLICE_X108Y133_A5Q;
  assign CLBLM_R_X103Y76_SLICE_X163Y76_B2 = 1'b1;
  assign CLBLM_R_X103Y76_SLICE_X163Y76_B3 = 1'b1;
  assign CLBLM_R_X103Y76_SLICE_X163Y76_B4 = 1'b1;
  assign CLBLM_L_X72Y132_SLICE_X108Y132_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y132_SLICE_X108Y132_C2 = CLBLL_R_X73Y132_SLICE_X110Y132_BO6;
  assign CLBLM_L_X72Y132_SLICE_X108Y132_C3 = CLBLM_L_X72Y132_SLICE_X108Y132_DQ;
  assign CLBLM_L_X72Y132_SLICE_X108Y132_C4 = CLBLL_R_X73Y132_SLICE_X110Y132_AO6;
  assign CLBLM_L_X72Y132_SLICE_X108Y132_C5 = CLBLL_R_X71Y132_SLICE_X107Y132_AO6;
  assign CLBLM_L_X72Y132_SLICE_X108Y132_C6 = CLBLM_L_X72Y132_SLICE_X108Y132_CQ;
  assign CLBLM_R_X103Y76_SLICE_X163Y76_B5 = 1'b1;
  assign CLBLM_L_X72Y132_SLICE_X108Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X103Y76_SLICE_X163Y76_B6 = 1'b1;
  assign CLBLM_L_X72Y132_SLICE_X108Y132_D1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y132_SLICE_X108Y132_D2 = CLBLM_L_X72Y133_SLICE_X108Y133_DO5;
  assign CLBLM_L_X72Y132_SLICE_X108Y132_D3 = CLBLM_L_X72Y132_SLICE_X108Y132_DQ;
  assign CLBLM_L_X72Y132_SLICE_X108Y132_D4 = CLBLL_R_X73Y132_SLICE_X110Y132_AO6;
  assign CLBLM_L_X72Y132_SLICE_X108Y132_D5 = CLBLL_R_X73Y132_SLICE_X110Y132_BO6;
  assign CLBLM_L_X72Y132_SLICE_X108Y132_D6 = CLBLM_L_X72Y133_SLICE_X108Y133_CQ;
  assign CLBLM_L_X72Y132_SLICE_X108Y132_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X67Y98_SLICE_X101Y98_A1 = CLBLM_R_X67Y98_SLICE_X100Y98_BQ;
  assign CLBLM_R_X67Y98_SLICE_X101Y98_A2 = 1'b1;
  assign CLBLM_R_X67Y98_SLICE_X101Y98_A3 = 1'b1;
  assign CLBLM_R_X67Y98_SLICE_X101Y98_A4 = CLBLM_R_X67Y98_SLICE_X100Y98_B5Q;
  assign CLBLM_R_X67Y98_SLICE_X101Y98_A5 = CLBLM_R_X67Y98_SLICE_X100Y98_AQ;
  assign CLBLM_R_X67Y98_SLICE_X101Y98_A6 = 1'b1;
  assign CLBLM_R_X103Y76_SLICE_X163Y76_C1 = 1'b1;
  assign CLBLM_R_X103Y76_SLICE_X163Y76_C2 = 1'b1;
  assign CLBLM_R_X67Y98_SLICE_X101Y98_B1 = CLBLM_R_X67Y98_SLICE_X100Y98_A5Q;
  assign CLBLM_R_X67Y98_SLICE_X101Y98_B2 = 1'b1;
  assign CLBLM_R_X67Y98_SLICE_X101Y98_B3 = 1'b1;
  assign CLBLM_R_X67Y98_SLICE_X101Y98_B4 = 1'b1;
  assign CLBLM_R_X67Y98_SLICE_X101Y98_B5 = CLBLM_L_X68Y101_SLICE_X102Y101_BQ;
  assign CLBLM_R_X67Y98_SLICE_X101Y98_B6 = 1'b1;
  assign CLBLM_R_X103Y76_SLICE_X163Y76_C3 = 1'b1;
  assign CLBLM_R_X103Y76_SLICE_X163Y76_C4 = 1'b1;
  assign CLBLM_R_X67Y98_SLICE_X101Y98_C1 = CLBLM_L_X68Y101_SLICE_X102Y101_BQ;
  assign CLBLM_R_X67Y98_SLICE_X101Y98_C2 = CLBLM_R_X67Y98_SLICE_X100Y98_A5Q;
  assign CLBLM_R_X67Y98_SLICE_X101Y98_C3 = 1'b1;
  assign CLBLM_R_X67Y98_SLICE_X101Y98_C4 = 1'b1;
  assign CLBLM_R_X67Y98_SLICE_X101Y98_C5 = 1'b1;
  assign CLBLM_R_X67Y98_SLICE_X101Y98_C6 = 1'b1;
  assign CLBLM_R_X103Y76_SLICE_X163Y76_C5 = 1'b1;
  assign CLBLM_R_X67Y98_SLICE_X101Y98_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X103Y76_SLICE_X163Y76_C6 = 1'b1;
  assign CLBLM_R_X67Y98_SLICE_X101Y98_D1 = CLBLM_R_X67Y98_SLICE_X101Y98_CO5;
  assign CLBLM_R_X67Y98_SLICE_X101Y98_D2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y98_SLICE_X101Y98_D3 = CLBLM_R_X67Y98_SLICE_X101Y98_DQ;
  assign CLBLM_R_X67Y98_SLICE_X101Y98_D4 = CLBLM_R_X67Y98_SLICE_X101Y98_AO5;
  assign CLBLM_R_X67Y98_SLICE_X101Y98_D5 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X67Y98_SLICE_X101Y98_D6 = CLBLM_R_X67Y97_SLICE_X101Y97_BQ;
  assign CLBLM_R_X67Y98_SLICE_X101Y98_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X103Y76_SLICE_X163Y76_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X67Y98_SLICE_X100Y98_A1 = CLBLM_R_X67Y98_SLICE_X100Y98_B5Q;
  assign CLBLM_R_X67Y98_SLICE_X100Y98_A2 = CLBLM_R_X67Y98_SLICE_X100Y98_A5Q;
  assign CLBLM_R_X67Y98_SLICE_X100Y98_A3 = CLBLM_R_X67Y98_SLICE_X100Y98_AQ;
  assign CLBLM_R_X67Y98_SLICE_X100Y98_A4 = 1'b1;
  assign CLBLM_R_X67Y98_SLICE_X100Y98_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y98_SLICE_X100Y98_A6 = 1'b1;
  assign CLBLM_R_X67Y98_SLICE_X100Y98_B1 = CLBLM_R_X67Y98_SLICE_X100Y98_B5Q;
  assign CLBLM_R_X67Y98_SLICE_X100Y98_B2 = CLBLM_R_X67Y98_SLICE_X100Y98_BQ;
  assign CLBLM_R_X67Y98_SLICE_X100Y98_B3 = CLBLM_R_X67Y98_SLICE_X100Y98_AQ;
  assign CLBLM_R_X67Y98_SLICE_X100Y98_B4 = 1'b1;
  assign CLBLM_R_X67Y98_SLICE_X100Y98_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y98_SLICE_X100Y98_B6 = 1'b1;
  assign CLBLM_R_X67Y98_SLICE_X100Y98_C1 = 1'b1;
  assign CLBLM_R_X67Y98_SLICE_X100Y98_C2 = CLBLM_R_X67Y98_SLICE_X100Y98_AQ;
  assign CLBLM_R_X67Y98_SLICE_X100Y98_C3 = CLBLM_R_X67Y98_SLICE_X100Y98_BQ;
  assign CLBLM_R_X67Y98_SLICE_X100Y98_C4 = 1'b1;
  assign CLBLM_R_X67Y98_SLICE_X100Y98_C5 = 1'b1;
  assign CLBLM_R_X67Y98_SLICE_X100Y98_C6 = 1'b1;
  assign CLBLM_R_X103Y76_SLICE_X163Y76_D1 = 1'b1;
  assign CLBLM_R_X67Y98_SLICE_X100Y98_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X103Y76_SLICE_X163Y76_D2 = 1'b1;
  assign CLBLM_R_X67Y98_SLICE_X100Y98_D1 = 1'b1;
  assign CLBLM_R_X67Y98_SLICE_X100Y98_D2 = 1'b1;
  assign CLBLM_R_X67Y98_SLICE_X100Y98_D3 = 1'b1;
  assign CLBLM_R_X67Y98_SLICE_X100Y98_D4 = 1'b1;
  assign CLBLM_R_X67Y98_SLICE_X100Y98_D5 = 1'b1;
  assign CLBLM_R_X67Y98_SLICE_X100Y98_D6 = 1'b1;
  assign CLBLM_R_X103Y76_SLICE_X163Y76_D3 = 1'b1;
  assign CLBLM_R_X103Y76_SLICE_X163Y76_D4 = 1'b1;
  assign CLBLM_R_X67Y98_SLICE_X100Y98_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X103Y76_SLICE_X163Y76_D5 = 1'b1;
  assign CLBLM_R_X103Y76_SLICE_X163Y76_D6 = 1'b1;
  assign CLBLM_R_X103Y76_SLICE_X163Y76_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X103Y76_SLICE_X162Y76_A1 = CLBLM_R_X103Y75_SLICE_X162Y75_BQ;
  assign CLBLM_R_X103Y76_SLICE_X162Y76_A2 = CLBLM_R_X103Y76_SLICE_X162Y76_BQ;
  assign CLBLM_R_X103Y76_SLICE_X162Y76_A3 = CLBLL_R_X79Y104_SLICE_X122Y104_AQ;
  assign CLBLM_R_X103Y76_SLICE_X162Y76_A4 = CLBLM_R_X103Y75_SLICE_X163Y75_AQ;
  assign CLBLM_R_X103Y76_SLICE_X162Y76_A5 = CLBLM_R_X103Y75_SLICE_X162Y75_AO6;
  assign CLBLM_R_X103Y76_SLICE_X162Y76_A6 = CLBLM_R_X103Y76_SLICE_X163Y76_AQ;
  assign CLBLM_L_X78Y130_SLICE_X120Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOB33_X0Y85_IOB_X0Y86_O = CLBLM_L_X70Y100_SLICE_X105Y100_CQ;
  assign LIOB33_X0Y85_IOB_X0Y85_O = CLBLM_L_X60Y94_SLICE_X90Y94_BQ;
  assign CLBLM_R_X103Y76_SLICE_X162Y76_AX = CLBLL_R_X79Y104_SLICE_X122Y104_AQ;
  assign CLBLM_R_X103Y76_SLICE_X162Y76_B2 = 1'b1;
  assign CLBLM_R_X103Y76_SLICE_X162Y76_B3 = 1'b1;
  assign CLBLM_L_X72Y133_SLICE_X109Y133_A1 = 1'b1;
  assign CLBLM_L_X72Y133_SLICE_X109Y133_A2 = CLBLL_R_X73Y132_SLICE_X111Y132_AO5;
  assign CLBLM_L_X72Y133_SLICE_X109Y133_A3 = CLBLL_R_X73Y131_SLICE_X110Y131_AQ;
  assign CLBLM_L_X72Y133_SLICE_X109Y133_A4 = CLBLM_L_X74Y133_SLICE_X112Y133_AQ;
  assign CLBLM_L_X72Y133_SLICE_X109Y133_A5 = CLBLM_L_X74Y132_SLICE_X112Y132_CQ;
  assign CLBLM_L_X72Y133_SLICE_X109Y133_A6 = 1'b1;
  assign CLBLM_R_X103Y76_SLICE_X162Y76_B4 = 1'b1;
  assign CLBLM_R_X103Y76_SLICE_X162Y76_B5 = 1'b1;
  assign RIOB33_X105Y173_IOB_X1Y173_O = 1'b1;
  assign CLBLM_L_X72Y133_SLICE_X109Y133_B1 = CLBLM_L_X72Y133_SLICE_X108Y133_A5Q;
  assign CLBLM_L_X72Y133_SLICE_X109Y133_B2 = CLBLM_L_X72Y133_SLICE_X109Y133_BQ;
  assign CLBLM_L_X72Y133_SLICE_X109Y133_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y133_SLICE_X109Y133_B4 = CLBLL_R_X73Y132_SLICE_X110Y132_BO6;
  assign CLBLM_L_X72Y133_SLICE_X109Y133_B5 = CLBLM_L_X72Y133_SLICE_X108Y133_AQ;
  assign CLBLM_L_X72Y133_SLICE_X109Y133_B6 = CLBLL_R_X73Y133_SLICE_X110Y133_BQ;
  assign CLBLM_R_X103Y76_SLICE_X162Y76_B6 = 1'b1;
  assign LIOB33_X0Y115_IOB_X0Y115_O = CLBLM_R_X67Y118_SLICE_X100Y118_A5Q;
  assign LIOB33_X0Y115_IOB_X0Y116_O = CLBLM_L_X76Y118_SLICE_X117Y118_CQ;
  assign CLBLM_L_X72Y133_SLICE_X109Y133_C1 = CLBLL_R_X71Y134_SLICE_X106Y134_AQ;
  assign CLBLM_L_X72Y133_SLICE_X109Y133_C2 = CLBLM_L_X70Y136_SLICE_X105Y136_CO6;
  assign CLBLM_L_X72Y133_SLICE_X109Y133_C3 = CLBLM_L_X74Y134_SLICE_X113Y134_CQ;
  assign CLBLM_L_X72Y133_SLICE_X109Y133_C4 = CLBLL_R_X73Y133_SLICE_X111Y133_BO6;
  assign CLBLM_L_X68Y121_SLICE_X103Y121_A1 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X103Y121_A2 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X103Y121_A3 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X103Y121_A4 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X103Y121_A5 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X103Y121_A6 = 1'b1;
  assign CLBLM_L_X72Y133_SLICE_X109Y133_C5 = CLBLL_R_X73Y133_SLICE_X110Y133_A5Q;
  assign CLBLM_L_X72Y133_SLICE_X109Y133_C6 = CLBLM_L_X74Y134_SLICE_X113Y134_A5Q;
  assign CLBLM_L_X68Y121_SLICE_X103Y121_B1 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X103Y121_B2 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X103Y121_B3 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X103Y121_B4 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X103Y121_B5 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X103Y121_B6 = 1'b1;
  assign CLBLM_L_X72Y133_SLICE_X109Y133_D1 = CLBLM_L_X60Y94_SLICE_X90Y94_AQ;
  assign CLBLM_L_X72Y133_SLICE_X109Y133_D2 = CLBLM_L_X70Y136_SLICE_X105Y136_CO6;
  assign CLBLM_L_X72Y133_SLICE_X109Y133_D3 = CLBLM_L_X74Y134_SLICE_X113Y134_CQ;
  assign CLBLM_L_X68Y121_SLICE_X103Y121_C1 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X103Y121_C2 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X103Y121_C3 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X103Y121_C4 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X103Y121_C5 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X103Y121_C6 = 1'b1;
  assign CLBLM_L_X72Y133_SLICE_X108Y133_A1 = CLBLM_L_X72Y133_SLICE_X108Y133_A5Q;
  assign CLBLM_L_X72Y133_SLICE_X108Y133_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y133_SLICE_X108Y133_A3 = CLBLM_L_X72Y133_SLICE_X108Y133_AQ;
  assign CLBLM_L_X72Y133_SLICE_X108Y133_A4 = CLBLL_R_X73Y132_SLICE_X110Y132_BO6;
  assign CLBLM_L_X72Y133_SLICE_X108Y133_A5 = CLBLL_R_X71Y132_SLICE_X107Y132_AQ;
  assign CLBLM_L_X72Y133_SLICE_X108Y133_A6 = 1'b1;
  assign CLBLM_R_X103Y76_SLICE_X162Y76_C3 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X103Y121_D1 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X103Y121_D2 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X103Y121_D3 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X103Y121_D4 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X103Y121_D5 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X103Y121_D6 = 1'b1;
  assign CLBLM_L_X72Y133_SLICE_X108Y133_B1 = CLBLM_L_X72Y133_SLICE_X108Y133_A5Q;
  assign CLBLM_L_X72Y133_SLICE_X108Y133_B2 = CLBLL_R_X73Y132_SLICE_X110Y132_BO6;
  assign CLBLM_L_X72Y133_SLICE_X108Y133_B3 = CLBLM_L_X72Y133_SLICE_X108Y133_AQ;
  assign CLBLM_L_X72Y133_SLICE_X108Y133_B4 = 1'b1;
  assign CLBLM_L_X72Y133_SLICE_X108Y133_B5 = 1'b1;
  assign CLBLM_L_X72Y133_SLICE_X108Y133_B6 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X102Y121_A1 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X102Y121_A2 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X102Y121_A3 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X102Y121_A4 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X102Y121_A5 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X102Y121_A6 = 1'b1;
  assign CLBLM_L_X72Y133_SLICE_X108Y133_C1 = CLBLL_R_X73Y132_SLICE_X110Y132_AO6;
  assign CLBLM_L_X72Y133_SLICE_X108Y133_C2 = CLBLM_L_X72Y133_SLICE_X108Y133_CQ;
  assign CLBLM_L_X72Y133_SLICE_X108Y133_C3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y121_SLICE_X102Y121_AX = CLBLM_L_X72Y121_SLICE_X108Y121_AQ;
  assign CLBLM_L_X72Y133_SLICE_X108Y133_C4 = CLBLL_R_X71Y132_SLICE_X107Y132_AQ;
  assign CLBLM_L_X68Y121_SLICE_X102Y121_B1 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X102Y121_B2 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X102Y121_B3 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X102Y121_B4 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X102Y121_B5 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X102Y121_B6 = 1'b1;
  assign CLBLM_L_X72Y133_SLICE_X108Y133_D1 = CLBLL_R_X71Y132_SLICE_X107Y132_AQ;
  assign CLBLM_L_X72Y133_SLICE_X108Y133_D2 = 1'b1;
  assign CLBLM_L_X72Y133_SLICE_X108Y133_D3 = CLBLL_R_X73Y132_SLICE_X110Y132_BO6;
  assign CLBLM_L_X68Y121_SLICE_X102Y121_C1 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X102Y121_C2 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X102Y121_C3 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X102Y121_C4 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X102Y121_C5 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X102Y121_C6 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X102Y121_CE = CLBLM_L_X76Y109_SLICE_X116Y109_AO6;
  assign CLBLM_L_X72Y133_SLICE_X108Y133_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X68Y121_SLICE_X102Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X67Y99_SLICE_X101Y99_A1 = 1'b1;
  assign CLBLM_R_X67Y99_SLICE_X101Y99_A2 = 1'b1;
  assign CLBLM_R_X67Y99_SLICE_X101Y99_A3 = 1'b1;
  assign CLBLM_R_X67Y99_SLICE_X101Y99_A4 = 1'b1;
  assign CLBLM_R_X67Y99_SLICE_X101Y99_A5 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X102Y121_D1 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X102Y121_D2 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X102Y121_D3 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X102Y121_D4 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X102Y121_D5 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X102Y121_D6 = 1'b1;
  assign CLBLM_R_X67Y99_SLICE_X101Y99_A6 = 1'b1;
  assign CLBLM_R_X67Y99_SLICE_X101Y99_B1 = 1'b1;
  assign CLBLM_L_X68Y121_SLICE_X102Y121_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X67Y99_SLICE_X101Y99_B2 = 1'b1;
  assign CLBLM_R_X67Y99_SLICE_X101Y99_B3 = 1'b1;
  assign CLBLM_R_X67Y99_SLICE_X101Y99_B4 = 1'b1;
  assign CLBLM_R_X67Y99_SLICE_X101Y99_B5 = 1'b1;
  assign CLBLM_R_X67Y99_SLICE_X101Y99_B6 = 1'b1;
  assign CLBLM_R_X67Y99_SLICE_X101Y99_C1 = 1'b1;
  assign CLBLM_R_X67Y99_SLICE_X101Y99_C2 = 1'b1;
  assign CLBLM_R_X67Y99_SLICE_X101Y99_C3 = 1'b1;
  assign CLBLM_R_X67Y99_SLICE_X101Y99_C4 = 1'b1;
  assign CLBLM_R_X67Y99_SLICE_X101Y99_C5 = 1'b1;
  assign CLBLM_R_X67Y99_SLICE_X101Y99_C6 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_T1 = 1'b1;
  assign CLBLM_L_X78Y130_SLICE_X120Y130_D1 = CLBLM_L_X78Y130_SLICE_X120Y130_BQ;
  assign CLBLM_R_X67Y99_SLICE_X101Y99_D1 = 1'b1;
  assign CLBLM_R_X67Y99_SLICE_X101Y99_D2 = 1'b1;
  assign CLBLM_R_X67Y99_SLICE_X101Y99_D3 = 1'b1;
  assign CLBLM_R_X67Y99_SLICE_X101Y99_D4 = 1'b1;
  assign CLBLM_R_X67Y99_SLICE_X101Y99_D5 = 1'b1;
  assign CLBLM_R_X67Y99_SLICE_X101Y99_D6 = 1'b1;
  assign CLBLM_R_X67Y99_SLICE_X100Y99_A1 = CLBLM_R_X67Y101_SLICE_X101Y101_DO6;
  assign CLBLM_R_X67Y99_SLICE_X100Y99_A2 = CLBLM_R_X67Y101_SLICE_X100Y101_DO6;
  assign CLBLM_R_X67Y99_SLICE_X100Y99_A3 = CLBLM_R_X67Y99_SLICE_X100Y99_AQ;
  assign CLBLM_R_X67Y99_SLICE_X100Y99_A4 = CLBLM_R_X67Y100_SLICE_X100Y100_CQ;
  assign CLBLM_R_X67Y99_SLICE_X100Y99_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y99_SLICE_X100Y99_A6 = CLBLM_R_X67Y99_SLICE_X100Y99_CO6;
  assign CLBLM_R_X67Y99_SLICE_X100Y99_B1 = CLBLM_R_X67Y99_SLICE_X100Y99_DO6;
  assign CLBLM_R_X67Y99_SLICE_X100Y99_B2 = CLBLM_R_X67Y99_SLICE_X100Y99_BQ;
  assign CLBLM_R_X67Y99_SLICE_X100Y99_B3 = CLBLM_R_X67Y99_SLICE_X100Y99_AQ;
  assign CLBLM_R_X67Y99_SLICE_X100Y99_B4 = 1'b1;
  assign CLBLM_R_X67Y99_SLICE_X100Y99_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y99_SLICE_X100Y99_B6 = CLBLM_R_X67Y99_SLICE_X100Y99_CO6;
  assign CLBLM_R_X67Y99_SLICE_X100Y99_C1 = CLBLM_R_X67Y100_SLICE_X100Y100_BQ;
  assign CLBLM_R_X67Y99_SLICE_X100Y99_C2 = CLBLM_R_X67Y99_SLICE_X100Y99_AQ;
  assign CLBLM_R_X67Y99_SLICE_X100Y99_C3 = CLBLM_R_X67Y99_SLICE_X100Y99_BQ;
  assign CLBLM_R_X67Y99_SLICE_X100Y99_C4 = 1'b1;
  assign CLBLM_R_X67Y99_SLICE_X100Y99_C5 = CLBLM_R_X67Y103_SLICE_X100Y103_BQ;
  assign CLBLM_R_X67Y99_SLICE_X100Y99_C6 = CLBLM_R_X67Y100_SLICE_X100Y100_CQ;
  assign CLBLM_R_X67Y99_SLICE_X100Y99_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X67Y99_SLICE_X100Y99_D1 = CLBLM_R_X67Y101_SLICE_X100Y101_DO6;
  assign CLBLM_R_X67Y99_SLICE_X100Y99_D2 = CLBLM_R_X67Y99_SLICE_X100Y99_AQ;
  assign CLBLM_R_X67Y99_SLICE_X100Y99_D3 = 1'b1;
  assign CLBLM_R_X67Y99_SLICE_X100Y99_D4 = 1'b1;
  assign CLBLM_R_X67Y99_SLICE_X100Y99_D5 = CLBLM_R_X67Y101_SLICE_X101Y101_DO6;
  assign CLBLM_R_X67Y99_SLICE_X100Y99_D6 = CLBLM_R_X67Y100_SLICE_X100Y100_CQ;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_D1 = RIOB33_X105Y57_IOB_X1Y58_I;
  assign CLBLM_R_X67Y99_SLICE_X100Y99_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign LIOI3_TBYTESRC_X0Y81_OLOGIC_X0Y81_T1 = 1'b1;
  assign LIOB33_X0Y87_IOB_X0Y88_O = CLBLM_L_X60Y94_SLICE_X90Y94_CQ;
  assign LIOB33_X0Y87_IOB_X0Y87_O = CLBLM_R_X63Y97_SLICE_X94Y97_B5Q;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_T1 = 1'b1;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_A2 = CLBLL_R_X75Y127_SLICE_X114Y127_A5Q;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_A3 = CLBLL_R_X75Y127_SLICE_X114Y127_AQ;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_A4 = CLBLL_R_X73Y127_SLICE_X110Y127_A5Q;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_A5 = CLBLL_R_X75Y128_SLICE_X115Y128_CO6;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_A6 = 1'b1;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_B2 = CLBLL_R_X75Y127_SLICE_X114Y127_BQ;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_B3 = CLBLL_R_X73Y127_SLICE_X110Y127_A5Q;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_B4 = CLBLL_R_X75Y128_SLICE_X114Y128_BO6;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_B5 = CLBLL_R_X73Y127_SLICE_X111Y127_AQ;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_B6 = CLBLL_R_X75Y127_SLICE_X114Y127_CO6;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_C1 = CLBLL_R_X75Y127_SLICE_X114Y127_A5Q;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_C2 = CLBLL_R_X73Y127_SLICE_X110Y127_A5Q;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_C3 = 1'b1;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_C4 = CLBLL_R_X75Y128_SLICE_X115Y128_CO6;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_C5 = 1'b1;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_C6 = 1'b1;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOB33_X105Y175_IOB_X1Y176_O = CLBLL_R_X73Y119_SLICE_X110Y119_AQ;
  assign RIOB33_X105Y175_IOB_X1Y175_O = 1'b1;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_D1 = CLBLL_R_X75Y127_SLICE_X114Y127_A5Q;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_D2 = CLBLL_R_X75Y127_SLICE_X114Y127_AQ;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_D3 = CLBLL_R_X75Y127_SLICE_X114Y127_DQ;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_D4 = CLBLL_R_X75Y128_SLICE_X115Y128_CO6;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_D5 = CLBLL_R_X75Y128_SLICE_X114Y128_CQ;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_D6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y134_SLICE_X109Y134_A1 = CLBLM_L_X74Y133_SLICE_X112Y133_CQ;
  assign CLBLM_L_X72Y134_SLICE_X109Y134_A2 = CLBLM_L_X74Y134_SLICE_X113Y134_AQ;
  assign CLBLM_L_X72Y134_SLICE_X109Y134_A3 = CLBLL_R_X73Y131_SLICE_X110Y131_AQ;
  assign CLBLM_L_X72Y134_SLICE_X109Y134_A4 = 1'b1;
  assign CLBLM_L_X72Y134_SLICE_X109Y134_A5 = CLBLL_R_X73Y132_SLICE_X111Y132_AO5;
  assign CLBLM_L_X72Y134_SLICE_X109Y134_A6 = 1'b1;
  assign CLBLM_L_X72Y134_SLICE_X109Y134_B1 = CLBLM_L_X74Y133_SLICE_X112Y133_CQ;
  assign CLBLM_L_X72Y134_SLICE_X109Y134_B2 = CLBLM_L_X74Y132_SLICE_X112Y132_CQ;
  assign CLBLM_L_X72Y134_SLICE_X109Y134_B3 = 1'b1;
  assign CLBLM_L_X72Y134_SLICE_X109Y134_B4 = CLBLL_R_X73Y132_SLICE_X111Y132_AO5;
  assign CLBLM_L_X72Y134_SLICE_X109Y134_B5 = CLBLM_L_X74Y134_SLICE_X113Y134_AQ;
  assign CLBLM_L_X72Y134_SLICE_X109Y134_B6 = 1'b1;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_A1 = CLBLM_L_X60Y104_SLICE_X90Y104_AQ;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_A2 = CLBLM_L_X62Y105_SLICE_X93Y105_A5Q;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_A3 = CLBLL_R_X75Y127_SLICE_X115Y127_AQ;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_A5 = CLBLL_R_X77Y130_SLICE_X118Y130_DO5;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_A6 = CLBLM_L_X76Y128_SLICE_X117Y128_CO6;
  assign CLBLM_L_X72Y134_SLICE_X109Y134_C1 = 1'b1;
  assign CLBLM_L_X72Y134_SLICE_X109Y134_C2 = 1'b1;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_B1 = CLBLL_R_X75Y128_SLICE_X115Y128_DO6;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_B2 = CLBLL_R_X75Y127_SLICE_X115Y127_BQ;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_B3 = CLBLM_L_X74Y129_SLICE_X112Y129_AQ;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_B4 = CLBLM_L_X74Y129_SLICE_X112Y129_A5Q;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_B6 = CLBLM_L_X72Y127_SLICE_X108Y127_DQ;
  assign CLBLM_L_X72Y134_SLICE_X109Y134_C4 = 1'b1;
  assign CLBLM_L_X72Y134_SLICE_X109Y134_C5 = 1'b1;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_C1 = CLBLL_R_X75Y127_SLICE_X115Y127_BQ;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_C2 = CLBLL_R_X75Y127_SLICE_X115Y127_CQ;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_C3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_C4 = CLBLM_L_X72Y127_SLICE_X108Y127_DQ;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_C5 = CLBLM_L_X74Y128_SLICE_X113Y128_BO5;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_C6 = 1'b1;
  assign CLBLM_L_X72Y134_SLICE_X109Y134_D1 = 1'b1;
  assign CLBLM_L_X72Y134_SLICE_X109Y134_D2 = 1'b1;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X72Y134_SLICE_X109Y134_D3 = 1'b1;
  assign CLBLM_L_X72Y134_SLICE_X109Y134_D4 = 1'b1;
  assign CLBLM_L_X72Y134_SLICE_X109Y134_D5 = 1'b1;
  assign CLBLM_L_X72Y134_SLICE_X108Y134_A1 = 1'b1;
  assign CLBLM_L_X72Y134_SLICE_X108Y134_A2 = CLBLM_L_X72Y133_SLICE_X109Y133_BQ;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_D1 = CLBLM_L_X74Y129_SLICE_X112Y129_AQ;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_D2 = CLBLL_R_X75Y127_SLICE_X115Y127_CQ;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_D3 = CLBLL_R_X75Y127_SLICE_X115Y127_DQ;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_D4 = CLBLM_L_X74Y129_SLICE_X112Y129_A5Q;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_D5 = CLBLL_R_X75Y128_SLICE_X115Y128_DO6;
  assign CLBLL_R_X73Y106_SLICE_X110Y106_B4 = CLBLM_L_X74Y107_SLICE_X112Y107_CQ;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_D6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y134_SLICE_X108Y134_A3 = CLBLM_L_X72Y134_SLICE_X108Y134_AQ;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y134_SLICE_X108Y134_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y134_SLICE_X108Y134_A6 = CLBLM_L_X72Y133_SLICE_X108Y133_BO5;
  assign CLBLM_L_X72Y134_SLICE_X108Y134_B1 = 1'b1;
  assign CLBLM_L_X72Y134_SLICE_X108Y134_B2 = 1'b1;
  assign CLBLM_L_X72Y134_SLICE_X108Y134_B3 = 1'b1;
  assign CLBLM_L_X72Y134_SLICE_X108Y134_B4 = 1'b1;
  assign CLBLM_L_X72Y134_SLICE_X108Y134_B5 = 1'b1;
  assign CLBLM_L_X72Y134_SLICE_X108Y134_B6 = 1'b1;
  assign CLBLM_L_X72Y134_SLICE_X108Y134_C1 = 1'b1;
  assign CLBLM_L_X72Y134_SLICE_X108Y134_C2 = 1'b1;
  assign CLBLM_L_X72Y134_SLICE_X108Y134_C3 = 1'b1;
  assign CLBLM_L_X72Y134_SLICE_X108Y134_C4 = 1'b1;
  assign CLBLM_L_X72Y134_SLICE_X108Y134_C5 = 1'b1;
  assign CLBLM_L_X72Y134_SLICE_X108Y134_C6 = 1'b1;
  assign LIOI3_X0Y65_OLOGIC_X0Y66_D1 = CLBLM_R_X65Y110_SLICE_X98Y110_A5Q;
  assign CLBLM_L_X72Y134_SLICE_X108Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_T1 = 1'b1;
  assign CLBLM_L_X72Y134_SLICE_X108Y134_D1 = 1'b1;
  assign CLBLM_L_X72Y134_SLICE_X108Y134_D2 = 1'b1;
  assign CLBLM_L_X72Y134_SLICE_X108Y134_D3 = 1'b1;
  assign CLBLM_L_X72Y134_SLICE_X108Y134_D4 = 1'b1;
  assign CLBLM_L_X72Y134_SLICE_X108Y134_D5 = 1'b1;
  assign CLBLM_L_X72Y134_SLICE_X108Y134_D6 = 1'b1;
  assign LIOI3_X0Y65_OLOGIC_X0Y66_T1 = 1'b1;
  assign RIOI3_X105Y109_OLOGIC_X1Y110_D1 = CLBLM_L_X72Y111_SLICE_X108Y111_C5Q;
  assign CLBLM_L_X72Y134_SLICE_X108Y134_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign LIOI3_X0Y65_OLOGIC_X0Y65_D1 = CLBLM_L_X72Y107_SLICE_X109Y107_BQ;
  assign CLBLM_R_X67Y100_SLICE_X101Y100_A1 = 1'b1;
  assign CLBLM_R_X67Y100_SLICE_X101Y100_A2 = 1'b1;
  assign CLBLM_R_X67Y100_SLICE_X101Y100_A3 = 1'b1;
  assign CLBLM_R_X67Y100_SLICE_X101Y100_A4 = 1'b1;
  assign CLBLM_R_X67Y100_SLICE_X101Y100_A5 = 1'b1;
  assign CLBLM_R_X67Y100_SLICE_X101Y100_A6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1 = CLBLL_R_X71Y119_SLICE_X106Y119_AQ;
  assign RIOI3_X105Y109_OLOGIC_X1Y110_T1 = 1'b1;
  assign CLBLM_R_X67Y100_SLICE_X101Y100_B1 = 1'b1;
  assign CLBLM_R_X67Y100_SLICE_X101Y100_B2 = 1'b1;
  assign CLBLM_R_X67Y100_SLICE_X101Y100_B3 = 1'b1;
  assign CLBLM_R_X67Y100_SLICE_X101Y100_B4 = 1'b1;
  assign CLBLM_R_X67Y100_SLICE_X101Y100_B5 = 1'b1;
  assign CLBLM_R_X67Y100_SLICE_X101Y100_B6 = 1'b1;
  assign LIOI3_X0Y65_OLOGIC_X0Y65_T1 = 1'b1;
  assign RIOI3_X105Y109_OLOGIC_X1Y109_D1 = CLBLL_R_X79Y104_SLICE_X122Y104_AQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1 = 1'b1;
  assign CLBLM_R_X67Y100_SLICE_X101Y100_C1 = 1'b1;
  assign CLBLM_R_X67Y100_SLICE_X101Y100_C2 = 1'b1;
  assign CLBLM_R_X67Y100_SLICE_X101Y100_C3 = 1'b1;
  assign CLBLM_R_X67Y100_SLICE_X101Y100_C4 = 1'b1;
  assign CLBLM_R_X67Y100_SLICE_X101Y100_C5 = 1'b1;
  assign CLBLM_R_X67Y100_SLICE_X101Y100_C6 = 1'b1;
  assign RIOI3_X105Y109_OLOGIC_X1Y109_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_D1 = CLBLM_L_X82Y130_SLICE_X128Y130_AQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1 = CLBLM_R_X63Y106_SLICE_X95Y106_AQ;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_T1 = 1'b1;
  assign CLBLM_R_X67Y100_SLICE_X101Y100_D1 = 1'b1;
  assign CLBLM_R_X67Y100_SLICE_X101Y100_D2 = 1'b1;
  assign CLBLM_R_X67Y100_SLICE_X101Y100_D3 = 1'b1;
  assign CLBLM_R_X67Y100_SLICE_X101Y100_D4 = 1'b1;
  assign CLBLM_R_X67Y100_SLICE_X101Y100_D5 = 1'b1;
  assign CLBLM_R_X67Y100_SLICE_X101Y100_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_D1 = CLBLL_R_X77Y125_SLICE_X118Y125_AQ;
  assign CLBLM_R_X67Y100_SLICE_X100Y100_A1 = CLBLM_R_X67Y99_SLICE_X100Y99_CO6;
  assign CLBLM_R_X67Y100_SLICE_X100Y100_A2 = CLBLM_R_X67Y100_SLICE_X100Y100_BQ;
  assign CLBLM_R_X67Y100_SLICE_X100Y100_A3 = CLBLM_R_X67Y100_SLICE_X100Y100_AQ;
  assign CLBLM_R_X67Y100_SLICE_X100Y100_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y100_SLICE_X100Y100_A5 = 1'b1;
  assign CLBLM_R_X67Y100_SLICE_X100Y100_A6 = CLBLM_R_X67Y103_SLICE_X100Y103_BQ;
  assign CLBLM_R_X67Y100_SLICE_X100Y100_AX = CLBLM_R_X63Y105_SLICE_X95Y105_AQ;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_T1 = 1'b1;
  assign CLBLM_R_X67Y100_SLICE_X100Y100_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y100_SLICE_X100Y100_B2 = CLBLM_R_X67Y100_SLICE_X100Y100_BQ;
  assign CLBLM_R_X67Y100_SLICE_X100Y100_B3 = CLBLL_R_X77Y104_SLICE_X119Y104_A5Q;
  assign CLBLM_R_X67Y100_SLICE_X100Y100_B4 = CLBLM_R_X63Y105_SLICE_X95Y105_AQ;
  assign CLBLM_R_X67Y100_SLICE_X100Y100_B5 = 1'b1;
  assign CLBLM_R_X67Y100_SLICE_X100Y100_B6 = CLBLM_R_X67Y100_SLICE_X100Y100_A5Q;
  assign CLBLM_R_X67Y100_SLICE_X100Y100_C1 = CLBLM_R_X67Y101_SLICE_X100Y101_DO6;
  assign CLBLM_R_X67Y100_SLICE_X100Y100_C2 = CLBLM_R_X67Y100_SLICE_X100Y100_CQ;
  assign CLBLM_R_X67Y100_SLICE_X100Y100_C3 = CLBLM_R_X67Y101_SLICE_X101Y101_DO6;
  assign CLBLM_R_X67Y100_SLICE_X100Y100_C4 = CLBLM_R_X67Y99_SLICE_X100Y99_CO6;
  assign CLBLM_R_X67Y100_SLICE_X100Y100_C5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y100_SLICE_X100Y100_C6 = CLBLM_R_X67Y101_SLICE_X101Y101_BQ;
  assign CLBLM_R_X67Y100_SLICE_X100Y100_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X67Y100_SLICE_X100Y100_D1 = 1'b1;
  assign CLBLM_R_X67Y100_SLICE_X100Y100_D2 = 1'b1;
  assign CLBLM_R_X67Y100_SLICE_X100Y100_D3 = 1'b1;
  assign CLBLM_R_X67Y100_SLICE_X100Y100_D4 = 1'b1;
  assign CLBLM_R_X67Y100_SLICE_X100Y100_D5 = 1'b1;
  assign CLBLM_R_X67Y100_SLICE_X100Y100_D6 = 1'b1;
  assign CLBLM_R_X67Y100_SLICE_X100Y100_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign LIOB33_X0Y89_IOB_X0Y90_O = CLBLM_R_X63Y103_SLICE_X94Y103_AQ;
  assign LIOB33_X0Y89_IOB_X0Y89_O = CLBLM_R_X63Y98_SLICE_X94Y98_BQ;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_A1 = CLBLM_L_X76Y128_SLICE_X116Y128_A5Q;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_A2 = CLBLL_R_X75Y130_SLICE_X115Y130_AQ;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_A3 = CLBLL_R_X75Y129_SLICE_X114Y129_DQ;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_A4 = CLBLM_L_X74Y129_SLICE_X113Y129_CO6;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_A5 = 1'b1;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_A6 = 1'b1;
  assign RIOB33_X105Y177_IOB_X1Y177_O = CLBLM_L_X72Y119_SLICE_X109Y119_BQ;
  assign RIOB33_X105Y177_IOB_X1Y178_O = CLBLL_R_X73Y119_SLICE_X110Y119_BQ;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_B1 = CLBLL_R_X77Y128_SLICE_X118Y128_B5Q;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_B2 = CLBLL_R_X75Y129_SLICE_X114Y129_BQ;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_B3 = CLBLM_L_X74Y129_SLICE_X113Y129_CO6;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_B4 = CLBLM_L_X76Y128_SLICE_X116Y128_A5Q;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_B5 = 1'b1;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_B6 = 1'b1;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_C1 = CLBLL_R_X75Y127_SLICE_X114Y127_A5Q;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_C2 = CLBLL_R_X75Y128_SLICE_X114Y128_CQ;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_C3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_C4 = CLBLL_R_X75Y128_SLICE_X115Y128_CO6;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_C5 = CLBLL_R_X75Y128_SLICE_X114Y128_BO5;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_C6 = CLBLL_R_X75Y127_SLICE_X114Y127_AQ;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_D1 = 1'b1;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_D2 = CLBLM_L_X74Y129_SLICE_X113Y129_CO6;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_D3 = CLBLM_L_X76Y130_SLICE_X116Y130_AQ;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_D4 = CLBLM_L_X76Y128_SLICE_X116Y128_A5Q;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_D5 = CLBLL_R_X77Y128_SLICE_X118Y128_B5Q;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_D6 = 1'b1;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_C5 = 1'b1;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_A1 = CLBLL_R_X75Y129_SLICE_X115Y129_BO6;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_A2 = CLBLL_R_X77Y128_SLICE_X118Y128_CQ;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_A3 = CLBLM_L_X76Y128_SLICE_X117Y128_B5Q;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_A4 = CLBLL_R_X77Y129_SLICE_X118Y129_CQ;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_A5 = CLBLL_R_X75Y127_SLICE_X115Y127_AQ;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_A6 = CLBLM_L_X76Y128_SLICE_X116Y128_DO6;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_BX = CLBLM_L_X74Y117_SLICE_X112Y117_AQ;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_C6 = CLBLM_R_X65Y105_SLICE_X98Y105_CQ;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_B1 = CLBLM_L_X76Y128_SLICE_X116Y128_DO6;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_B2 = CLBLL_R_X77Y128_SLICE_X118Y128_CQ;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_B3 = CLBLM_L_X76Y128_SLICE_X117Y128_B5Q;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_B4 = CLBLL_R_X77Y129_SLICE_X118Y129_CQ;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_B5 = CLBLM_L_X60Y104_SLICE_X90Y104_AQ;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_B6 = CLBLL_R_X75Y129_SLICE_X115Y129_CO6;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_C1 = CLBLL_R_X77Y129_SLICE_X118Y129_CQ;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_C2 = CLBLM_L_X62Y105_SLICE_X93Y105_A5Q;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_C3 = CLBLL_R_X75Y129_SLICE_X115Y129_DO6;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_C4 = CLBLM_L_X76Y128_SLICE_X116Y128_DO6;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_C5 = CLBLM_L_X76Y128_SLICE_X117Y128_B5Q;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_C6 = CLBLL_R_X77Y128_SLICE_X118Y128_CQ;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_D1 = CLBLL_R_X75Y130_SLICE_X114Y130_BO6;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_D2 = CLBLL_R_X77Y126_SLICE_X118Y126_AQ;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_D3 = CLBLL_R_X77Y129_SLICE_X118Y129_CQ;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_D4 = CLBLM_L_X76Y128_SLICE_X116Y128_DO6;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_D5 = CLBLM_L_X76Y128_SLICE_X117Y128_B5Q;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_D6 = CLBLL_R_X77Y128_SLICE_X118Y128_CQ;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_D2 = 1'b1;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_D3 = CLBLM_R_X65Y103_SLICE_X98Y103_DO6;
  assign CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_D4 = CLBLM_R_X65Y105_SLICE_X98Y105_AQ;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_D5 = CLBLM_R_X65Y105_SLICE_X98Y105_B5Q;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_D6 = CLBLM_R_X63Y106_SLICE_X95Y106_AQ;
  assign CLBLM_R_X67Y101_SLICE_X101Y101_A1 = CLBLM_R_X67Y99_SLICE_X100Y99_CO6;
  assign CLBLM_R_X67Y101_SLICE_X101Y101_A2 = CLBLM_R_X67Y103_SLICE_X100Y103_BQ;
  assign CLBLM_R_X67Y101_SLICE_X101Y101_A3 = CLBLM_R_X67Y100_SLICE_X100Y100_AQ;
  assign CLBLM_R_X67Y101_SLICE_X101Y101_A4 = CLBLM_R_X67Y101_SLICE_X101Y101_AQ;
  assign CLBLM_R_X67Y101_SLICE_X101Y101_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y101_SLICE_X101Y101_A6 = CLBLM_R_X67Y100_SLICE_X100Y100_BQ;
  assign CLBLM_R_X67Y101_SLICE_X101Y101_B1 = CLBLM_R_X67Y99_SLICE_X100Y99_CO6;
  assign CLBLM_R_X67Y101_SLICE_X101Y101_B2 = CLBLM_R_X67Y101_SLICE_X101Y101_BQ;
  assign CLBLM_R_X67Y101_SLICE_X101Y101_B3 = 1'b1;
  assign CLBLM_R_X67Y101_SLICE_X101Y101_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y101_SLICE_X101Y101_B5 = CLBLM_R_X67Y101_SLICE_X101Y101_CO6;
  assign CLBLM_R_X67Y101_SLICE_X101Y101_B6 = CLBLM_R_X67Y101_SLICE_X100Y101_CQ;
  assign CLBLM_R_X67Y101_SLICE_X101Y101_C1 = CLBLM_R_X67Y100_SLICE_X100Y100_AQ;
  assign CLBLM_R_X67Y101_SLICE_X101Y101_C2 = CLBLM_R_X67Y103_SLICE_X100Y103_BQ;
  assign CLBLM_R_X67Y101_SLICE_X101Y101_C3 = CLBLM_R_X67Y101_SLICE_X100Y101_AQ;
  assign CLBLM_R_X67Y101_SLICE_X101Y101_C4 = CLBLM_R_X67Y101_SLICE_X100Y101_CQ;
  assign CLBLM_R_X67Y101_SLICE_X101Y101_C5 = CLBLM_R_X67Y100_SLICE_X100Y100_BQ;
  assign CLBLM_R_X67Y101_SLICE_X101Y101_C6 = CLBLM_R_X67Y101_SLICE_X101Y101_AQ;
  assign CLBLM_R_X67Y101_SLICE_X101Y101_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X67Y101_SLICE_X101Y101_D1 = CLBLM_R_X67Y100_SLICE_X100Y100_AQ;
  assign CLBLM_R_X67Y101_SLICE_X101Y101_D2 = CLBLM_R_X67Y101_SLICE_X100Y101_AQ;
  assign CLBLM_R_X67Y101_SLICE_X101Y101_D3 = CLBLM_R_X67Y101_SLICE_X101Y101_BQ;
  assign CLBLM_R_X67Y101_SLICE_X101Y101_D4 = CLBLM_R_X67Y101_SLICE_X100Y101_CQ;
  assign CLBLM_R_X67Y101_SLICE_X101Y101_D5 = CLBLM_R_X67Y100_SLICE_X100Y100_BQ;
  assign CLBLM_R_X67Y101_SLICE_X101Y101_D6 = CLBLM_R_X67Y101_SLICE_X101Y101_AQ;
  assign CLBLM_R_X67Y101_SLICE_X101Y101_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X67Y101_SLICE_X100Y101_A1 = 1'b1;
  assign CLBLM_R_X67Y101_SLICE_X100Y101_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y101_SLICE_X100Y101_A3 = CLBLM_R_X67Y101_SLICE_X100Y101_AQ;
  assign CLBLM_R_X67Y101_SLICE_X100Y101_A4 = CLBLM_R_X67Y101_SLICE_X100Y101_BO6;
  assign CLBLM_R_X67Y101_SLICE_X100Y101_A5 = CLBLM_R_X67Y101_SLICE_X101Y101_AQ;
  assign CLBLM_R_X67Y101_SLICE_X100Y101_A6 = CLBLM_R_X67Y99_SLICE_X100Y99_CO6;
  assign CLBLM_R_X67Y101_SLICE_X100Y101_B1 = CLBLM_R_X67Y101_SLICE_X100Y101_AQ;
  assign CLBLM_R_X67Y101_SLICE_X100Y101_B2 = CLBLM_R_X67Y101_SLICE_X101Y101_AQ;
  assign CLBLM_R_X67Y101_SLICE_X100Y101_B3 = CLBLM_R_X67Y100_SLICE_X100Y100_AQ;
  assign CLBLM_R_X67Y101_SLICE_X100Y101_B4 = CLBLM_R_X67Y103_SLICE_X100Y103_BQ;
  assign CLBLM_R_X67Y101_SLICE_X100Y101_B5 = CLBLM_R_X67Y100_SLICE_X100Y100_BQ;
  assign CLBLM_R_X67Y101_SLICE_X100Y101_B6 = 1'b1;
  assign CLBLM_R_X67Y101_SLICE_X100Y101_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y101_SLICE_X100Y101_C2 = CLBLM_R_X67Y101_SLICE_X100Y101_CQ;
  assign CLBLM_R_X67Y101_SLICE_X100Y101_C3 = 1'b1;
  assign CLBLM_R_X67Y101_SLICE_X100Y101_C4 = CLBLM_R_X67Y99_SLICE_X100Y99_CO6;
  assign CLBLM_R_X67Y101_SLICE_X100Y101_C5 = CLBLM_R_X67Y101_SLICE_X100Y101_BO5;
  assign CLBLM_R_X67Y101_SLICE_X100Y101_C6 = CLBLM_R_X67Y101_SLICE_X100Y101_AQ;
  assign RIOI3_X105Y67_OLOGIC_X1Y68_D1 = CLBLM_R_X103Y67_SLICE_X163Y67_CQ;
  assign CLBLM_R_X67Y101_SLICE_X100Y101_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X67Y101_SLICE_X100Y101_D1 = CLBLM_R_X67Y100_SLICE_X100Y100_AQ;
  assign CLBLM_R_X67Y101_SLICE_X100Y101_D2 = CLBLM_R_X67Y101_SLICE_X100Y101_CQ;
  assign CLBLM_R_X67Y101_SLICE_X100Y101_D3 = CLBLM_R_X67Y103_SLICE_X100Y103_BQ;
  assign CLBLM_R_X67Y101_SLICE_X100Y101_D4 = CLBLM_R_X67Y101_SLICE_X101Y101_AQ;
  assign CLBLM_R_X67Y101_SLICE_X100Y101_D5 = CLBLM_R_X67Y101_SLICE_X100Y101_AQ;
  assign CLBLM_R_X67Y101_SLICE_X100Y101_D6 = CLBLM_R_X67Y101_SLICE_X101Y101_BQ;
  assign LIOB33_X0Y91_IOB_X0Y91_O = CLBLM_L_X60Y99_SLICE_X90Y99_DQ;
  assign LIOB33_X0Y91_IOB_X0Y92_O = CLBLM_L_X62Y95_SLICE_X92Y95_CQ;
  assign CLBLM_R_X67Y101_SLICE_X100Y101_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign RIOB33_X105Y179_IOB_X1Y180_O = CLBLM_R_X67Y118_SLICE_X101Y118_AQ;
  assign RIOB33_X105Y179_IOB_X1Y179_O = CLBLM_L_X72Y119_SLICE_X108Y119_CQ;
  assign RIOI3_X105Y67_OLOGIC_X1Y68_T1 = 1'b1;
  assign CLBLL_R_X71Y109_SLICE_X107Y109_C3 = 1'b1;
  assign CLBLL_R_X71Y109_SLICE_X107Y109_C4 = 1'b1;
  assign CLBLL_R_X75Y129_SLICE_X114Y129_A1 = CLBLL_R_X75Y130_SLICE_X114Y130_CO6;
  assign CLBLL_R_X75Y129_SLICE_X114Y129_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y129_SLICE_X114Y129_A3 = CLBLL_R_X75Y129_SLICE_X114Y129_AQ;
  assign CLBLL_R_X71Y109_SLICE_X107Y109_C5 = 1'b1;
  assign CLBLL_R_X75Y129_SLICE_X114Y129_A4 = CLBLM_L_X76Y130_SLICE_X116Y130_A5Q;
  assign CLBLL_R_X75Y129_SLICE_X114Y129_A6 = CLBLM_L_X76Y130_SLICE_X116Y130_BQ;
  assign CLBLL_R_X75Y129_SLICE_X114Y129_A5 = CLBLL_R_X75Y129_SLICE_X114Y129_CO5;
  assign CLBLL_R_X75Y129_SLICE_X114Y129_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y129_SLICE_X114Y129_B2 = CLBLL_R_X75Y129_SLICE_X114Y129_BQ;
  assign CLBLL_R_X75Y129_SLICE_X114Y129_B3 = CLBLL_R_X75Y130_SLICE_X114Y130_AQ;
  assign CLBLL_R_X75Y129_SLICE_X114Y129_B4 = CLBLM_L_X76Y130_SLICE_X116Y130_BQ;
  assign CLBLL_R_X75Y129_SLICE_X114Y129_B5 = CLBLL_R_X75Y129_SLICE_X115Y129_AQ;
  assign CLBLL_R_X75Y129_SLICE_X114Y129_B6 = CLBLL_R_X75Y129_SLICE_X114Y129_CO6;
  assign CLBLL_R_X75Y129_SLICE_X114Y129_C1 = CLBLL_R_X77Y128_SLICE_X118Y128_CQ;
  assign CLBLL_R_X75Y129_SLICE_X114Y129_C2 = 1'b1;
  assign CLBLL_R_X75Y129_SLICE_X114Y129_C3 = CLBLL_R_X77Y129_SLICE_X118Y129_CQ;
  assign CLBLL_R_X75Y129_SLICE_X114Y129_C4 = 1'b1;
  assign CLBLL_R_X75Y129_SLICE_X114Y129_C5 = CLBLM_L_X76Y127_SLICE_X116Y127_AQ;
  assign CLBLL_R_X75Y129_SLICE_X114Y129_C6 = 1'b1;
  assign CLBLL_R_X75Y129_SLICE_X114Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X75Y129_SLICE_X114Y129_D1 = CLBLL_R_X75Y129_SLICE_X114Y129_CO5;
  assign CLBLL_R_X75Y129_SLICE_X114Y129_D2 = CLBLL_R_X75Y129_SLICE_X114Y129_AQ;
  assign CLBLL_R_X75Y129_SLICE_X114Y129_D3 = CLBLL_R_X75Y129_SLICE_X114Y129_DQ;
  assign CLBLL_R_X75Y129_SLICE_X114Y129_D4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y129_SLICE_X114Y129_D5 = CLBLL_R_X75Y130_SLICE_X114Y130_AQ;
  assign CLBLL_R_X75Y129_SLICE_X114Y129_D6 = CLBLM_L_X76Y130_SLICE_X116Y130_BQ;
  assign CLBLL_R_X75Y129_SLICE_X114Y129_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X75Y129_SLICE_X115Y129_A1 = CLBLL_R_X75Y129_SLICE_X114Y129_CO6;
  assign CLBLL_R_X75Y129_SLICE_X115Y129_A2 = CLBLL_R_X75Y130_SLICE_X115Y130_AQ;
  assign CLBLL_R_X75Y129_SLICE_X115Y129_A3 = CLBLL_R_X75Y129_SLICE_X115Y129_AQ;
  assign CLBLL_R_X75Y129_SLICE_X115Y129_A4 = CLBLM_L_X76Y129_SLICE_X116Y129_AO6;
  assign CLBLL_R_X75Y129_SLICE_X115Y129_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y129_SLICE_X115Y129_A6 = CLBLM_L_X76Y130_SLICE_X116Y130_CO6;
  assign CLBLL_R_X75Y129_SLICE_X115Y129_B1 = CLBLL_R_X77Y130_SLICE_X118Y130_AQ;
  assign CLBLL_R_X75Y129_SLICE_X115Y129_B2 = CLBLM_L_X76Y130_SLICE_X116Y130_DQ;
  assign CLBLL_R_X75Y129_SLICE_X115Y129_B3 = CLBLM_L_X76Y125_SLICE_X117Y125_BQ;
  assign CLBLL_R_X75Y129_SLICE_X115Y129_B4 = CLBLL_R_X75Y129_SLICE_X114Y129_DQ;
  assign CLBLL_R_X75Y129_SLICE_X115Y129_B5 = CLBLM_L_X78Y131_SLICE_X120Y131_AQ;
  assign CLBLL_R_X75Y129_SLICE_X115Y129_B6 = CLBLL_R_X77Y129_SLICE_X119Y129_BQ;
  assign CLBLL_R_X75Y129_SLICE_X115Y129_C1 = CLBLL_R_X75Y130_SLICE_X115Y130_AQ;
  assign CLBLL_R_X75Y129_SLICE_X115Y129_C2 = CLBLL_R_X77Y129_SLICE_X119Y129_BQ;
  assign CLBLL_R_X75Y129_SLICE_X115Y129_C3 = CLBLM_L_X76Y130_SLICE_X116Y130_DQ;
  assign CLBLL_R_X75Y129_SLICE_X115Y129_C4 = CLBLM_L_X78Y131_SLICE_X120Y131_AQ;
  assign CLBLL_R_X75Y129_SLICE_X115Y129_C5 = CLBLL_R_X77Y130_SLICE_X118Y130_AQ;
  assign CLBLL_R_X75Y129_SLICE_X115Y129_C6 = CLBLM_L_X76Y125_SLICE_X117Y125_BQ;
  assign CLBLL_R_X75Y129_SLICE_X115Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X75Y129_SLICE_X115Y129_D1 = CLBLM_L_X78Y131_SLICE_X120Y131_AQ;
  assign CLBLL_R_X75Y129_SLICE_X115Y129_D2 = CLBLM_L_X76Y125_SLICE_X117Y125_BQ;
  assign CLBLL_R_X75Y129_SLICE_X115Y129_D3 = CLBLM_L_X76Y130_SLICE_X116Y130_DQ;
  assign CLBLL_R_X75Y129_SLICE_X115Y129_D4 = CLBLL_R_X77Y129_SLICE_X119Y129_BQ;
  assign CLBLL_R_X75Y129_SLICE_X115Y129_D5 = CLBLL_R_X77Y130_SLICE_X118Y130_AQ;
  assign CLBLL_R_X75Y129_SLICE_X115Y129_D6 = CLBLL_R_X75Y129_SLICE_X114Y129_BQ;
  assign CLBLL_R_X75Y129_SLICE_X115Y129_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_D1 = CLBLL_L_X2Y131_SLICE_X0Y131_AO6;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_A1 = CLBLL_R_X73Y118_SLICE_X111Y118_A5Q;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_A2 = CLBLL_R_X73Y118_SLICE_X110Y118_BQ;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_A3 = CLBLL_R_X73Y119_SLICE_X110Y119_CO6;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_A5 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_A6 = CLBLL_R_X73Y119_SLICE_X110Y119_A5Q;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_B1 = CLBLL_R_X73Y118_SLICE_X111Y118_A5Q;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_B2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_B3 = CLBLL_R_X73Y118_SLICE_X110Y118_AQ;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_B4 = CLBLL_R_X73Y119_SLICE_X111Y119_AQ;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_B5 = CLBLL_R_X73Y119_SLICE_X110Y119_CO6;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_B6 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_C1 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_C2 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_C3 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_C4 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_C5 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_C6 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_D1 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_D2 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_D3 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_D4 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_D5 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_D6 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_T1 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_A1 = CLBLL_R_X73Y119_SLICE_X110Y119_B5Q;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_A2 = CLBLL_R_X73Y118_SLICE_X111Y118_BQ;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_A3 = CLBLL_R_X73Y119_SLICE_X110Y119_CO6;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_A5 = CLBLL_R_X73Y118_SLICE_X111Y118_A5Q;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_A6 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_B1 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_B2 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_B3 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_B4 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_B5 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_B6 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_BX = CLBLL_R_X73Y118_SLICE_X110Y118_B5Q;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_C1 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_C2 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_C3 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_C4 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_C5 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_C6 = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_D1 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOB33_X0Y93_IOB_X0Y93_O = CLBLM_L_X62Y95_SLICE_X92Y95_BQ;
  assign LIOB33_X0Y93_IOB_X0Y94_O = CLBLM_L_X62Y106_SLICE_X92Y106_AQ;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_D1 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_D2 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_D3 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_D4 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_D5 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_D6 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_D1 = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_T1 = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_D1 = 1'b1;
  assign LIOI3_X0Y67_OLOGIC_X0Y68_D1 = CLBLL_R_X71Y134_SLICE_X106Y134_AQ;
  assign LIOI3_SING_X0Y99_OLOGIC_X0Y99_D1 = RIOB33_X105Y61_IOB_X1Y62_I;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_T1 = 1'b1;
  assign RIOB33_X105Y181_IOB_X1Y182_O = CLBLL_R_X77Y128_SLICE_X119Y128_BQ;
  assign RIOB33_X105Y181_IOB_X1Y181_O = CLBLL_R_X75Y133_SLICE_X114Y133_BQ;
  assign LIOI3_X0Y67_OLOGIC_X0Y68_T1 = 1'b1;
  assign RIOI3_X105Y111_OLOGIC_X1Y112_D1 = CLBLL_R_X71Y100_SLICE_X106Y100_BQ;
  assign LIOI3_X0Y67_OLOGIC_X0Y67_D1 = CLBLM_L_X72Y103_SLICE_X109Y103_AQ;
  assign RIOI3_X105Y111_OLOGIC_X1Y112_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1 = CLBLM_L_X70Y134_SLICE_X104Y134_CO5;
  assign LIOI3_X0Y67_OLOGIC_X0Y67_T1 = 1'b1;
  assign RIOI3_X105Y111_OLOGIC_X1Y111_D1 = CLBLM_L_X62Y107_SLICE_X93Y107_BQ;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1 = CLBLL_R_X77Y124_SLICE_X118Y124_AO6;
  assign RIOI3_X105Y111_OLOGIC_X1Y111_T1 = 1'b1;
  assign CLBLL_R_X75Y130_SLICE_X114Y130_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y130_SLICE_X114Y130_A2 = CLBLL_R_X77Y129_SLICE_X118Y129_CQ;
  assign CLBLL_R_X75Y130_SLICE_X114Y130_A3 = CLBLL_R_X75Y130_SLICE_X114Y130_AQ;
  assign CLBLL_R_X75Y130_SLICE_X114Y130_A4 = CLBLM_L_X76Y130_SLICE_X116Y130_A5Q;
  assign CLBLL_R_X75Y130_SLICE_X114Y130_A5 = CLBLL_R_X77Y128_SLICE_X118Y128_CQ;
  assign CLBLL_R_X75Y130_SLICE_X114Y130_A6 = CLBLM_L_X76Y127_SLICE_X116Y127_AQ;
  assign LIOI3_SING_X0Y99_OLOGIC_X0Y99_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1 = CLBLM_L_X62Y107_SLICE_X92Y107_AO5;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1 = 1'b1;
  assign CLBLL_R_X75Y130_SLICE_X114Y130_B1 = CLBLM_L_X78Y131_SLICE_X120Y131_AQ;
  assign CLBLL_R_X75Y130_SLICE_X114Y130_B2 = CLBLM_L_X76Y130_SLICE_X116Y130_AQ;
  assign CLBLL_R_X75Y130_SLICE_X114Y130_B3 = CLBLM_L_X76Y130_SLICE_X116Y130_DQ;
  assign CLBLL_R_X75Y130_SLICE_X114Y130_B4 = CLBLM_L_X76Y125_SLICE_X117Y125_BQ;
  assign CLBLL_R_X75Y130_SLICE_X114Y130_B5 = CLBLL_R_X77Y130_SLICE_X118Y130_AQ;
  assign CLBLL_R_X75Y130_SLICE_X114Y130_B6 = CLBLL_R_X77Y129_SLICE_X119Y129_BQ;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1 = 1'b0;
  assign CLBLL_R_X75Y130_SLICE_X114Y130_C1 = CLBLM_L_X76Y128_SLICE_X117Y128_AQ;
  assign CLBLL_R_X75Y130_SLICE_X114Y130_C2 = 1'b1;
  assign CLBLL_R_X75Y130_SLICE_X114Y130_C3 = CLBLL_R_X75Y129_SLICE_X114Y129_DQ;
  assign CLBLL_R_X75Y130_SLICE_X114Y130_C4 = CLBLL_R_X77Y129_SLICE_X119Y129_BQ;
  assign CLBLL_R_X75Y130_SLICE_X114Y130_C5 = CLBLM_L_X78Y131_SLICE_X120Y131_AQ;
  assign CLBLL_R_X75Y130_SLICE_X114Y130_C6 = CLBLL_R_X77Y130_SLICE_X118Y130_AQ;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1 = 1'b1;
  assign CLBLL_R_X75Y130_SLICE_X114Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X75Y130_SLICE_X114Y130_D1 = CLBLM_L_X76Y128_SLICE_X117Y128_AQ;
  assign CLBLL_R_X75Y130_SLICE_X114Y130_D2 = CLBLL_R_X75Y130_SLICE_X115Y130_AQ;
  assign CLBLL_R_X75Y130_SLICE_X114Y130_D3 = 1'b1;
  assign CLBLL_R_X75Y130_SLICE_X114Y130_D4 = CLBLL_R_X77Y129_SLICE_X119Y129_BQ;
  assign CLBLL_R_X75Y130_SLICE_X114Y130_D5 = CLBLM_L_X78Y131_SLICE_X120Y131_AQ;
  assign CLBLL_R_X75Y130_SLICE_X114Y130_D6 = CLBLL_R_X77Y130_SLICE_X118Y130_AQ;
  assign CLBLM_R_X63Y122_SLICE_X95Y122_B4 = 1'b1;
  assign CLBLL_R_X75Y130_SLICE_X114Y130_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X75Y130_SLICE_X115Y130_A1 = CLBLL_R_X75Y130_SLICE_X115Y130_CQ;
  assign CLBLL_R_X75Y130_SLICE_X115Y130_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y130_SLICE_X115Y130_A3 = CLBLL_R_X75Y130_SLICE_X115Y130_AQ;
  assign CLBLL_R_X75Y130_SLICE_X115Y130_A4 = CLBLL_R_X75Y130_SLICE_X115Y130_BO6;
  assign CLBLL_R_X75Y130_SLICE_X115Y130_A5 = CLBLL_R_X75Y130_SLICE_X114Y130_AQ;
  assign CLBLL_R_X75Y130_SLICE_X115Y130_A6 = CLBLM_L_X76Y130_SLICE_X116Y130_BQ;
  assign CLBLL_R_X75Y130_SLICE_X115Y130_B1 = 1'b1;
  assign CLBLL_R_X75Y130_SLICE_X115Y130_B2 = CLBLL_R_X77Y128_SLICE_X118Y128_CQ;
  assign CLBLL_R_X75Y130_SLICE_X115Y130_B3 = CLBLM_L_X76Y127_SLICE_X116Y127_AQ;
  assign CLBLL_R_X75Y130_SLICE_X115Y130_B4 = 1'b1;
  assign CLBLL_R_X75Y130_SLICE_X115Y130_B5 = CLBLL_R_X77Y129_SLICE_X118Y129_CQ;
  assign CLBLL_R_X75Y130_SLICE_X115Y130_B6 = 1'b1;
  assign CLBLL_R_X75Y130_SLICE_X115Y130_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y130_SLICE_X115Y130_C2 = CLBLL_R_X75Y130_SLICE_X115Y130_CQ;
  assign CLBLL_R_X75Y130_SLICE_X115Y130_C3 = CLBLL_R_X75Y130_SLICE_X114Y130_DO6;
  assign CLBLL_R_X75Y130_SLICE_X115Y130_C4 = CLBLM_L_X76Y130_SLICE_X116Y130_CO6;
  assign CLBLL_R_X75Y130_SLICE_X115Y130_C5 = CLBLL_R_X75Y129_SLICE_X114Y129_DQ;
  assign CLBLL_R_X75Y130_SLICE_X115Y130_C6 = CLBLL_R_X75Y130_SLICE_X115Y130_BO6;
  assign CLBLL_R_X75Y130_SLICE_X115Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X75Y130_SLICE_X115Y130_D1 = 1'b1;
  assign CLBLL_R_X75Y130_SLICE_X115Y130_D2 = 1'b1;
  assign CLBLL_R_X75Y130_SLICE_X115Y130_D3 = 1'b1;
  assign CLBLL_R_X75Y130_SLICE_X115Y130_D4 = 1'b1;
  assign CLBLL_R_X75Y130_SLICE_X115Y130_D5 = 1'b1;
  assign CLBLL_R_X75Y130_SLICE_X115Y130_D6 = 1'b1;
  assign CLBLL_R_X75Y130_SLICE_X115Y130_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_A2 = CLBLL_R_X73Y119_SLICE_X110Y119_A5Q;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_A3 = CLBLL_R_X73Y118_SLICE_X111Y118_A5Q;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_A4 = CLBLM_L_X72Y119_SLICE_X109Y119_AQ;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_A5 = CLBLL_R_X73Y119_SLICE_X110Y119_CO6;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_A6 = CLBLM_L_X72Y113_SLICE_X108Y113_AQ;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_AX = CLBLL_R_X73Y119_SLICE_X110Y119_BQ;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_B1 = CLBLM_L_X72Y113_SLICE_X108Y113_AQ;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_B2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_B3 = CLBLL_R_X73Y118_SLICE_X111Y118_A5Q;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_B4 = CLBLM_L_X72Y119_SLICE_X109Y119_AQ;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_B5 = CLBLL_R_X73Y119_SLICE_X110Y119_CO6;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_B6 = 1'b1;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_C1 = CLBLL_R_X73Y119_SLICE_X111Y119_AQ;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_C2 = CLBLL_R_X73Y119_SLICE_X110Y119_AQ;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_C3 = CLBLL_R_X73Y119_SLICE_X110Y119_BQ;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_C4 = CLBLL_R_X73Y119_SLICE_X110Y119_A5Q;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_C5 = 1'b1;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_C6 = CLBLM_L_X72Y113_SLICE_X108Y113_AQ;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_D1 = 1'b1;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_D2 = 1'b1;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_D3 = 1'b1;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_D4 = 1'b1;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_D5 = 1'b1;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_D6 = 1'b1;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X67Y103_SLICE_X101Y103_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y103_SLICE_X101Y103_A2 = CLBLM_L_X68Y102_SLICE_X102Y102_CQ;
  assign CLBLM_R_X67Y103_SLICE_X101Y103_A3 = CLBLM_R_X67Y103_SLICE_X101Y103_AQ;
  assign CLBLM_R_X67Y103_SLICE_X101Y103_A4 = CLBLM_L_X68Y101_SLICE_X102Y101_BQ;
  assign CLBLM_R_X67Y103_SLICE_X101Y103_A5 = CLBLM_R_X67Y98_SLICE_X100Y98_B5Q;
  assign CLBLM_R_X67Y103_SLICE_X101Y103_A6 = CLBLM_R_X67Y98_SLICE_X100Y98_A5Q;
  assign CLBLM_R_X67Y103_SLICE_X101Y103_B1 = 1'b1;
  assign CLBLM_R_X67Y103_SLICE_X101Y103_B2 = 1'b1;
  assign CLBLM_R_X67Y103_SLICE_X101Y103_B3 = 1'b1;
  assign CLBLM_R_X67Y103_SLICE_X101Y103_B4 = 1'b1;
  assign CLBLM_R_X67Y103_SLICE_X101Y103_B5 = 1'b1;
  assign CLBLM_R_X67Y103_SLICE_X101Y103_B6 = 1'b1;
  assign CLBLM_R_X67Y103_SLICE_X101Y103_C1 = 1'b1;
  assign CLBLM_R_X67Y103_SLICE_X101Y103_C2 = 1'b1;
  assign CLBLM_R_X67Y103_SLICE_X101Y103_C3 = 1'b1;
  assign CLBLM_R_X67Y103_SLICE_X101Y103_C4 = 1'b1;
  assign CLBLM_R_X67Y103_SLICE_X101Y103_C5 = 1'b1;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_A1 = 1'b1;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_A2 = 1'b1;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_A3 = 1'b1;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_A4 = 1'b1;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_A5 = 1'b1;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_A6 = 1'b1;
  assign CLBLM_R_X67Y103_SLICE_X101Y103_C6 = 1'b1;
  assign CLBLM_R_X67Y103_SLICE_X101Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_AX = CLBLL_R_X73Y119_SLICE_X110Y119_AQ;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_B1 = 1'b1;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_B2 = 1'b1;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_B3 = 1'b1;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_B4 = 1'b1;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_B5 = 1'b1;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_B6 = 1'b1;
  assign CLBLM_R_X67Y103_SLICE_X101Y103_D1 = 1'b1;
  assign CLBLM_R_X67Y103_SLICE_X101Y103_D2 = 1'b1;
  assign CLBLM_R_X67Y103_SLICE_X101Y103_D3 = 1'b1;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_C1 = 1'b1;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_C2 = 1'b1;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_C3 = 1'b1;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_C4 = 1'b1;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_C5 = 1'b1;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_C6 = 1'b1;
  assign CLBLM_R_X67Y103_SLICE_X100Y103_A1 = CLBLM_R_X67Y103_SLICE_X100Y103_B5Q;
  assign CLBLM_R_X67Y103_SLICE_X100Y103_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X67Y103_SLICE_X100Y103_A3 = CLBLM_L_X68Y103_SLICE_X102Y103_B5Q;
  assign CLBLM_R_X67Y103_SLICE_X100Y103_A4 = CLBLM_L_X68Y99_SLICE_X102Y99_AO5;
  assign CLBLM_R_X67Y103_SLICE_X100Y103_A5 = CLBLM_L_X68Y103_SLICE_X102Y103_DQ;
  assign CLBLM_R_X67Y103_SLICE_X100Y103_A6 = 1'b1;
  assign CLBLM_R_X67Y103_SLICE_X100Y103_AX = CLBLL_R_X77Y104_SLICE_X119Y104_A5Q;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_D1 = 1'b1;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_D2 = 1'b1;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_D3 = 1'b1;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_D4 = 1'b1;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_D5 = 1'b1;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_D6 = 1'b1;
  assign CLBLM_R_X67Y103_SLICE_X100Y103_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y103_SLICE_X100Y103_B2 = CLBLM_R_X67Y103_SLICE_X100Y103_BQ;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X67Y103_SLICE_X100Y103_B3 = CLBLM_R_X67Y103_SLICE_X100Y103_AQ;
  assign CLBLM_R_X67Y103_SLICE_X100Y103_B4 = CLBLL_R_X77Y104_SLICE_X119Y104_A5Q;
  assign CLBLM_R_X67Y103_SLICE_X100Y103_B5 = CLBLM_R_X63Y105_SLICE_X95Y105_AQ;
  assign CLBLM_R_X67Y103_SLICE_X100Y103_B6 = 1'b1;
  assign CLBLM_R_X67Y103_SLICE_X100Y103_BX = CLBLM_R_X67Y103_SLICE_X100Y103_AO5;
  assign CLBLM_R_X67Y103_SLICE_X100Y103_C6 = 1'b1;
  assign CLBLM_R_X67Y103_SLICE_X100Y103_C1 = 1'b1;
  assign CLBLM_R_X67Y103_SLICE_X100Y103_C2 = 1'b1;
  assign CLBLM_R_X67Y103_SLICE_X100Y103_C3 = 1'b1;
  assign CLBLM_R_X67Y103_SLICE_X100Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X67Y103_SLICE_X100Y103_C4 = 1'b1;
  assign CLBLM_R_X67Y103_SLICE_X100Y103_C5 = 1'b1;
  assign CLBLM_R_X67Y103_SLICE_X100Y103_D1 = 1'b1;
  assign CLBLM_R_X67Y103_SLICE_X100Y103_D2 = 1'b1;
  assign CLBLM_R_X67Y103_SLICE_X100Y103_D3 = 1'b1;
  assign CLBLM_R_X67Y103_SLICE_X100Y103_D4 = 1'b1;
  assign CLBLM_R_X67Y103_SLICE_X100Y103_D5 = 1'b1;
  assign CLBLM_R_X67Y103_SLICE_X100Y103_D6 = 1'b1;
  assign CLBLM_R_X67Y103_SLICE_X100Y103_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign LIOB33_X0Y165_IOB_X0Y166_O = CLBLL_L_X2Y131_SLICE_X0Y131_AO6;
  assign LIOB33_X0Y165_IOB_X0Y165_O = CLBLL_L_X34Y123_SLICE_X50Y123_AO6;
  assign RIOB33_X105Y145_IOB_X1Y146_O = CLBLM_R_X63Y97_SLICE_X94Y97_AQ;
  assign RIOB33_X105Y145_IOB_X1Y145_O = CLBLL_R_X75Y107_SLICE_X114Y107_AQ;
  assign LIOB33_X0Y97_IOB_X0Y98_O = CLBLM_L_X68Y97_SLICE_X103Y97_AQ;
  assign LIOB33_X0Y97_IOB_X0Y97_O = CLBLM_L_X62Y103_SLICE_X92Y103_A5Q;
  assign RIOB33_X105Y185_IOB_X1Y186_O = 1'b0;
  assign RIOB33_X105Y185_IOB_X1Y185_O = CLBLL_R_X71Y117_SLICE_X106Y117_A5Q;
  assign CLBLM_L_X74Y131_SLICE_X113Y131_A1 = 1'b1;
  assign CLBLM_L_X74Y131_SLICE_X113Y131_A5 = 1'b1;
  assign CLBLM_L_X74Y131_SLICE_X113Y131_A6 = 1'b1;
  assign CLBLM_L_X74Y131_SLICE_X113Y131_B6 = 1'b1;
  assign CLBLM_L_X70Y100_SLICE_X104Y100_C5 = CLBLM_L_X70Y103_SLICE_X105Y103_CO6;
  assign CLBLM_L_X74Y131_SLICE_X113Y131_C1 = 1'b1;
  assign CLBLM_L_X74Y131_SLICE_X113Y131_C2 = 1'b1;
  assign CLBLM_L_X74Y131_SLICE_X113Y131_C3 = 1'b1;
  assign CLBLM_L_X74Y131_SLICE_X113Y131_C4 = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_D1 = 1'b1;
  assign CLBLM_L_X74Y131_SLICE_X113Y131_C5 = 1'b1;
  assign RIOI3_X105Y91_OLOGIC_X1Y91_D1 = CLBLM_L_X68Y98_SLICE_X103Y98_AQ;
  assign CLBLM_L_X74Y131_SLICE_X113Y131_C6 = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_T1 = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_T1 = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_D1 = 1'b1;
  assign LIOI3_X0Y71_OLOGIC_X0Y72_D1 = CLBLM_L_X60Y104_SLICE_X90Y104_AQ;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_T1 = 1'b1;
  assign LIOI3_X0Y71_OLOGIC_X0Y72_T1 = 1'b1;
  assign RIOI3_X105Y115_OLOGIC_X1Y116_D1 = CLBLM_L_X68Y95_SLICE_X102Y95_AQ;
  assign LIOI3_X0Y71_OLOGIC_X0Y71_D1 = CLBLM_L_X60Y94_SLICE_X90Y94_AQ;
  assign CLBLM_L_X74Y131_SLICE_X113Y131_D1 = 1'b1;
  assign RIOI3_X105Y115_OLOGIC_X1Y116_T1 = 1'b1;
  assign CLBLM_L_X74Y131_SLICE_X113Y131_D2 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1 = CLBLM_L_X64Y106_SLICE_X97Y106_AO6;
  assign RIOI3_X105Y91_OLOGIC_X1Y91_T1 = 1'b1;
  assign CLBLM_L_X74Y131_SLICE_X113Y131_D3 = 1'b1;
  assign CLBLM_L_X70Y100_SLICE_X104Y100_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign LIOI3_X0Y71_OLOGIC_X0Y71_T1 = 1'b1;
  assign RIOI3_X105Y115_OLOGIC_X1Y115_D1 = CLBLM_L_X62Y100_SLICE_X92Y100_AQ;
  assign CLBLM_L_X74Y131_SLICE_X113Y131_D4 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1 = 1'b1;
  assign CLBLM_L_X74Y131_SLICE_X113Y131_D5 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1 = CLBLL_R_X71Y117_SLICE_X106Y117_B5Q;
  assign CLBLM_L_X74Y131_SLICE_X113Y131_D6 = 1'b1;
  assign RIOI3_X105Y115_OLOGIC_X1Y115_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1 = 1'b1;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_A2 = CLBLL_R_X73Y122_SLICE_X110Y122_BQ;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_A3 = CLBLL_R_X73Y121_SLICE_X110Y121_AQ;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_A4 = CLBLL_R_X75Y128_SLICE_X114Y128_AO5;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_A5 = CLBLL_R_X73Y122_SLICE_X111Y122_AQ;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_A6 = CLBLL_R_X73Y122_SLICE_X110Y122_AO6;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1 = 1'b1;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_B1 = CLBLL_R_X75Y128_SLICE_X114Y128_AO5;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_B2 = CLBLL_R_X73Y121_SLICE_X110Y121_BQ;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_B3 = CLBLL_R_X75Y128_SLICE_X115Y128_BO6;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_B4 = CLBLL_R_X73Y122_SLICE_X110Y122_DO5;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_B6 = CLBLL_R_X73Y122_SLICE_X110Y122_CQ;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1 = CLBLL_R_X73Y108_SLICE_X110Y108_AQ;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_C1 = CLBLL_R_X73Y121_SLICE_X111Y121_AQ;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_C2 = CLBLL_R_X73Y121_SLICE_X111Y121_CO6;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_C3 = CLBLM_L_X72Y122_SLICE_X109Y122_AQ;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_C4 = CLBLM_L_X72Y122_SLICE_X109Y122_A5Q;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_C5 = CLBLL_R_X73Y121_SLICE_X110Y121_DO6;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_C6 = CLBLL_R_X73Y122_SLICE_X110Y122_BQ;
  assign LIOB33_X0Y101_IOB_X0Y101_O = RIOB33_X105Y57_IOB_X1Y58_I;
  assign LIOB33_X0Y101_IOB_X0Y102_O = RIOB33_X105Y59_IOB_X1Y59_I;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1 = 1'b1;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_D1 = CLBLL_R_X73Y123_SLICE_X111Y123_AQ;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_D2 = CLBLL_R_X73Y121_SLICE_X110Y121_AQ;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_D3 = CLBLM_L_X72Y122_SLICE_X109Y122_AQ;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_D4 = CLBLM_L_X72Y122_SLICE_X109Y122_A5Q;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_D5 = CLBLL_R_X73Y121_SLICE_X110Y121_BQ;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_D6 = 1'b1;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y131_SLICE_X112Y131_A4 = 1'b1;
  assign RIOB33_X105Y167_IOB_X1Y168_O = 1'b1;
  assign CLBLM_L_X74Y131_SLICE_X112Y131_A5 = 1'b1;
  assign CLBLM_R_X67Y105_SLICE_X101Y105_A1 = CLBLM_L_X68Y105_SLICE_X102Y105_AO5;
  assign CLBLM_R_X67Y105_SLICE_X101Y105_A2 = CLBLM_R_X67Y105_SLICE_X100Y105_BO6;
  assign CLBLM_R_X67Y105_SLICE_X101Y105_A3 = CLBLM_R_X65Y105_SLICE_X99Y105_BO5;
  assign CLBLM_L_X74Y131_SLICE_X112Y131_A6 = 1'b1;
  assign CLBLM_R_X67Y105_SLICE_X101Y105_A4 = CLBLM_R_X67Y105_SLICE_X101Y105_DO6;
  assign CLBLM_R_X67Y105_SLICE_X101Y105_A5 = CLBLM_R_X67Y105_SLICE_X100Y105_DO5;
  assign CLBLM_R_X67Y105_SLICE_X101Y105_A6 = CLBLM_R_X67Y105_SLICE_X101Y105_CO6;
  assign RIOB33_X105Y187_IOB_X1Y187_O = CLBLL_R_X73Y108_SLICE_X110Y108_AQ;
  assign RIOB33_X105Y187_IOB_X1Y188_O = CLBLL_R_X71Y117_SLICE_X106Y117_B5Q;
  assign CLBLM_R_X67Y105_SLICE_X101Y105_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y105_SLICE_X101Y105_B2 = CLBLM_L_X72Y104_SLICE_X108Y104_CQ;
  assign CLBLM_R_X67Y105_SLICE_X101Y105_B3 = CLBLM_L_X72Y105_SLICE_X109Y105_B5Q;
  assign CLBLM_R_X67Y105_SLICE_X101Y105_B4 = CLBLM_R_X67Y108_SLICE_X100Y108_BO6;
  assign CLBLM_R_X67Y105_SLICE_X101Y105_B5 = CLBLL_R_X71Y109_SLICE_X106Y109_AQ;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_A1 = CLBLM_L_X74Y122_SLICE_X112Y122_A5Q;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_A2 = CLBLL_R_X73Y122_SLICE_X110Y122_AO6;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_A3 = CLBLL_R_X73Y121_SLICE_X111Y121_AQ;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_A4 = CLBLL_R_X75Y128_SLICE_X114Y128_AO5;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_A6 = CLBLL_R_X73Y121_SLICE_X111Y121_BQ;
  assign CLBLM_R_X67Y105_SLICE_X101Y105_B6 = CLBLL_R_X71Y108_SLICE_X106Y108_D5Q;
  assign CLBLM_L_X74Y131_SLICE_X112Y131_AX = CLBLL_R_X73Y131_SLICE_X111Y131_AQ;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_B2 = CLBLL_R_X73Y121_SLICE_X111Y121_BQ;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_B3 = CLBLL_R_X73Y122_SLICE_X111Y122_AO6;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_B4 = CLBLL_R_X73Y121_SLICE_X110Y121_BQ;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_B5 = CLBLL_R_X75Y128_SLICE_X115Y128_BO6;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_B6 = CLBLL_R_X75Y128_SLICE_X114Y128_AO5;
  assign CLBLM_R_X67Y105_SLICE_X101Y105_C3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y105_SLICE_X101Y105_C4 = CLBLM_L_X68Y103_SLICE_X102Y103_DQ;
  assign CLBLM_L_X74Y131_SLICE_X112Y131_B1 = 1'b1;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_C1 = CLBLL_R_X73Y123_SLICE_X111Y123_AQ;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_C2 = CLBLL_R_X73Y122_SLICE_X110Y122_CQ;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_C3 = CLBLL_R_X73Y121_SLICE_X111Y121_BQ;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_C4 = CLBLM_L_X72Y122_SLICE_X109Y122_A5Q;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_C5 = CLBLM_L_X72Y122_SLICE_X109Y122_AQ;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_C6 = 1'b1;
  assign CLBLM_L_X74Y131_SLICE_X112Y131_B2 = 1'b1;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y131_SLICE_X112Y131_B3 = 1'b1;
  assign CLBLM_R_X67Y105_SLICE_X101Y105_D2 = CLBLM_R_X67Y105_SLICE_X100Y105_AO6;
  assign CLBLM_R_X67Y105_SLICE_X101Y105_D3 = CLBLM_R_X67Y105_SLICE_X100Y105_CO5;
  assign CLBLM_R_X67Y105_SLICE_X101Y105_D4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y131_SLICE_X112Y131_B4 = 1'b1;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_D1 = 1'b1;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_D2 = 1'b1;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_D3 = 1'b1;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_D4 = 1'b1;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_D5 = 1'b1;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_D6 = 1'b1;
  assign CLBLM_L_X74Y131_SLICE_X112Y131_B5 = 1'b1;
  assign CLBLM_R_X67Y105_SLICE_X100Y105_A1 = CLBLM_R_X67Y105_SLICE_X100Y105_DO6;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y131_SLICE_X112Y131_B6 = 1'b1;
  assign CLBLM_R_X67Y105_SLICE_X100Y105_A5 = CLBLM_R_X65Y101_SLICE_X99Y101_AO6;
  assign CLBLM_R_X67Y105_SLICE_X100Y105_A6 = CLBLM_R_X67Y108_SLICE_X100Y108_BO6;
  assign CLBLM_R_X67Y105_SLICE_X100Y105_B1 = CLBLM_R_X67Y105_SLICE_X100Y105_DO6;
  assign CLBLM_R_X67Y105_SLICE_X100Y105_B2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y105_SLICE_X100Y105_B3 = CLBLM_R_X67Y103_SLICE_X100Y103_AO6;
  assign CLBLM_R_X67Y105_SLICE_X100Y105_B4 = CLBLM_R_X67Y108_SLICE_X100Y108_BO6;
  assign CLBLM_R_X67Y105_SLICE_X100Y105_B5 = CLBLM_R_X65Y105_SLICE_X99Y105_AO6;
  assign CLBLM_R_X67Y105_SLICE_X100Y105_B6 = CLBLM_R_X67Y105_SLICE_X100Y105_CO6;
  assign CLBLM_R_X67Y105_SLICE_X100Y105_C1 = CLBLL_R_X71Y109_SLICE_X106Y109_AQ;
  assign CLBLM_R_X67Y105_SLICE_X100Y105_C2 = CLBLM_R_X65Y100_SLICE_X99Y100_CQ;
  assign CLBLM_R_X67Y105_SLICE_X100Y105_C3 = CLBLL_R_X71Y108_SLICE_X106Y108_D5Q;
  assign CLBLM_R_X67Y105_SLICE_X100Y105_C4 = CLBLM_R_X65Y100_SLICE_X99Y100_A5Q;
  assign CLBLM_R_X67Y105_SLICE_X100Y105_C5 = 1'b1;
  assign CLBLM_R_X67Y105_SLICE_X100Y105_C6 = 1'b1;
  assign CLBLM_R_X67Y105_SLICE_X100Y105_D1 = CLBLM_L_X72Y105_SLICE_X109Y105_B5Q;
  assign CLBLM_R_X67Y105_SLICE_X100Y105_D2 = CLBLM_R_X65Y105_SLICE_X98Y105_CQ;
  assign CLBLM_R_X67Y105_SLICE_X100Y105_D3 = CLBLM_L_X72Y104_SLICE_X108Y104_CQ;
  assign CLBLM_L_X74Y131_SLICE_X112Y131_C1 = 1'b1;
  assign CLBLM_R_X67Y105_SLICE_X100Y105_D4 = CLBLM_R_X65Y106_SLICE_X99Y106_C5Q;
  assign CLBLM_R_X67Y105_SLICE_X100Y105_D5 = 1'b1;
  assign CLBLM_R_X67Y105_SLICE_X100Y105_D6 = 1'b1;
  assign CLBLM_L_X74Y131_SLICE_X112Y131_C2 = 1'b1;
  assign CLBLM_L_X74Y131_SLICE_X112Y131_C3 = 1'b1;
  assign CLBLM_L_X74Y131_SLICE_X112Y131_C4 = 1'b1;
  assign CLBLM_L_X74Y131_SLICE_X112Y131_C5 = 1'b1;
  assign CLBLM_L_X74Y131_SLICE_X112Y131_C6 = 1'b1;
  assign CLBLL_R_X75Y133_SLICE_X114Y133_A1 = CLBLM_L_X74Y132_SLICE_X112Y132_C5Q;
  assign CLBLL_R_X75Y133_SLICE_X114Y133_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y133_SLICE_X114Y133_A3 = CLBLL_R_X75Y133_SLICE_X115Y133_AO6;
  assign CLBLL_R_X75Y133_SLICE_X114Y133_A4 = CLBLL_R_X75Y133_SLICE_X115Y133_BQ;
  assign CLBLL_R_X75Y133_SLICE_X114Y133_A5 = CLBLM_L_X74Y131_SLICE_X112Y131_AQ;
  assign CLBLL_R_X75Y133_SLICE_X114Y133_A6 = CLBLL_R_X75Y134_SLICE_X115Y134_AQ;
  assign CLBLM_L_X74Y131_SLICE_X112Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X75Y133_SLICE_X114Y133_B1 = CLBLL_R_X75Y133_SLICE_X114Y133_DO6;
  assign CLBLL_R_X75Y133_SLICE_X114Y133_B2 = CLBLM_L_X74Y129_SLICE_X112Y129_BQ;
  assign CLBLL_R_X75Y133_SLICE_X114Y133_B3 = CLBLM_L_X74Y132_SLICE_X112Y132_C5Q;
  assign CLBLL_R_X75Y133_SLICE_X114Y133_B4 = CLBLL_R_X79Y135_SLICE_X122Y135_AQ;
  assign CLBLL_R_X75Y133_SLICE_X114Y133_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y133_SLICE_X114Y133_B6 = CLBLL_R_X75Y133_SLICE_X114Y133_CO6;
  assign CLBLL_R_X75Y133_SLICE_X114Y133_C1 = CLBLL_R_X75Y133_SLICE_X114Y133_BQ;
  assign CLBLL_R_X75Y133_SLICE_X114Y133_C2 = CLBLM_L_X70Y136_SLICE_X105Y136_A5Q;
  assign CLBLL_R_X75Y133_SLICE_X114Y133_C3 = CLBLL_R_X75Y133_SLICE_X114Y133_AQ;
  assign CLBLL_R_X75Y133_SLICE_X114Y133_C4 = CLBLL_R_X75Y134_SLICE_X115Y134_AQ;
  assign CLBLL_R_X75Y133_SLICE_X114Y133_C5 = 1'b1;
  assign CLBLL_R_X75Y133_SLICE_X114Y133_C6 = 1'b1;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_A2 = CLBLM_L_X76Y124_SLICE_X116Y124_DQ;
  assign CLBLL_R_X75Y133_SLICE_X114Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X75Y133_SLICE_X114Y133_D1 = CLBLM_L_X74Y131_SLICE_X112Y131_AQ;
  assign CLBLL_R_X75Y133_SLICE_X114Y133_D2 = CLBLM_L_X74Y132_SLICE_X112Y132_C5Q;
  assign CLBLL_R_X75Y133_SLICE_X114Y133_D3 = CLBLL_R_X75Y133_SLICE_X115Y133_AQ;
  assign CLBLL_R_X75Y133_SLICE_X114Y133_D4 = CLBLL_R_X75Y134_SLICE_X115Y134_AQ;
  assign CLBLL_R_X75Y133_SLICE_X114Y133_D5 = CLBLM_L_X76Y133_SLICE_X116Y133_BQ;
  assign CLBLL_R_X75Y133_SLICE_X114Y133_D6 = CLBLL_R_X75Y133_SLICE_X115Y133_BQ;
  assign CLBLM_L_X74Y131_SLICE_X112Y131_D1 = 1'b1;
  assign CLBLL_R_X75Y133_SLICE_X114Y133_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y131_SLICE_X112Y131_D2 = 1'b1;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_A3 = CLBLL_R_X75Y122_SLICE_X115Y122_A5Q;
  assign CLBLM_L_X74Y131_SLICE_X112Y131_D3 = 1'b1;
  assign CLBLM_L_X74Y131_SLICE_X112Y131_D4 = 1'b1;
  assign CLBLM_L_X74Y131_SLICE_X112Y131_D5 = 1'b1;
  assign CLBLM_L_X74Y131_SLICE_X112Y131_D6 = 1'b1;
  assign CLBLL_R_X75Y133_SLICE_X115Y133_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y133_SLICE_X115Y133_A2 = CLBLL_R_X75Y134_SLICE_X114Y134_CO5;
  assign CLBLL_R_X75Y133_SLICE_X115Y133_A3 = CLBLL_R_X75Y133_SLICE_X115Y133_AQ;
  assign CLBLL_R_X75Y133_SLICE_X115Y133_A4 = CLBLL_R_X75Y134_SLICE_X115Y134_BO6;
  assign CLBLL_R_X75Y133_SLICE_X115Y133_A5 = CLBLM_L_X76Y133_SLICE_X116Y133_BQ;
  assign CLBLL_R_X75Y133_SLICE_X115Y133_A6 = 1'b1;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_A4 = CLBLL_R_X75Y124_SLICE_X115Y124_AQ;
  assign CLBLL_R_X75Y133_SLICE_X115Y133_B1 = 1'b1;
  assign CLBLL_R_X75Y133_SLICE_X115Y133_B2 = 1'b1;
  assign CLBLL_R_X75Y133_SLICE_X115Y133_B3 = 1'b1;
  assign CLBLL_R_X75Y133_SLICE_X115Y133_B4 = 1'b1;
  assign CLBLL_R_X75Y133_SLICE_X115Y133_B5 = 1'b1;
  assign CLBLL_R_X75Y133_SLICE_X115Y133_B6 = 1'b1;
  assign CLBLL_R_X75Y133_SLICE_X115Y133_BX = CLBLM_L_X74Y129_SLICE_X112Y129_BQ;
  assign LIOI3_X0Y51_OLOGIC_X0Y52_D1 = CLBLM_L_X68Y95_SLICE_X102Y95_A5Q;
  assign CLBLL_R_X75Y133_SLICE_X115Y133_C1 = 1'b1;
  assign CLBLL_R_X75Y133_SLICE_X115Y133_C2 = 1'b1;
  assign CLBLL_R_X75Y133_SLICE_X115Y133_C3 = 1'b1;
  assign CLBLL_R_X75Y133_SLICE_X115Y133_C4 = 1'b1;
  assign CLBLL_R_X75Y133_SLICE_X115Y133_C5 = 1'b1;
  assign CLBLL_R_X75Y133_SLICE_X115Y133_C6 = 1'b1;
  assign CLBLM_L_X74Y131_SLICE_X112Y131_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_A5 = CLBLM_L_X76Y122_SLICE_X116Y122_A5Q;
  assign CLBLL_R_X75Y133_SLICE_X115Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X75Y133_SLICE_X115Y133_D1 = 1'b1;
  assign CLBLL_R_X75Y133_SLICE_X115Y133_D2 = 1'b1;
  assign CLBLL_R_X75Y133_SLICE_X115Y133_D3 = 1'b1;
  assign CLBLL_R_X75Y133_SLICE_X115Y133_D4 = 1'b1;
  assign CLBLL_R_X75Y133_SLICE_X115Y133_D5 = 1'b1;
  assign CLBLL_R_X75Y133_SLICE_X115Y133_D6 = 1'b1;
  assign CLBLL_R_X75Y133_SLICE_X115Y133_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign LIOB33_X0Y103_IOB_X0Y104_O = RIOB33_X105Y53_IOB_X1Y53_I;
  assign LIOB33_X0Y103_IOB_X0Y103_O = RIOB33_X105Y55_IOB_X1Y56_I;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_A6 = 1'b1;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_A1 = CLBLM_L_X74Y122_SLICE_X112Y122_A5Q;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_A2 = CLBLM_L_X74Y122_SLICE_X112Y122_AQ;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_A3 = 1'b1;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_A4 = 1'b1;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_A5 = CLBLL_R_X75Y128_SLICE_X115Y128_BO6;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_A6 = 1'b1;
  assign CLBLM_L_X72Y134_SLICE_X109Y134_C3 = 1'b1;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_B1 = CLBLL_R_X73Y123_SLICE_X111Y123_CQ;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_B2 = CLBLL_R_X73Y122_SLICE_X110Y122_BQ;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_B4 = 1'b1;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_B5 = CLBLL_R_X75Y128_SLICE_X114Y128_AO5;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_B6 = CLBLL_R_X73Y122_SLICE_X110Y122_AO5;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_C1 = CLBLL_R_X73Y122_SLICE_X111Y122_AQ;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_C2 = CLBLL_R_X73Y122_SLICE_X110Y122_CQ;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_C3 = CLBLL_R_X75Y128_SLICE_X114Y128_AO5;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_C4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_C5 = CLBLL_R_X73Y122_SLICE_X110Y122_DO6;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_C6 = CLBLL_R_X73Y121_SLICE_X110Y121_AQ;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOB33_X105Y189_IOB_X1Y189_O = 1'b0;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_D1 = CLBLL_R_X73Y122_SLICE_X111Y122_AQ;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_D2 = CLBLM_L_X74Y122_SLICE_X112Y122_A5Q;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_D3 = 1'b1;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_D4 = CLBLL_R_X75Y128_SLICE_X115Y128_BO6;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_D5 = 1'b1;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_D6 = 1'b1;
  assign RIOB33_X105Y189_IOB_X1Y190_O = CLBLM_L_X76Y128_SLICE_X116Y128_C5Q;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_A1 = CLBLL_R_X75Y128_SLICE_X115Y128_BO6;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_A2 = CLBLM_L_X74Y122_SLICE_X112Y122_AQ;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_A3 = CLBLL_R_X73Y122_SLICE_X111Y122_AQ;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_A5 = CLBLL_R_X73Y123_SLICE_X110Y123_BQ;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_A6 = 1'b1;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_B2 = CLBLL_R_X73Y124_SLICE_X111Y124_BQ;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_B3 = CLBLL_R_X71Y124_SLICE_X106Y124_CO6;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_B4 = CLBLM_L_X72Y122_SLICE_X109Y122_AQ;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_B5 = CLBLM_L_X72Y122_SLICE_X109Y122_A5Q;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_B6 = CLBLL_R_X73Y122_SLICE_X111Y122_BQ;
  assign RIOB33_SING_X105Y149_IOB_X1Y149_O = CLBLM_L_X76Y111_SLICE_X116Y111_BQ;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_C2 = CLBLL_R_X73Y122_SLICE_X111Y122_CQ;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_C3 = CLBLM_L_X74Y122_SLICE_X112Y122_A5Q;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_C4 = CLBLL_R_X73Y122_SLICE_X111Y122_BQ;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_C5 = CLBLL_R_X75Y128_SLICE_X115Y128_BO6;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_C6 = CLBLM_L_X74Y122_SLICE_X112Y122_AQ;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_D1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_D2 = CLBLL_R_X73Y122_SLICE_X111Y122_CQ;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_D3 = CLBLL_R_X73Y122_SLICE_X111Y122_DQ;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_D4 = CLBLL_R_X73Y122_SLICE_X111Y122_BQ;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_D5 = CLBLL_R_X73Y122_SLICE_X110Y122_AO5;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_D6 = 1'b1;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_D5 = CLBLL_R_X77Y122_SLICE_X119Y122_AO5;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_D6 = CLBLM_L_X78Y122_SLICE_X121Y122_BQ;
  assign CLBLL_R_X75Y134_SLICE_X114Y134_A1 = 1'b1;
  assign CLBLL_R_X75Y134_SLICE_X114Y134_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y134_SLICE_X114Y134_A3 = CLBLL_R_X75Y134_SLICE_X114Y134_AQ;
  assign CLBLL_R_X75Y134_SLICE_X114Y134_A4 = CLBLM_L_X76Y134_SLICE_X117Y134_BQ;
  assign CLBLL_R_X75Y134_SLICE_X114Y134_A5 = CLBLL_R_X75Y134_SLICE_X114Y134_CO5;
  assign CLBLL_R_X75Y134_SLICE_X114Y134_A6 = CLBLL_R_X75Y133_SLICE_X115Y133_AQ;
  assign CLBLL_R_X75Y134_SLICE_X114Y134_AX = CLBLL_R_X75Y134_SLICE_X114Y134_BO6;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_T1 = 1'b1;
  assign CLBLL_R_X75Y134_SLICE_X114Y134_B1 = CLBLL_R_X75Y134_SLICE_X114Y134_A5Q;
  assign CLBLL_R_X75Y134_SLICE_X114Y134_B2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X75Y134_SLICE_X114Y134_B3 = CLBLL_R_X75Y134_SLICE_X114Y134_AQ;
  assign CLBLL_R_X75Y134_SLICE_X114Y134_B4 = CLBLL_R_X75Y133_SLICE_X115Y133_AQ;
  assign CLBLL_R_X75Y134_SLICE_X114Y134_B5 = CLBLL_R_X75Y134_SLICE_X114Y134_CO5;
  assign CLBLL_R_X75Y134_SLICE_X114Y134_B6 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_B4 = 1'b1;
  assign CLBLL_R_X75Y134_SLICE_X114Y134_C1 = CLBLL_R_X75Y133_SLICE_X115Y133_BQ;
  assign CLBLL_R_X75Y134_SLICE_X114Y134_C2 = CLBLL_R_X75Y134_SLICE_X115Y134_AQ;
  assign CLBLL_R_X75Y134_SLICE_X114Y134_C3 = CLBLM_L_X76Y133_SLICE_X116Y133_BQ;
  assign CLBLL_R_X75Y134_SLICE_X114Y134_C4 = CLBLM_L_X74Y132_SLICE_X112Y132_C5Q;
  assign CLBLL_R_X75Y134_SLICE_X114Y134_C5 = CLBLL_R_X75Y133_SLICE_X115Y133_AQ;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_B5 = 1'b1;
  assign CLBLL_R_X75Y134_SLICE_X114Y134_C6 = 1'b1;
  assign CLBLL_R_X75Y134_SLICE_X114Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_B6 = 1'b1;
  assign CLBLL_R_X75Y134_SLICE_X114Y134_D1 = 1'b1;
  assign CLBLL_R_X75Y134_SLICE_X114Y134_D2 = CLBLM_L_X74Y134_SLICE_X112Y134_BQ;
  assign CLBLL_R_X75Y134_SLICE_X114Y134_D3 = CLBLM_L_X74Y134_SLICE_X112Y134_CQ;
  assign CLBLL_R_X75Y134_SLICE_X114Y134_D4 = 1'b1;
  assign CLBLL_R_X75Y134_SLICE_X114Y134_D5 = 1'b1;
  assign CLBLL_R_X75Y134_SLICE_X114Y134_D6 = CLBLM_L_X74Y132_SLICE_X112Y132_C5Q;
  assign CLBLL_R_X75Y134_SLICE_X114Y134_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_C3 = 1'b1;
  assign CLBLL_R_X75Y134_SLICE_X115Y134_A1 = CLBLL_R_X75Y133_SLICE_X115Y133_BQ;
  assign CLBLL_R_X75Y134_SLICE_X115Y134_A2 = CLBLM_L_X76Y134_SLICE_X117Y134_BQ;
  assign CLBLL_R_X75Y134_SLICE_X115Y134_A3 = CLBLM_L_X76Y133_SLICE_X116Y133_AQ;
  assign CLBLL_R_X75Y134_SLICE_X115Y134_A4 = CLBLM_L_X76Y134_SLICE_X116Y134_BQ;
  assign CLBLL_R_X75Y134_SLICE_X115Y134_A5 = CLBLM_L_X74Y132_SLICE_X112Y132_C5Q;
  assign CLBLL_R_X75Y134_SLICE_X115Y134_A6 = 1'b1;
  assign CLBLL_R_X75Y134_SLICE_X115Y134_AX = CLBLL_R_X79Y135_SLICE_X122Y135_AQ;
  assign CLBLL_R_X75Y134_SLICE_X115Y134_B1 = CLBLL_R_X75Y134_SLICE_X115Y134_DO6;
  assign CLBLL_R_X75Y134_SLICE_X115Y134_B2 = CLBLL_R_X75Y134_SLICE_X115Y134_AQ;
  assign CLBLL_R_X75Y134_SLICE_X115Y134_B3 = CLBLL_R_X75Y133_SLICE_X115Y133_BQ;
  assign CLBLL_R_X75Y134_SLICE_X115Y134_B4 = CLBLL_R_X75Y134_SLICE_X114Y134_BO5;
  assign CLBLL_R_X75Y134_SLICE_X115Y134_B5 = CLBLM_L_X76Y133_SLICE_X116Y133_BQ;
  assign CLBLL_R_X75Y134_SLICE_X115Y134_B6 = CLBLM_L_X74Y132_SLICE_X112Y132_C5Q;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_B6 = 1'b1;
  assign CLBLL_R_X75Y134_SLICE_X115Y134_C1 = CLBLL_R_X75Y133_SLICE_X114Y133_BQ;
  assign CLBLL_R_X75Y134_SLICE_X115Y134_C2 = CLBLL_R_X75Y133_SLICE_X115Y133_AQ;
  assign CLBLL_R_X75Y134_SLICE_X115Y134_C3 = CLBLL_R_X75Y134_SLICE_X114Y134_DO6;
  assign CLBLL_R_X75Y134_SLICE_X115Y134_C4 = CLBLL_R_X75Y134_SLICE_X115Y134_AO5;
  assign CLBLL_R_X75Y134_SLICE_X115Y134_C5 = CLBLM_L_X76Y133_SLICE_X116Y133_BQ;
  assign CLBLL_R_X75Y134_SLICE_X115Y134_C6 = CLBLL_R_X75Y134_SLICE_X115Y134_DO5;
  assign LIOB33_X0Y105_IOB_X0Y105_O = RIOB33_X105Y53_IOB_X1Y54_I;
  assign LIOB33_X0Y105_IOB_X0Y106_O = RIOB33_X105Y59_IOB_X1Y60_I;
  assign CLBLL_R_X75Y134_SLICE_X115Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X75Y134_SLICE_X115Y134_D1 = CLBLM_L_X76Y134_SLICE_X116Y134_AQ;
  assign CLBLL_R_X75Y134_SLICE_X115Y134_D2 = 1'b1;
  assign CLBLL_R_X75Y134_SLICE_X115Y134_D3 = CLBLM_L_X76Y134_SLICE_X117Y134_AQ;
  assign CLBLL_R_X75Y134_SLICE_X115Y134_D4 = CLBLL_R_X75Y133_SLICE_X115Y133_BQ;
  assign CLBLL_R_X75Y134_SLICE_X115Y134_D5 = CLBLL_R_X75Y134_SLICE_X115Y134_AQ;
  assign CLBLL_R_X75Y134_SLICE_X115Y134_D6 = 1'b1;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE = 1'b1;
  assign CLBLL_R_X75Y134_SLICE_X115Y134_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_CE = 1'b1;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_A1 = 1'b1;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_A2 = 1'b1;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_A3 = 1'b1;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_A4 = 1'b1;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_A5 = 1'b1;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_A6 = 1'b1;
  assign RIOB33_X105Y191_IOB_X1Y192_O = CLBLM_L_X72Y118_SLICE_X109Y118_A5Q;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_AX = CLBLL_R_X75Y124_SLICE_X114Y124_C5Q;
  assign RIOB33_X105Y191_IOB_X1Y191_O = CLBLM_L_X68Y109_SLICE_X102Y109_AQ;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_B1 = 1'b1;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_B2 = 1'b1;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_B3 = 1'b1;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_B4 = 1'b1;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_B5 = 1'b1;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_B6 = 1'b1;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_BX = CLBLM_L_X74Y122_SLICE_X112Y122_AQ;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_C1 = 1'b1;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_C2 = 1'b1;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_C3 = 1'b1;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_C4 = 1'b1;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_C5 = 1'b1;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_C6 = 1'b1;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_CE = CLBLM_L_X76Y109_SLICE_X116Y109_AO6;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_D6 = 1'b1;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_CX = CLBLL_R_X73Y123_SLICE_X111Y123_AQ;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_D1 = CLBLM_L_X64Y105_SLICE_X97Y105_DO6;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_D1 = 1'b1;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_D2 = 1'b1;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_D3 = 1'b1;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_D4 = 1'b1;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_D5 = 1'b1;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_D6 = 1'b1;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_T1 = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_D1 = 1'b1;
  assign LIOI3_X0Y73_OLOGIC_X0Y74_D1 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_A1 = CLBLL_R_X73Y123_SLICE_X111Y123_AQ;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_A2 = CLBLL_R_X71Y124_SLICE_X106Y124_CO6;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_A3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_A4 = CLBLM_L_X72Y122_SLICE_X109Y122_AQ;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_A5 = 1'b1;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_A6 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_A4 = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_T1 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_A5 = 1'b1;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_B1 = CLBLM_L_X74Y122_SLICE_X112Y122_A5Q;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_B2 = CLBLL_R_X73Y123_SLICE_X111Y123_BQ;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_B3 = CLBLM_L_X74Y122_SLICE_X112Y122_AQ;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_B4 = CLBLL_R_X75Y128_SLICE_X115Y128_BO6;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_B6 = CLBLM_L_X74Y128_SLICE_X113Y128_AO5;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_A6 = 1'b1;
  assign LIOI3_X0Y73_OLOGIC_X0Y74_T1 = 1'b1;
  assign RIOI3_X105Y117_OLOGIC_X1Y118_D1 = CLBLM_L_X70Y136_SLICE_X105Y136_A5Q;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_C1 = CLBLM_L_X74Y122_SLICE_X112Y122_AQ;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_C2 = CLBLL_R_X73Y123_SLICE_X111Y123_CQ;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_C3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_C4 = CLBLL_R_X73Y123_SLICE_X111Y123_BQ;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_C5 = CLBLM_L_X74Y122_SLICE_X112Y122_A5Q;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_C6 = CLBLL_R_X75Y128_SLICE_X115Y128_BO6;
  assign LIOI3_X0Y73_OLOGIC_X0Y73_D1 = CLBLM_L_X62Y105_SLICE_X93Y105_A5Q;
  assign RIOI3_X105Y117_OLOGIC_X1Y118_T1 = 1'b1;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_D1 = CLBLM_L_X76Y125_SLICE_X116Y125_AQ;
  assign LIOI3_X0Y73_OLOGIC_X0Y73_T1 = 1'b1;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_D1 = CLBLM_L_X74Y122_SLICE_X112Y122_AQ;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_D2 = CLBLM_L_X74Y122_SLICE_X112Y122_A5Q;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_D3 = CLBLL_R_X73Y123_SLICE_X111Y123_DQ;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_D4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_D5 = CLBLL_R_X73Y122_SLICE_X111Y122_DQ;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_D6 = CLBLL_R_X75Y128_SLICE_X115Y128_BO6;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_T1 = 1'b1;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_C1 = CLBLM_L_X76Y124_SLICE_X116Y124_AO6;
  assign RIOI3_X105Y117_OLOGIC_X1Y117_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_D1 = CLBLM_R_X63Y122_SLICE_X95Y122_CQ;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_B3 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_B4 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_B5 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_T1 = 1'b1;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_B6 = 1'b1;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_C2 = CLBLM_L_X76Y122_SLICE_X116Y122_C5Q;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_T1 = 1'b1;
  assign RIOB33_X105Y101_IOB_X1Y101_O = CLBLM_L_X72Y109_SLICE_X109Y109_DQ;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOI3_X105Y117_OLOGIC_X1Y117_D1 = CLBLL_R_X73Y118_SLICE_X111Y118_AQ;
  assign LIOB33_X0Y71_IOB_X0Y72_O = CLBLM_L_X60Y104_SLICE_X90Y104_AQ;
  assign LIOB33_X0Y107_IOB_X0Y108_O = CLBLM_L_X70Y110_SLICE_X104Y110_CQ;
  assign LIOB33_X0Y107_IOB_X0Y107_O = RIOB33_X105Y55_IOB_X1Y55_I;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_D6 = 1'b1;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_A2 = CLBLM_L_X74Y127_SLICE_X112Y127_BQ;
  assign RIOB33_X105Y193_IOB_X1Y194_O = CLBLM_L_X76Y129_SLICE_X116Y129_CQ;
  assign RIOB33_X105Y193_IOB_X1Y193_O = 1'b0;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_A1 = CLBLM_L_X72Y124_SLICE_X108Y124_BO6;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_A2 = CLBLL_R_X73Y126_SLICE_X110Y126_AQ;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_A3 = CLBLL_R_X73Y124_SLICE_X110Y124_AQ;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_A4 = CLBLL_R_X73Y124_SLICE_X110Y124_BO6;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_A6 = CLBLM_L_X74Y126_SLICE_X112Y126_CO6;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_AX = CLBLL_R_X73Y124_SLICE_X110Y124_CO6;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_B1 = CLBLM_L_X72Y124_SLICE_X108Y124_BO6;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_B2 = CLBLL_R_X73Y124_SLICE_X110Y124_BQ;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_B4 = CLBLL_R_X73Y125_SLICE_X110Y125_AQ;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_B5 = CLBLL_R_X73Y124_SLICE_X110Y124_A5Q;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_B6 = 1'b1;
  assign LIOB33_X0Y167_IOB_X0Y168_O = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_C2 = CLBLM_L_X72Y124_SLICE_X108Y124_BO6;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_C3 = 1'b1;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_C4 = CLBLL_R_X73Y124_SLICE_X110Y124_A5Q;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_C5 = CLBLM_L_X72Y124_SLICE_X109Y124_AQ;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_C6 = 1'b1;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOB33_X105Y101_IOB_X1Y102_O = CLBLL_R_X73Y131_SLICE_X111Y131_AQ;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_D1 = 1'b1;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_D2 = 1'b1;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_D3 = 1'b1;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_D4 = 1'b1;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_D5 = 1'b1;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_D6 = 1'b1;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign LIOB33_X0Y167_IOB_X0Y167_O = CLBLL_L_X34Y126_SLICE_X50Y126_AO6;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_A2 = CLBLL_R_X73Y123_SLICE_X111Y123_AQ;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_A3 = CLBLL_R_X73Y124_SLICE_X111Y124_AQ;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_A4 = CLBLM_L_X72Y122_SLICE_X109Y122_AQ;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_A5 = CLBLM_L_X72Y123_SLICE_X108Y123_AQ;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_A6 = CLBLL_R_X71Y124_SLICE_X106Y124_CO6;
  assign CLBLM_R_X67Y108_SLICE_X101Y108_A1 = CLBLM_L_X68Y109_SLICE_X102Y109_A5Q;
  assign CLBLM_R_X67Y108_SLICE_X101Y108_A2 = CLBLM_L_X68Y108_SLICE_X102Y108_A5Q;
  assign CLBLM_R_X67Y108_SLICE_X101Y108_A3 = CLBLM_L_X68Y108_SLICE_X102Y108_AQ;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_B1 = 1'b1;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_B2 = CLBLL_R_X73Y124_SLICE_X111Y124_BQ;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_B3 = CLBLL_R_X73Y124_SLICE_X111Y124_AQ;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_B4 = CLBLL_R_X73Y123_SLICE_X111Y123_AO5;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_B5 = CLBLL_R_X73Y123_SLICE_X111Y123_CQ;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_B6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y108_SLICE_X101Y108_B1 = CLBLM_R_X67Y109_SLICE_X100Y109_BQ;
  assign CLBLM_R_X67Y108_SLICE_X101Y108_B2 = CLBLM_R_X67Y108_SLICE_X101Y108_BQ;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_C1 = 1'b1;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_C2 = 1'b1;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_C3 = 1'b1;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_C4 = 1'b1;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_C5 = 1'b1;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_C6 = 1'b1;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_A2 = CLBLM_L_X64Y97_SLICE_X96Y97_AQ;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_A3 = CLBLM_R_X63Y96_SLICE_X95Y96_AQ;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_A4 = CLBLM_L_X64Y97_SLICE_X97Y97_BO5;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_A5 = CLBLM_R_X63Y99_SLICE_X94Y99_BO5;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_A6 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_D1 = 1'b1;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_D2 = 1'b1;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_D3 = 1'b1;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_D4 = 1'b1;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_D5 = 1'b1;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_D6 = 1'b1;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_B3 = CLBLM_R_X63Y99_SLICE_X94Y99_BO5;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_B4 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_B5 = CLBLM_R_X63Y96_SLICE_X95Y96_BQ;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_B6 = CLBLM_L_X64Y97_SLICE_X96Y97_CQ;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_C1 = CLBLM_L_X64Y97_SLICE_X97Y97_BO5;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_C2 = CLBLM_R_X63Y96_SLICE_X95Y96_CQ;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_C3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_C4 = CLBLM_R_X63Y99_SLICE_X94Y99_CO6;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_C5 = CLBLM_R_X63Y96_SLICE_X95Y96_AQ;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_C6 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X67Y108_SLICE_X100Y108_A1 = CLBLM_R_X67Y108_SLICE_X101Y108_AO6;
  assign CLBLM_R_X67Y108_SLICE_X100Y108_A2 = CLBLM_L_X72Y105_SLICE_X108Y105_AQ;
  assign CLBLM_R_X67Y108_SLICE_X100Y108_A3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_D1 = CLBLM_R_X63Y96_SLICE_X95Y96_BQ;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_D2 = CLBLM_R_X63Y99_SLICE_X94Y99_CO6;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_D3 = CLBLM_R_X63Y96_SLICE_X95Y96_DQ;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_D4 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_D5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_D6 = CLBLM_L_X64Y98_SLICE_X96Y98_AO6;
  assign CLBLM_R_X67Y108_SLICE_X100Y108_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X67Y108_SLICE_X100Y108_B2 = CLBLM_R_X67Y108_SLICE_X100Y108_DQ;
  assign CLBLM_R_X67Y108_SLICE_X100Y108_B3 = CLBLL_R_X71Y109_SLICE_X106Y109_AQ;
  assign CLBLM_R_X67Y108_SLICE_X100Y108_B4 = CLBLL_R_X71Y108_SLICE_X106Y108_D5Q;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_A1 = CLBLM_R_X63Y99_SLICE_X94Y99_BO6;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_A2 = CLBLM_L_X64Y97_SLICE_X96Y97_BQ;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_A3 = CLBLM_R_X63Y96_SLICE_X94Y96_AQ;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_A4 = CLBLM_L_X64Y97_SLICE_X97Y97_BO6;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_A6 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X67Y108_SLICE_X100Y108_C1 = CLBLM_R_X67Y108_SLICE_X100Y108_C5Q;
  assign CLBLM_R_X67Y108_SLICE_X100Y108_C2 = CLBLM_R_X67Y108_SLICE_X100Y108_CQ;
  assign CLBLM_R_X67Y108_SLICE_X100Y108_C3 = CLBLM_R_X67Y108_SLICE_X101Y108_AO6;
  assign CLBLM_R_X67Y108_SLICE_X100Y108_C4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_B2 = CLBLM_R_X63Y96_SLICE_X94Y96_BQ;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_B3 = CLBLM_R_X63Y96_SLICE_X94Y96_AQ;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_B4 = CLBLM_L_X64Y97_SLICE_X97Y97_BO6;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_B5 = CLBLM_R_X63Y99_SLICE_X94Y99_BO5;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_B6 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X67Y108_SLICE_X100Y108_D1 = CLBLM_R_X67Y111_SLICE_X100Y111_CO5;
  assign CLBLM_R_X67Y108_SLICE_X100Y108_D2 = CLBLM_R_X67Y108_SLICE_X100Y108_AQ;
  assign CLBLM_R_X67Y108_SLICE_X100Y108_D3 = CLBLM_R_X67Y108_SLICE_X100Y108_DQ;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_C1 = 1'b1;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_C2 = 1'b1;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_C3 = 1'b1;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_C4 = 1'b1;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_C5 = 1'b1;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_C6 = 1'b1;
  assign CLBLM_R_X67Y108_SLICE_X100Y108_D6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y108_SLICE_X100Y108_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign RIOI3_X105Y101_OLOGIC_X1Y102_D1 = CLBLL_R_X73Y131_SLICE_X111Y131_AQ;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_D1 = 1'b1;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_D2 = 1'b1;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_D3 = 1'b1;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_D4 = 1'b1;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_D5 = 1'b1;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_D6 = 1'b1;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_A4 = CLBLM_L_X74Y127_SLICE_X113Y127_A5Q;
  assign LIOB33_X0Y109_IOB_X0Y110_O = CLBLL_R_X77Y129_SLICE_X118Y129_AQ;
  assign LIOB33_X0Y109_IOB_X0Y109_O = CLBLL_R_X75Y133_SLICE_X114Y133_AQ;
  assign RIOB33_X105Y195_IOB_X1Y196_O = 1'b0;
  assign RIOB33_X105Y195_IOB_X1Y195_O = CLBLL_R_X73Y104_SLICE_X110Y104_AQ;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_A1 = CLBLL_R_X73Y125_SLICE_X110Y125_BO6;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_A2 = CLBLL_R_X73Y124_SLICE_X110Y124_BQ;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_A3 = CLBLL_R_X73Y126_SLICE_X111Y126_CQ;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_A4 = CLBLM_L_X72Y124_SLICE_X109Y124_AQ;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_A5 = CLBLL_R_X73Y126_SLICE_X110Y126_AQ;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_A6 = CLBLL_R_X73Y125_SLICE_X110Y125_CO6;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_AX = CLBLL_R_X73Y124_SLICE_X110Y124_A5Q;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_B1 = CLBLM_L_X74Y126_SLICE_X112Y126_AQ;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_B2 = CLBLL_R_X73Y124_SLICE_X110Y124_BQ;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_B3 = 1'b1;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_B4 = CLBLL_R_X73Y126_SLICE_X111Y126_DQ;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_B5 = CLBLL_R_X73Y124_SLICE_X110Y124_A5Q;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_B6 = CLBLM_L_X72Y124_SLICE_X109Y124_AQ;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_C1 = CLBLL_R_X73Y124_SLICE_X110Y124_A5Q;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_C2 = 1'b1;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_C3 = CLBLL_R_X73Y126_SLICE_X111Y126_AQ;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_C4 = CLBLM_L_X72Y124_SLICE_X109Y124_AQ;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_C5 = CLBLM_L_X74Y126_SLICE_X112Y126_DQ;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_C6 = CLBLL_R_X73Y124_SLICE_X110Y124_BQ;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_CE = CLBLM_L_X76Y109_SLICE_X116Y109_AO6;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_D1 = CLBLL_R_X73Y123_SLICE_X110Y123_BQ;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_D2 = CLBLM_L_X72Y127_SLICE_X109Y127_BQ;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_D3 = CLBLL_R_X73Y125_SLICE_X110Y125_AQ;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_D4 = CLBLM_L_X74Y125_SLICE_X112Y125_BO6;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_D5 = 1'b1;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_D6 = CLBLM_L_X72Y127_SLICE_X109Y127_AQ;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign RIOB33_X105Y147_IOB_X1Y148_O = CLBLM_L_X62Y103_SLICE_X92Y103_B5Q;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_A1 = CLBLM_L_X70Y125_SLICE_X104Y125_BQ;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_A2 = CLBLM_L_X70Y125_SLICE_X105Y125_CO6;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_A3 = CLBLL_R_X75Y124_SLICE_X114Y124_AQ;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_A4 = CLBLM_L_X74Y125_SLICE_X112Y125_AO6;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_A6 = 1'b1;
  assign CLBLM_R_X67Y109_SLICE_X101Y109_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y109_SLICE_X101Y109_A2 = CLBLM_R_X67Y109_SLICE_X101Y109_BQ;
  assign CLBLM_R_X67Y109_SLICE_X101Y109_A3 = CLBLM_R_X67Y109_SLICE_X101Y109_AQ;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_B1 = CLBLM_L_X74Y126_SLICE_X113Y126_AQ;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_B2 = CLBLL_R_X73Y125_SLICE_X111Y125_BQ;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_B3 = CLBLM_L_X72Y125_SLICE_X109Y125_BQ;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_B4 = CLBLL_R_X75Y128_SLICE_X115Y128_AO6;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_B6 = CLBLM_L_X74Y126_SLICE_X113Y126_A5Q;
  assign CLBLM_R_X67Y109_SLICE_X101Y109_A4 = CLBLM_R_X67Y111_SLICE_X101Y111_B5Q;
  assign CLBLM_R_X67Y109_SLICE_X101Y109_A5 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X67Y109_SLICE_X101Y109_A6 = CLBLM_R_X65Y110_SLICE_X99Y110_AO5;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_C2 = CLBLL_R_X73Y125_SLICE_X111Y125_CQ;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_C3 = CLBLL_R_X73Y126_SLICE_X111Y126_BO5;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_C4 = CLBLL_R_X73Y125_SLICE_X111Y125_BQ;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_C5 = 1'b1;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_C6 = CLBLM_L_X72Y125_SLICE_X109Y125_BQ;
  assign CLBLM_R_X67Y109_SLICE_X101Y109_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y109_SLICE_X101Y109_B4 = CLBLM_R_X67Y111_SLICE_X101Y111_DO5;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_A1 = CLBLM_R_X63Y96_SLICE_X95Y96_AQ;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_A2 = CLBLM_R_X63Y97_SLICE_X94Y97_B5Q;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_A3 = CLBLM_R_X63Y97_SLICE_X95Y97_AQ;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_A4 = CLBLM_R_X63Y99_SLICE_X95Y99_BQ;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_A5 = CLBLM_R_X63Y99_SLICE_X95Y99_B5Q;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_D1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_D2 = CLBLL_R_X73Y125_SLICE_X111Y125_CQ;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_D3 = CLBLL_R_X73Y125_SLICE_X111Y125_DQ;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_D4 = CLBLM_L_X74Y126_SLICE_X113Y126_AQ;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_D5 = CLBLM_L_X74Y126_SLICE_X113Y126_A5Q;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_D6 = CLBLL_R_X75Y128_SLICE_X115Y128_AO6;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_A6 = CLBLM_L_X64Y97_SLICE_X96Y97_DQ;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_AX = CLBLM_R_X63Y98_SLICE_X94Y98_AQ;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_B1 = CLBLM_L_X64Y97_SLICE_X96Y97_CQ;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_B2 = CLBLM_L_X64Y97_SLICE_X97Y97_CQ;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_B3 = CLBLM_R_X63Y98_SLICE_X94Y98_AQ;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_B4 = CLBLM_R_X63Y99_SLICE_X95Y99_BQ;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_B5 = CLBLM_R_X63Y99_SLICE_X95Y99_B5Q;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_B6 = CLBLM_R_X63Y97_SLICE_X94Y97_CQ;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_C1 = CLBLM_R_X63Y99_SLICE_X95Y99_B5Q;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_C2 = CLBLM_L_X60Y92_SLICE_X90Y92_BQ;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_C3 = CLBLM_L_X64Y97_SLICE_X97Y97_DQ;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_C4 = CLBLM_R_X63Y97_SLICE_X94Y97_B5Q;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_C5 = CLBLM_R_X63Y99_SLICE_X95Y99_BQ;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_C6 = CLBLM_R_X63Y97_SLICE_X94Y97_BQ;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X67Y109_SLICE_X100Y109_A1 = CLBLM_R_X67Y111_SLICE_X100Y111_AQ;
  assign CLBLM_R_X67Y109_SLICE_X100Y109_A2 = 1'b1;
  assign CLBLM_R_X67Y109_SLICE_X100Y109_A3 = CLBLM_R_X67Y109_SLICE_X100Y109_AQ;
  assign CLBLM_R_X67Y109_SLICE_X100Y109_A4 = CLBLM_L_X68Y109_SLICE_X102Y109_CO6;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_D1 = CLBLM_R_X63Y97_SLICE_X95Y97_AO6;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_D2 = CLBLM_R_X63Y98_SLICE_X94Y98_AQ;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_D3 = CLBLM_L_X64Y97_SLICE_X97Y97_A5Q;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_D4 = CLBLM_R_X63Y99_SLICE_X95Y99_BQ;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_D5 = CLBLM_R_X63Y99_SLICE_X95Y99_B5Q;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_D6 = CLBLM_L_X64Y97_SLICE_X96Y97_AQ;
  assign CLBLM_R_X67Y109_SLICE_X100Y109_B1 = CLBLM_R_X67Y111_SLICE_X100Y111_AQ;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X67Y109_SLICE_X100Y109_B2 = CLBLM_R_X67Y109_SLICE_X100Y109_BQ;
  assign CLBLM_R_X67Y109_SLICE_X100Y109_B3 = CLBLM_R_X67Y109_SLICE_X100Y109_AQ;
  assign CLBLM_R_X67Y109_SLICE_X100Y109_B4 = 1'b1;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_A1 = CLBLM_L_X64Y97_SLICE_X97Y97_A5Q;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_A2 = CLBLM_R_X63Y99_SLICE_X95Y99_B5Q;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_A3 = CLBLM_L_X64Y97_SLICE_X96Y97_BQ;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_A4 = CLBLM_R_X63Y99_SLICE_X95Y99_BQ;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_A5 = CLBLM_R_X63Y97_SLICE_X94Y97_CQ;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_A6 = 1'b1;
  assign CLBLM_R_X67Y109_SLICE_X100Y109_C1 = CLBLM_R_X67Y111_SLICE_X101Y111_B5Q;
  assign CLBLM_R_X67Y109_SLICE_X100Y109_C2 = CLBLM_R_X67Y109_SLICE_X100Y109_CQ;
  assign CLBLM_R_X67Y109_SLICE_X100Y109_C3 = CLBLM_R_X67Y111_SLICE_X101Y111_A5Q;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_AX = CLBLM_R_X63Y97_SLICE_X95Y97_AQ;
  assign CLBLM_R_X67Y109_SLICE_X100Y109_C4 = CLBLM_R_X67Y111_SLICE_X100Y111_A5Q;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_B2 = CLBLM_R_X63Y97_SLICE_X94Y97_BQ;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_B3 = CLBLM_L_X64Y97_SLICE_X97Y97_BO6;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_B4 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_B5 = CLBLM_L_X62Y97_SLICE_X93Y97_BQ;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_B6 = CLBLM_R_X63Y99_SLICE_X94Y99_A5Q;
  assign CLBLM_R_X67Y109_SLICE_X100Y109_D1 = CLBLM_R_X65Y111_SLICE_X98Y111_AQ;
  assign CLBLM_R_X67Y109_SLICE_X100Y109_D2 = CLBLM_L_X68Y109_SLICE_X102Y109_A5Q;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_BX = CLBLM_R_X63Y97_SLICE_X94Y97_AQ;
  assign CLBLM_R_X67Y109_SLICE_X100Y109_D3 = CLBLM_L_X76Y111_SLICE_X116Y111_AQ;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_C1 = CLBLM_L_X62Y97_SLICE_X93Y97_BQ;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_C2 = CLBLM_R_X63Y99_SLICE_X95Y99_BQ;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_C3 = CLBLM_R_X63Y98_SLICE_X94Y98_BQ;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_C4 = CLBLM_L_X62Y97_SLICE_X93Y97_AQ;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_C5 = CLBLM_R_X63Y99_SLICE_X95Y99_B5Q;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_C6 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_R_X67Y109_SLICE_X100Y109_D6 = 1'b1;
  assign CLBLM_R_X67Y109_SLICE_X100Y109_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_T1 = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_D1 = 1'b1;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_CX = CLBLM_R_X63Y97_SLICE_X94Y97_B5Q;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_D1 = CLBLM_R_X63Y97_SLICE_X95Y97_AQ;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_D2 = CLBLM_L_X64Y98_SLICE_X96Y98_BQ;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_D3 = CLBLM_R_X63Y97_SLICE_X95Y97_BO6;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_D4 = CLBLM_R_X63Y97_SLICE_X94Y97_AO5;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_D5 = CLBLM_L_X62Y99_SLICE_X93Y99_AQ;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_D6 = CLBLM_R_X63Y96_SLICE_X95Y96_BQ;
  assign LIOI3_X0Y75_OLOGIC_X0Y76_D1 = CLBLM_L_X60Y99_SLICE_X90Y99_AQ;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_T1 = 1'b1;
  assign LIOB33_X0Y111_IOB_X0Y112_O = CLBLM_L_X64Y99_SLICE_X97Y99_B5Q;
  assign LIOB33_X0Y111_IOB_X0Y111_O = CLBLM_R_X65Y106_SLICE_X99Y106_DQ;
  assign LIOI3_X0Y75_OLOGIC_X0Y76_T1 = 1'b1;
  assign RIOI3_X105Y121_OLOGIC_X1Y122_D1 = CLBLM_R_X63Y98_SLICE_X94Y98_AQ;
  assign LIOI3_X0Y75_OLOGIC_X0Y75_D1 = CLBLM_L_X60Y101_SLICE_X90Y101_BQ;
  assign RIOI3_X105Y121_OLOGIC_X1Y122_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_D1 = CLBLM_L_X74Y120_SLICE_X112Y120_AO6;
  assign LIOI3_X0Y75_OLOGIC_X0Y75_T1 = 1'b1;
  assign CLBLM_L_X76Y118_SLICE_X117Y118_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign RIOI3_X105Y121_OLOGIC_X1Y121_D1 = CLBLM_L_X70Y100_SLICE_X104Y100_A5Q;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_T1 = 1'b1;
  assign RIOB33_X105Y197_IOB_X1Y198_O = CLBLM_L_X80Y132_SLICE_X124Y132_AQ;
  assign RIOB33_X105Y197_IOB_X1Y197_O = CLBLL_R_X79Y135_SLICE_X122Y135_AQ;
  assign RIOI3_X105Y121_OLOGIC_X1Y121_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_D1 = CLBLL_R_X73Y131_SLICE_X110Y131_AQ;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_T1 = 1'b1;
  assign CLBLM_L_X76Y118_SLICE_X116Y118_A5 = CLBLM_L_X76Y118_SLICE_X117Y118_AQ;
  assign CLBLM_L_X76Y118_SLICE_X116Y118_A6 = 1'b1;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_A1 = CLBLL_R_X73Y126_SLICE_X111Y126_DQ;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_A2 = CLBLL_R_X73Y126_SLICE_X111Y126_BO6;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_A3 = CLBLL_R_X73Y126_SLICE_X110Y126_AQ;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_A4 = CLBLM_L_X74Y126_SLICE_X113Y126_A5Q;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_A6 = CLBLL_R_X75Y128_SLICE_X114Y128_AO6;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_AX = CLBLL_R_X73Y126_SLICE_X110Y126_CO5;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_B1 = CLBLL_R_X73Y127_SLICE_X110Y127_CO6;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_B2 = CLBLL_R_X73Y126_SLICE_X110Y126_BQ;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_B3 = CLBLL_R_X71Y126_SLICE_X106Y126_CO6;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_B4 = CLBLL_R_X73Y127_SLICE_X110Y127_AQ;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_B6 = CLBLL_R_X73Y126_SLICE_X110Y126_CO6;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_C1 = CLBLL_R_X71Y126_SLICE_X106Y126_CO6;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_C2 = CLBLL_R_X71Y127_SLICE_X107Y127_AQ;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_C3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_C4 = CLBLL_R_X73Y126_SLICE_X110Y126_A5Q;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_C5 = CLBLM_L_X74Y127_SLICE_X112Y127_AQ;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_C6 = 1'b1;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_D1 = CLBLL_R_X71Y126_SLICE_X106Y126_CO6;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_D2 = CLBLL_R_X71Y127_SLICE_X107Y127_DQ;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_D3 = CLBLL_R_X73Y126_SLICE_X110Y126_DQ;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_D4 = CLBLL_R_X73Y126_SLICE_X110Y126_A5Q;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_D5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_D6 = CLBLM_L_X72Y126_SLICE_X109Y126_AQ;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X76Y118_SLICE_X116Y118_C1 = 1'b1;
  assign CLBLM_L_X76Y118_SLICE_X116Y118_C2 = 1'b1;
  assign CLBLM_L_X76Y118_SLICE_X116Y118_C5 = 1'b1;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_A1 = CLBLM_L_X74Y126_SLICE_X112Y126_A5Q;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_A2 = CLBLL_R_X73Y126_SLICE_X111Y126_CQ;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_A3 = CLBLL_R_X73Y126_SLICE_X111Y126_AQ;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_A4 = CLBLL_R_X73Y126_SLICE_X111Y126_BO6;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_A6 = CLBLL_R_X75Y128_SLICE_X114Y128_AO6;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_B1 = CLBLM_L_X74Y126_SLICE_X113Y126_AQ;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_B2 = CLBLM_L_X74Y126_SLICE_X113Y126_A5Q;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_B3 = 1'b1;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_B4 = 1'b1;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_B5 = CLBLL_R_X75Y128_SLICE_X115Y128_AO6;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_B6 = 1'b1;
  assign CLBLM_R_X67Y110_SLICE_X101Y110_A1 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X67Y110_SLICE_X101Y110_A2 = CLBLM_R_X65Y110_SLICE_X99Y110_AO6;
  assign CLBLM_R_X67Y110_SLICE_X101Y110_A3 = CLBLM_R_X67Y110_SLICE_X101Y110_AQ;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_C2 = CLBLL_R_X73Y126_SLICE_X111Y126_CQ;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_C3 = CLBLM_L_X74Y126_SLICE_X113Y126_CQ;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_C4 = CLBLL_R_X75Y128_SLICE_X114Y128_AO6;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_C5 = CLBLL_R_X73Y126_SLICE_X111Y126_BO5;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_C6 = 1'b1;
  assign CLBLM_R_X67Y110_SLICE_X101Y110_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X67Y110_SLICE_X101Y110_B2 = CLBLM_R_X67Y110_SLICE_X101Y110_BQ;
  assign CLBLM_R_X67Y110_SLICE_X101Y110_B3 = CLBLM_R_X67Y110_SLICE_X101Y110_AQ;
  assign CLBLM_R_X67Y110_SLICE_X101Y110_B4 = CLBLM_R_X67Y111_SLICE_X101Y111_CO5;
  assign CLBLM_R_X67Y110_SLICE_X101Y110_B5 = CLBLM_R_X65Y110_SLICE_X99Y110_AO6;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_A1 = CLBLM_R_X63Y97_SLICE_X94Y97_DO6;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_D1 = CLBLL_R_X75Y128_SLICE_X115Y128_AO6;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_D2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_D3 = CLBLL_R_X73Y126_SLICE_X111Y126_DQ;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_D4 = CLBLM_L_X74Y126_SLICE_X112Y126_DQ;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_D5 = CLBLM_L_X74Y126_SLICE_X112Y126_CO6;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_D6 = CLBLL_R_X75Y128_SLICE_X114Y128_AO6;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_A2 = CLBLM_R_X63Y97_SLICE_X95Y97_DO6;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_A3 = CLBLM_R_X63Y98_SLICE_X94Y98_CO6;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_A4 = CLBLM_R_X63Y98_SLICE_X95Y98_BO6;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_A5 = CLBLM_L_X64Y103_SLICE_X97Y103_CO6;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_A6 = CLBLM_R_X63Y98_SLICE_X95Y98_CO6;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_B1 = CLBLM_R_X63Y99_SLICE_X95Y99_DO6;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_B2 = CLBLM_R_X63Y98_SLICE_X94Y98_BO6;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_B3 = CLBLM_R_X63Y99_SLICE_X95Y99_AO6;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_B4 = CLBLM_L_X64Y98_SLICE_X96Y98_CO6;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_B5 = CLBLM_R_X63Y97_SLICE_X94Y97_AO6;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_B6 = CLBLM_L_X64Y99_SLICE_X96Y99_CQ;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_C3 = CLBLM_R_X63Y97_SLICE_X95Y97_CO6;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_C4 = CLBLM_L_X64Y97_SLICE_X97Y97_A5Q;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_C5 = CLBLM_R_X63Y96_SLICE_X95Y96_DQ;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_C6 = CLBLM_R_X63Y99_SLICE_X95Y99_BQ;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_C1 = CLBLM_R_X63Y97_SLICE_X94Y97_AQ;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_C2 = CLBLM_R_X63Y99_SLICE_X95Y99_B5Q;
  assign CLBLM_R_X67Y110_SLICE_X100Y110_A1 = CLBLM_R_X67Y111_SLICE_X101Y111_DO6;
  assign CLBLM_R_X67Y110_SLICE_X100Y110_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y110_SLICE_X100Y110_A3 = CLBLM_R_X67Y110_SLICE_X100Y110_AQ;
  assign CLBLM_R_X67Y110_SLICE_X100Y110_A4 = CLBLM_R_X67Y110_SLICE_X101Y110_BQ;
  assign CLBLM_R_X67Y110_SLICE_X100Y110_A5 = CLBLM_R_X65Y110_SLICE_X99Y110_AO6;
  assign CLBLM_L_X76Y118_SLICE_X116Y118_D3 = 1'b1;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_D1 = 1'b1;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_D2 = 1'b1;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_D3 = 1'b1;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_D4 = 1'b1;
  assign CLBLM_L_X76Y118_SLICE_X116Y118_D4 = 1'b1;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_D5 = 1'b1;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_D6 = 1'b1;
  assign CLBLM_L_X76Y118_SLICE_X116Y118_D5 = 1'b1;
  assign CLBLM_R_X67Y110_SLICE_X100Y110_B2 = CLBLM_R_X67Y110_SLICE_X100Y110_BQ;
  assign CLBLM_R_X67Y110_SLICE_X100Y110_B3 = CLBLM_R_X67Y110_SLICE_X100Y110_AQ;
  assign CLBLM_R_X67Y110_SLICE_X100Y110_B4 = CLBLM_R_X67Y111_SLICE_X101Y111_DO5;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_A1 = CLBLM_L_X62Y99_SLICE_X93Y99_AQ;
  assign CLBLM_L_X76Y118_SLICE_X116Y118_D6 = 1'b1;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_A2 = CLBLM_R_X63Y98_SLICE_X94Y98_BQ;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_A3 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_A4 = CLBLM_L_X64Y97_SLICE_X97Y97_A5Q;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_A5 = CLBLM_L_X76Y111_SLICE_X116Y111_BQ;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_A6 = 1'b1;
  assign CLBLM_R_X67Y110_SLICE_X100Y110_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y110_SLICE_X100Y110_C2 = CLBLM_R_X67Y110_SLICE_X100Y110_CQ;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_AX = CLBLM_L_X60Y92_SLICE_X90Y92_BQ;
  assign CLBLM_R_X67Y110_SLICE_X100Y110_C4 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_B1 = CLBLM_L_X62Y99_SLICE_X93Y99_AQ;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_B2 = CLBLM_R_X63Y99_SLICE_X95Y99_BQ;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_B3 = CLBLM_L_X64Y97_SLICE_X97Y97_A5Q;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_B4 = CLBLM_R_X63Y99_SLICE_X95Y99_B5Q;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_B5 = CLBLM_R_X63Y96_SLICE_X94Y96_AQ;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_B6 = 1'b1;
  assign CLBLM_R_X67Y110_SLICE_X100Y110_D1 = CLBLM_L_X68Y108_SLICE_X102Y108_AQ;
  assign CLBLM_R_X67Y110_SLICE_X100Y110_D2 = CLBLM_L_X68Y108_SLICE_X102Y108_A5Q;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_BX = CLBLM_L_X76Y111_SLICE_X116Y111_BQ;
  assign CLBLM_L_X76Y118_SLICE_X116Y118_DX = CLBLM_L_X76Y118_SLICE_X116Y118_AQ;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_C1 = CLBLM_R_X63Y98_SLICE_X94Y98_AO6;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_C2 = CLBLM_R_X63Y97_SLICE_X94Y97_CO6;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_C3 = CLBLM_L_X62Y98_SLICE_X93Y98_BQ;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_C4 = CLBLM_R_X63Y98_SLICE_X94Y98_BQ;
  assign CLBLM_L_X76Y118_SLICE_X116Y118_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_C5 = CLBLM_R_X63Y98_SLICE_X94Y98_BO5;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_C6 = CLBLM_R_X63Y98_SLICE_X94Y98_DO6;
  assign CLBLM_R_X67Y110_SLICE_X100Y110_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign LIOB33_X0Y113_IOB_X0Y113_O = CLBLM_R_X63Y122_SLICE_X95Y122_CQ;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_D1 = CLBLM_L_X76Y111_SLICE_X116Y111_BQ;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_D2 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_D3 = CLBLM_L_X62Y98_SLICE_X93Y98_CQ;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_D4 = CLBLM_R_X63Y99_SLICE_X95Y99_B5Q;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_D5 = CLBLM_L_X62Y98_SLICE_X93Y98_AQ;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_D6 = CLBLM_R_X63Y99_SLICE_X95Y99_BQ;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_A1 = CLBLL_R_X75Y127_SLICE_X114Y127_A5Q;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_A2 = CLBLL_R_X73Y127_SLICE_X111Y127_BO6;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_A3 = CLBLL_R_X73Y127_SLICE_X110Y127_AQ;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_A4 = CLBLL_R_X75Y128_SLICE_X114Y128_BO6;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_A5 = CLBLL_R_X73Y127_SLICE_X110Y127_BQ;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_A6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_AX = CLBLL_R_X73Y127_SLICE_X110Y127_CO5;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_B1 = CLBLL_R_X75Y128_SLICE_X115Y128_CO6;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_B2 = CLBLL_R_X73Y127_SLICE_X110Y127_BQ;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_B3 = CLBLL_R_X73Y127_SLICE_X110Y127_DQ;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_B4 = CLBLL_R_X75Y128_SLICE_X114Y128_BO6;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_B6 = CLBLL_R_X73Y127_SLICE_X110Y127_CO6;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_D1 = RIOB33_X105Y53_IOB_X1Y53_I;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_C2 = CLBLL_R_X75Y128_SLICE_X115Y128_CO6;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_C3 = CLBLL_R_X75Y127_SLICE_X114Y127_AQ;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_C4 = CLBLL_R_X73Y127_SLICE_X110Y127_A5Q;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_C5 = CLBLM_L_X72Y127_SLICE_X109Y127_AQ;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_C6 = 1'b1;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_D1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_D2 = CLBLL_R_X75Y127_SLICE_X114Y127_BQ;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_D3 = CLBLL_R_X73Y127_SLICE_X110Y127_DQ;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_D4 = CLBLL_R_X75Y128_SLICE_X114Y128_BO6;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_D5 = CLBLL_R_X75Y128_SLICE_X115Y128_CO6;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_D6 = CLBLL_R_X75Y127_SLICE_X114Y127_CO5;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_A1 = CLBLL_R_X73Y127_SLICE_X110Y127_A5Q;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_A2 = CLBLL_R_X75Y128_SLICE_X114Y128_BO6;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_A3 = CLBLL_R_X73Y127_SLICE_X111Y127_AQ;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_A4 = CLBLL_R_X73Y127_SLICE_X111Y127_BO6;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_A5 = CLBLL_R_X73Y127_SLICE_X111Y127_CQ;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_A6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_B1 = CLBLL_R_X75Y127_SLICE_X114Y127_A5Q;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_B2 = CLBLL_R_X75Y128_SLICE_X115Y128_CO6;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_B3 = 1'b1;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_B4 = 1'b1;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_B5 = CLBLL_R_X75Y127_SLICE_X114Y127_AQ;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_B6 = 1'b1;
  assign CLBLM_R_X67Y111_SLICE_X101Y111_A1 = CLBLM_R_X67Y111_SLICE_X101Y111_AQ;
  assign CLBLM_R_X67Y111_SLICE_X101Y111_A2 = CLBLM_R_X67Y111_SLICE_X101Y111_A5Q;
  assign CLBLM_R_X67Y111_SLICE_X101Y111_A3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_C2 = CLBLL_R_X73Y127_SLICE_X111Y127_CQ;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_C3 = CLBLL_R_X75Y127_SLICE_X114Y127_DQ;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_C4 = CLBLL_R_X75Y128_SLICE_X114Y128_BO6;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_C5 = CLBLL_R_X73Y127_SLICE_X111Y127_BO5;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_C6 = 1'b1;
  assign CLBLM_R_X67Y111_SLICE_X101Y111_A4 = CLBLM_R_X67Y111_SLICE_X101Y111_B5Q;
  assign CLBLM_R_X67Y111_SLICE_X101Y111_A5 = 1'b1;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X67Y111_SLICE_X101Y111_A6 = 1'b1;
  assign CLBLM_R_X67Y111_SLICE_X101Y111_B1 = CLBLM_R_X67Y111_SLICE_X101Y111_AQ;
  assign CLBLM_R_X67Y111_SLICE_X101Y111_B2 = CLBLM_R_X67Y111_SLICE_X101Y111_BQ;
  assign CLBLM_R_X67Y111_SLICE_X101Y111_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_D1 = 1'b1;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_D2 = 1'b1;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_D3 = 1'b1;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_D4 = 1'b1;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_D5 = 1'b1;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_D6 = 1'b1;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_A1 = CLBLM_R_X63Y99_SLICE_X95Y99_B5Q;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_A2 = CLBLM_R_X63Y99_SLICE_X95Y99_BQ;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_A3 = CLBLM_L_X60Y92_SLICE_X90Y92_BQ;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_A4 = CLBLM_L_X64Y103_SLICE_X97Y103_CO6;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_A5 = CLBLM_L_X64Y97_SLICE_X97Y97_A5Q;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_A6 = 1'b1;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_B1 = CLBLM_R_X63Y99_SLICE_X95Y99_B5Q;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_B2 = CLBLM_R_X63Y99_SLICE_X95Y99_BQ;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_B4 = CLBLM_L_X64Y103_SLICE_X97Y103_CO6;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_B5 = CLBLM_R_X63Y99_SLICE_X94Y99_D5Q;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_B6 = 1'b1;
  assign CLBLM_R_X67Y111_SLICE_X101Y111_D1 = 1'b1;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_C1 = CLBLM_R_X63Y99_SLICE_X94Y99_D5Q;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_C2 = CLBLM_L_X64Y103_SLICE_X97Y103_CO6;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_C3 = CLBLM_L_X64Y102_SLICE_X97Y102_AQ;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_C4 = CLBLM_R_X63Y99_SLICE_X95Y99_BQ;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_C5 = CLBLM_R_X63Y99_SLICE_X94Y99_DQ;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_C6 = CLBLM_R_X63Y99_SLICE_X95Y99_B5Q;
  assign CLBLM_R_X67Y111_SLICE_X100Y111_A1 = CLBLM_R_X67Y111_SLICE_X101Y111_B5Q;
  assign CLBLM_R_X67Y111_SLICE_X100Y111_A2 = CLBLM_R_X67Y111_SLICE_X100Y111_BQ;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X67Y111_SLICE_X100Y111_A3 = CLBLM_R_X67Y111_SLICE_X100Y111_AQ;
  assign CLBLM_R_X67Y111_SLICE_X100Y111_A4 = CLBLM_R_X67Y111_SLICE_X101Y111_A5Q;
  assign CLBLM_R_X67Y111_SLICE_X100Y111_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y111_SLICE_X100Y111_A6 = CLBLM_R_X67Y111_SLICE_X100Y111_A5Q;
  assign CLBLM_R_X67Y111_SLICE_X100Y111_AX = CLBLM_R_X67Y111_SLICE_X100Y111_CO6;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_D1 = 1'b1;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_D2 = 1'b1;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_D3 = 1'b1;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_D4 = CLBLM_R_X63Y99_SLICE_X95Y99_BQ;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_D5 = CLBLM_R_X63Y99_SLICE_X95Y99_B5Q;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_D6 = 1'b1;
  assign CLBLM_R_X67Y111_SLICE_X100Y111_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y111_SLICE_X100Y111_B2 = CLBLM_R_X67Y111_SLICE_X100Y111_BQ;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X67Y111_SLICE_X100Y111_B3 = CLBLM_R_X67Y111_SLICE_X101Y111_B5Q;
  assign CLBLM_R_X67Y111_SLICE_X100Y111_B4 = CLBLM_R_X67Y111_SLICE_X101Y111_A5Q;
  assign CLBLM_R_X67Y111_SLICE_X100Y111_B5 = CLBLL_R_X79Y99_SLICE_X122Y99_AO6;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_A1 = 1'b1;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_A2 = CLBLM_R_X63Y99_SLICE_X94Y99_A5Q;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_A3 = CLBLM_R_X63Y99_SLICE_X94Y99_AQ;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_A4 = CLBLM_L_X64Y99_SLICE_X96Y99_AQ;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_A6 = 1'b1;
  assign CLBLM_R_X67Y111_SLICE_X100Y111_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y111_SLICE_X100Y111_C2 = CLBLM_R_X67Y111_SLICE_X101Y111_A5Q;
  assign CLBLM_R_X67Y111_SLICE_X100Y111_C3 = CLBLM_R_X67Y111_SLICE_X101Y111_B5Q;
  assign CLBLM_R_X67Y111_SLICE_X100Y111_C4 = CLBLM_R_X67Y111_SLICE_X100Y111_A5Q;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_B1 = 1'b1;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_B2 = CLBLM_R_X63Y99_SLICE_X94Y99_A5Q;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_B3 = CLBLM_R_X63Y99_SLICE_X94Y99_AQ;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_B4 = 1'b1;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_B5 = CLBLM_L_X64Y99_SLICE_X96Y99_AQ;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_B6 = 1'b1;
  assign CLBLM_R_X67Y111_SLICE_X100Y111_D1 = 1'b1;
  assign CLBLM_R_X67Y111_SLICE_X100Y111_D2 = 1'b1;
  assign CLBLM_R_X67Y111_SLICE_X100Y111_D3 = 1'b1;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_C1 = CLBLM_L_X64Y99_SLICE_X96Y99_AQ;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_C2 = CLBLM_R_X63Y99_SLICE_X94Y99_AQ;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_C3 = 1'b1;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_C4 = 1'b1;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_C5 = 1'b1;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_C6 = 1'b1;
  assign CLBLM_R_X67Y111_SLICE_X100Y111_D6 = 1'b1;
  assign CLBLM_R_X67Y111_SLICE_X100Y111_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_D1 = CLBLM_R_X63Y98_SLICE_X94Y98_AO5;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_D2 = CLBLM_R_X63Y99_SLICE_X94Y99_D5Q;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_D3 = CLBLM_R_X63Y99_SLICE_X94Y99_DQ;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_D4 = CLBLM_L_X64Y97_SLICE_X97Y97_A5Q;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_D5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_D6 = 1'b1;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_A2 = CLBLL_R_X75Y127_SLICE_X114Y127_A5Q;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_A3 = CLBLL_R_X73Y128_SLICE_X110Y128_AQ;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_A4 = CLBLL_R_X73Y128_SLICE_X111Y128_BQ;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_A5 = CLBLL_R_X75Y127_SLICE_X114Y127_AQ;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_A6 = CLBLL_R_X75Y128_SLICE_X115Y128_CO6;
  assign LIOB33_X0Y147_IOB_X0Y148_O = CLBLL_R_X73Y134_SLICE_X110Y134_AO5;
  assign LIOI3_X0Y77_OLOGIC_X0Y78_D1 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_B1 = 1'b1;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_B2 = 1'b1;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_B3 = 1'b1;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_B4 = 1'b1;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_B5 = 1'b1;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_B6 = 1'b1;
  assign LIOI3_X0Y77_OLOGIC_X0Y78_T1 = 1'b1;
  assign RIOI3_X105Y123_OLOGIC_X1Y124_D1 = CLBLM_L_X68Y99_SLICE_X102Y99_AQ;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_C1 = 1'b1;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_C2 = 1'b1;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_C3 = 1'b1;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_C4 = 1'b1;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_C5 = 1'b1;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_C6 = 1'b1;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOB33_X0Y147_IOB_X0Y147_O = CLBLL_R_X71Y124_SLICE_X106Y124_BO6;
  assign LIOI3_X0Y77_OLOGIC_X0Y77_D1 = CLBLM_L_X60Y97_SLICE_X90Y97_BQ;
  assign RIOI3_X105Y123_OLOGIC_X1Y124_T1 = 1'b1;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_D1 = 1'b1;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_D2 = 1'b1;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_D3 = 1'b1;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_D4 = 1'b1;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_D5 = 1'b1;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_D6 = 1'b1;
  assign LIOI3_X0Y77_OLOGIC_X0Y77_T1 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_D4 = 1'b1;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1 = CLBLM_L_X70Y126_SLICE_X104Y126_DO6;
  assign RIOI3_X105Y123_OLOGIC_X1Y123_D1 = CLBLM_R_X63Y101_SLICE_X94Y101_AQ;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_D5 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_D6 = 1'b1;
  assign RIOI3_X105Y123_OLOGIC_X1Y123_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1 = CLBLM_L_X64Y106_SLICE_X97Y106_AO6;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_A1 = CLBLL_R_X73Y126_SLICE_X110Y126_DQ;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_A3 = CLBLL_R_X73Y128_SLICE_X111Y128_AQ;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_A4 = CLBLL_R_X75Y127_SLICE_X114Y127_A5Q;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_A5 = CLBLL_R_X75Y127_SLICE_X114Y127_AQ;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_A6 = CLBLL_R_X75Y128_SLICE_X115Y128_CO6;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1 = 1'b1;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_B1 = CLBLL_R_X73Y127_SLICE_X111Y127_BO5;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_B2 = CLBLL_R_X73Y128_SLICE_X111Y128_BQ;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_B3 = CLBLL_R_X73Y128_SLICE_X111Y128_AQ;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_B4 = 1'b1;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_B6 = CLBLL_R_X73Y126_SLICE_X110Y126_DQ;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_C1 = 1'b1;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_C2 = 1'b1;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_C3 = 1'b1;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_C4 = 1'b1;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_C5 = 1'b1;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_C6 = 1'b1;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_D1 = 1'b1;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_D2 = 1'b1;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_D3 = 1'b1;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_D4 = 1'b1;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_D5 = 1'b1;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_D6 = 1'b1;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign LIOB33_X0Y117_IOB_X0Y118_O = CLBLM_R_X67Y116_SLICE_X100Y116_AQ;
  assign LIOB33_X0Y117_IOB_X0Y117_O = CLBLM_L_X76Y125_SLICE_X116Y125_AQ;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_B6 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_BX = CLBLM_L_X72Y117_SLICE_X108Y117_AQ;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_C1 = CLBLM_L_X72Y130_SLICE_X108Y130_AQ;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_C3 = 1'b1;
  assign CLBLM_R_X67Y108_SLICE_X100Y108_A4 = CLBLM_R_X67Y108_SLICE_X100Y108_AQ;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_C2 = CLBLM_L_X72Y131_SLICE_X108Y131_CQ;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_C5 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_C6 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_CE = CLBLM_L_X76Y109_SLICE_X116Y109_AO6;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_C3 = CLBLM_L_X72Y131_SLICE_X108Y131_BQ;
  assign CLBLM_L_X68Y107_SLICE_X103Y107_D4 = CLBLM_L_X68Y109_SLICE_X103Y109_B5Q;
  assign CLBLM_L_X68Y107_SLICE_X103Y107_D5 = CLBLM_L_X68Y106_SLICE_X103Y106_BQ;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_C4 = CLBLM_L_X72Y134_SLICE_X109Y134_AO5;
  assign CLBLM_L_X68Y107_SLICE_X103Y107_D6 = CLBLM_L_X68Y109_SLICE_X103Y109_BQ;
  assign CLBLM_L_X76Y109_SLICE_X117Y109_A1 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X117Y109_A2 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X117Y109_A3 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X117Y109_A4 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X117Y109_A5 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X117Y109_A6 = 1'b1;
  assign LIOB33_X0Y169_IOB_X0Y170_O = CLBLM_L_X74Y120_SLICE_X112Y120_AO6;
  assign CLBLM_L_X76Y109_SLICE_X117Y109_B1 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X117Y109_B2 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X117Y109_B3 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X117Y109_B4 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X117Y109_B5 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X117Y109_B6 = 1'b1;
  assign LIOB33_X0Y169_IOB_X0Y169_O = CLBLL_R_X73Y131_SLICE_X110Y131_AQ;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_D4 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X117Y109_C1 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X117Y109_C2 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X117Y109_C3 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X117Y109_C4 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_D5 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X117Y109_C5 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X117Y109_C6 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X117Y109_D1 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X117Y109_D2 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X117Y109_D3 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X117Y109_D4 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X117Y109_D5 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X117Y109_D6 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_C6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign RIOB33_X105Y151_IOB_X1Y151_O = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X116Y109_A1 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X116Y109_A2 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X116Y109_A3 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X116Y109_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X76Y109_SLICE_X116Y109_A5 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X116Y109_A6 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X116Y109_B1 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X116Y109_B2 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X116Y109_B3 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X116Y109_B4 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X116Y109_B5 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X116Y109_B6 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X116Y109_C1 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X116Y109_C2 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X116Y109_C3 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X116Y109_C4 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X116Y109_C5 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X116Y109_C6 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X116Y109_D1 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X116Y109_D2 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X116Y109_D3 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X116Y109_D4 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X116Y109_D5 = 1'b1;
  assign CLBLM_L_X76Y109_SLICE_X116Y109_D6 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_D1 = 1'b1;
  assign LIOB33_X0Y119_IOB_X0Y120_O = CLBLL_R_X71Y119_SLICE_X106Y119_AQ;
  assign LIOB33_X0Y119_IOB_X0Y119_O = CLBLM_R_X63Y106_SLICE_X95Y106_AQ;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_A1 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_A2 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_A3 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_A4 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_A5 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_A6 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_B1 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_B2 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_B3 = 1'b1;
  assign CLBLM_L_X68Y107_SLICE_X102Y107_C5 = CLBLM_L_X68Y107_SLICE_X102Y107_DO6;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_B4 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_B5 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_B6 = 1'b1;
  assign CLBLM_L_X68Y107_SLICE_X102Y107_C6 = CLBLM_L_X72Y105_SLICE_X108Y105_CQ;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_C1 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_C2 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_C3 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_C4 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_C5 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_C6 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_T1 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_D1 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_D2 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_D3 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_D4 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_D5 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_D6 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_A1 = CLBLM_R_X63Y102_SLICE_X95Y102_DQ;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_A2 = CLBLM_L_X64Y101_SLICE_X96Y101_B5Q;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_A3 = CLBLM_L_X64Y101_SLICE_X96Y101_BQ;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_A4 = CLBLM_L_X64Y101_SLICE_X96Y101_A5Q;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_A5 = CLBLM_L_X60Y99_SLICE_X90Y99_CQ;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_A6 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_AX = CLBLM_L_X60Y99_SLICE_X90Y99_CQ;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_B1 = CLBLM_L_X64Y101_SLICE_X96Y101_B5Q;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_B2 = CLBLM_L_X64Y103_SLICE_X97Y103_DO6;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_B3 = CLBLM_L_X60Y99_SLICE_X90Y99_CQ;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_B4 = CLBLM_L_X64Y101_SLICE_X96Y101_A5Q;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_B5 = CLBLM_L_X64Y101_SLICE_X96Y101_BQ;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_B6 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_BX = CLBLM_R_X63Y103_SLICE_X94Y103_AQ;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_C1 = CLBLM_R_X63Y101_SLICE_X94Y101_BQ;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_C2 = CLBLM_R_X63Y101_SLICE_X94Y101_AQ;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_C3 = CLBLM_R_X63Y102_SLICE_X95Y102_BQ;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_C4 = CLBLM_L_X64Y101_SLICE_X96Y101_BQ;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_C5 = CLBLM_L_X64Y101_SLICE_X96Y101_B5Q;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_C6 = CLBLM_R_X63Y102_SLICE_X94Y102_AQ;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_D1 = CLBLM_L_X62Y101_SLICE_X93Y101_DO6;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_D2 = CLBLM_R_X63Y103_SLICE_X94Y103_CO6;
  assign CLBLM_L_X68Y107_SLICE_X102Y107_D4 = CLBLM_R_X65Y106_SLICE_X98Y106_CQ;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_D3 = CLBLM_L_X62Y101_SLICE_X93Y101_CO6;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_D4 = CLBLM_R_X63Y101_SLICE_X94Y101_AO5;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_D5 = CLBLM_R_X63Y103_SLICE_X94Y103_DO6;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_D6 = CLBLM_L_X64Y103_SLICE_X97Y103_DO6;
  assign CLBLM_L_X68Y107_SLICE_X102Y107_D5 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y102_SLICE_X113Y102_A1 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X113Y102_A2 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X113Y102_A3 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X113Y102_A4 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X113Y102_A5 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X113Y102_A6 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X113Y102_B1 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X113Y102_B2 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X113Y102_B3 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X113Y102_B4 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X113Y102_B5 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X113Y102_B6 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X113Y102_C1 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X113Y102_C2 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X113Y102_C3 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X113Y102_C4 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X113Y102_C5 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X113Y102_C6 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X113Y102_D1 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X113Y102_D2 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X113Y102_D3 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X113Y102_D4 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X113Y102_D5 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X113Y102_D6 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X112Y102_A1 = CLBLM_L_X72Y103_SLICE_X108Y103_DO5;
  assign CLBLM_L_X74Y102_SLICE_X112Y102_A2 = CLBLM_L_X72Y103_SLICE_X108Y103_CO6;
  assign CLBLM_L_X74Y102_SLICE_X112Y102_A3 = CLBLM_L_X74Y102_SLICE_X112Y102_AQ;
  assign CLBLM_L_X74Y102_SLICE_X112Y102_A4 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X74Y102_SLICE_X112Y102_A5 = CLBLL_R_X73Y101_SLICE_X110Y101_AQ;
  assign CLBLM_L_X74Y102_SLICE_X112Y102_A6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y102_SLICE_X112Y102_B1 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X112Y102_B2 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X112Y102_B3 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X112Y102_B4 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X112Y102_B5 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X112Y102_B6 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X112Y102_C1 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X112Y102_C2 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X112Y102_C3 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X112Y102_C4 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X112Y102_C5 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X112Y102_C6 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X112Y102_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOB33_X0Y121_IOB_X0Y122_O = RIOB33_X105Y51_IOB_X1Y52_I;
  assign LIOB33_X0Y121_IOB_X0Y121_O = CLBLL_R_X73Y123_SLICE_X110Y123_AQ;
  assign CLBLM_L_X74Y102_SLICE_X112Y102_D1 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X112Y102_D2 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X112Y102_D3 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X112Y102_D4 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X112Y102_D5 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X112Y102_D6 = 1'b1;
  assign CLBLM_L_X74Y102_SLICE_X112Y102_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_A1 = CLBLM_L_X64Y102_SLICE_X96Y102_A5Q;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_D6 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_A3 = CLBLM_R_X63Y102_SLICE_X95Y102_AQ;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_A4 = CLBLM_L_X64Y102_SLICE_X96Y102_AQ;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_A5 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_A6 = 1'b1;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_D1 = CLBLM_L_X60Y92_SLICE_X90Y92_BQ;
  assign LIOI3_TBYTESRC_X0Y81_OLOGIC_X0Y82_D1 = CLBLM_L_X62Y107_SLICE_X93Y107_A5Q;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_B1 = CLBLM_L_X64Y102_SLICE_X96Y102_A5Q;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_B2 = CLBLM_R_X63Y102_SLICE_X95Y102_BQ;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_B3 = CLBLM_L_X64Y102_SLICE_X96Y102_BO5;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_B4 = CLBLM_R_X63Y102_SLICE_X95Y102_CQ;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_B5 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_B6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_T1 = 1'b1;
  assign RIOI3_X105Y125_OLOGIC_X1Y126_D1 = CLBLM_L_X76Y127_SLICE_X116Y127_AQ;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_C1 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_C2 = CLBLM_L_X64Y102_SLICE_X96Y102_CQ;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_C3 = CLBLM_R_X63Y103_SLICE_X94Y103_AO5;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_C4 = CLBLM_L_X64Y102_SLICE_X96Y102_BO5;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_C5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_C6 = CLBLM_R_X63Y102_SLICE_X95Y102_CQ;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_X0Y79_OLOGIC_X0Y79_D1 = CLBLM_L_X64Y106_SLICE_X96Y106_A5Q;
  assign RIOI3_X105Y125_OLOGIC_X1Y126_T1 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_D1 = CLBLM_L_X62Y102_SLICE_X92Y102_CQ;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_D2 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_D3 = CLBLM_R_X63Y102_SLICE_X95Y102_DQ;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_D4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_D5 = CLBLM_R_X63Y103_SLICE_X95Y103_BO5;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_D6 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign LIOI3_X0Y79_OLOGIC_X0Y79_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign RIOI3_X105Y125_OLOGIC_X1Y125_D1 = CLBLM_L_X74Y129_SLICE_X112Y129_BQ;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_A1 = CLBLM_L_X62Y102_SLICE_X93Y102_AQ;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_A2 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_A3 = CLBLM_R_X63Y102_SLICE_X94Y102_AQ;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_A4 = CLBLM_R_X63Y102_SLICE_X95Y102_AO5;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_A5 = CLBLM_L_X64Y102_SLICE_X96Y102_BO5;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_A6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1 = 1'b1;
  assign RIOI3_X105Y125_OLOGIC_X1Y125_T1 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_B1 = CLBLM_L_X64Y102_SLICE_X96Y102_BO5;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_B2 = CLBLM_R_X63Y102_SLICE_X94Y102_BQ;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_B3 = CLBLM_R_X63Y102_SLICE_X94Y102_AQ;
  assign CLBLM_L_X74Y133_SLICE_X113Y133_A4 = CLBLM_L_X74Y135_SLICE_X113Y135_BQ;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_B4 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_B6 = CLBLM_R_X63Y103_SLICE_X94Y103_AO6;
  assign LIOI3_TBYTESRC_X0Y81_OLOGIC_X0Y82_T1 = 1'b1;
  assign CLBLM_L_X74Y133_SLICE_X113Y133_A5 = CLBLM_L_X74Y133_SLICE_X112Y133_CQ;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_C1 = CLBLM_R_X63Y102_SLICE_X95Y102_CQ;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_C2 = CLBLM_L_X64Y101_SLICE_X96Y101_BQ;
  assign CLBLM_L_X74Y133_SLICE_X113Y133_A6 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_C3 = CLBLM_L_X64Y101_SLICE_X96Y101_B5Q;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_C4 = CLBLM_R_X63Y103_SLICE_X94Y103_AQ;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_C5 = CLBLM_L_X62Y102_SLICE_X93Y102_AQ;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_C6 = CLBLM_L_X60Y99_SLICE_X90Y99_CQ;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_D1 = CLBLM_R_X63Y102_SLICE_X95Y102_AQ;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_D2 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_D3 = CLBLM_L_X64Y105_SLICE_X96Y105_C5Q;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_D4 = CLBLM_L_X64Y105_SLICE_X96Y105_CQ;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_D5 = CLBLM_L_X64Y102_SLICE_X96Y102_AQ;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_D6 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y133_SLICE_X113Y133_B1 = 1'b1;
  assign CLBLM_L_X76Y119_SLICE_X117Y119_D5 = 1'b1;
  assign CLBLM_L_X76Y119_SLICE_X117Y119_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y81_OLOGIC_X0Y81_D1 = CLBLM_L_X60Y99_SLICE_X90Y99_BQ;
  assign CLBLL_R_X73Y109_SLICE_X110Y109_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y109_SLICE_X110Y109_A6 = CLBLM_L_X72Y109_SLICE_X109Y109_B5Q;
  assign CLBLM_L_X76Y111_SLICE_X117Y111_A1 = 1'b1;
  assign CLBLM_L_X76Y111_SLICE_X117Y111_A2 = 1'b1;
  assign CLBLM_L_X76Y111_SLICE_X117Y111_A3 = 1'b1;
  assign CLBLM_L_X76Y111_SLICE_X117Y111_A4 = 1'b1;
  assign CLBLM_L_X76Y111_SLICE_X117Y111_A5 = 1'b1;
  assign CLBLM_L_X76Y111_SLICE_X117Y111_A6 = 1'b1;
  assign CLBLM_L_X76Y119_SLICE_X116Y119_A4 = CLBLL_R_X77Y127_SLICE_X118Y127_AQ;
  assign CLBLM_L_X76Y111_SLICE_X117Y111_B1 = 1'b1;
  assign CLBLM_L_X76Y111_SLICE_X117Y111_B2 = 1'b1;
  assign CLBLM_L_X76Y111_SLICE_X117Y111_B3 = 1'b1;
  assign CLBLM_L_X76Y111_SLICE_X117Y111_B4 = 1'b1;
  assign CLBLM_L_X76Y111_SLICE_X117Y111_B5 = 1'b1;
  assign CLBLM_L_X76Y111_SLICE_X117Y111_B6 = 1'b1;
  assign CLBLM_L_X74Y103_SLICE_X113Y103_A1 = CLBLM_L_X72Y103_SLICE_X108Y103_BO5;
  assign CLBLM_L_X74Y103_SLICE_X113Y103_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y103_SLICE_X113Y103_A3 = CLBLM_L_X74Y103_SLICE_X113Y103_AQ;
  assign CLBLM_L_X74Y103_SLICE_X113Y103_A4 = CLBLL_R_X73Y104_SLICE_X110Y104_DO6;
  assign CLBLM_L_X74Y103_SLICE_X113Y103_A5 = CLBLM_L_X74Y103_SLICE_X112Y103_AQ;
  assign CLBLL_R_X73Y131_SLICE_X110Y131_A1 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X110Y131_A2 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X110Y131_A3 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X110Y131_A4 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X110Y131_A5 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X110Y131_A6 = 1'b1;
  assign CLBLM_L_X74Y103_SLICE_X113Y103_A6 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLL_R_X73Y131_SLICE_X110Y131_AX = CLBLM_L_X70Y136_SLICE_X105Y136_A5Q;
  assign CLBLM_L_X74Y103_SLICE_X113Y103_B1 = CLBLL_R_X73Y104_SLICE_X110Y104_DO6;
  assign CLBLL_R_X73Y131_SLICE_X110Y131_B1 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X110Y131_B2 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X110Y131_B3 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X110Y131_B4 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X110Y131_B5 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X110Y131_B6 = 1'b1;
  assign CLBLM_L_X74Y103_SLICE_X113Y103_B3 = CLBLM_L_X74Y103_SLICE_X113Y103_AQ;
  assign CLBLM_L_X74Y103_SLICE_X113Y103_B4 = CLBLM_L_X72Y103_SLICE_X108Y103_DO6;
  assign CLBLM_L_X74Y103_SLICE_X113Y103_B6 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLL_R_X73Y131_SLICE_X110Y131_C1 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X110Y131_C2 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X110Y131_C3 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X110Y131_C4 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X110Y131_C5 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X110Y131_C6 = 1'b1;
  assign CLBLM_L_X74Y103_SLICE_X113Y103_C3 = CLBLL_R_X73Y104_SLICE_X110Y104_A5Q;
  assign CLBLM_L_X74Y103_SLICE_X113Y103_C4 = CLBLM_L_X62Y95_SLICE_X92Y95_AQ;
  assign CLBLL_R_X73Y131_SLICE_X110Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y103_SLICE_X113Y103_C6 = CLBLM_L_X72Y104_SLICE_X109Y104_BQ;
  assign CLBLM_L_X74Y103_SLICE_X113Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y103_SLICE_X113Y103_D1 = 1'b1;
  assign CLBLM_L_X74Y103_SLICE_X113Y103_D2 = CLBLM_L_X72Y104_SLICE_X109Y104_B5Q;
  assign CLBLL_R_X73Y131_SLICE_X110Y131_D1 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X110Y131_D2 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X110Y131_D3 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X110Y131_D4 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X110Y131_D5 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X110Y131_D6 = 1'b1;
  assign CLBLL_R_X77Y121_SLICE_X119Y121_B3 = CLBLL_R_X77Y121_SLICE_X119Y121_AQ;
  assign CLBLM_L_X74Y103_SLICE_X113Y103_D4 = CLBLM_L_X74Y103_SLICE_X113Y103_CO6;
  assign CLBLL_R_X73Y131_SLICE_X110Y131_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X77Y121_SLICE_X119Y121_B4 = CLBLL_R_X77Y122_SLICE_X119Y122_CQ;
  assign CLBLM_L_X74Y103_SLICE_X112Y103_A1 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X74Y103_SLICE_X112Y103_A2 = CLBLM_L_X72Y103_SLICE_X108Y103_BO6;
  assign CLBLM_L_X74Y103_SLICE_X112Y103_A3 = CLBLM_L_X74Y103_SLICE_X112Y103_AQ;
  assign CLBLL_R_X73Y109_SLICE_X110Y109_C1 = 1'b1;
  assign CLBLL_R_X77Y121_SLICE_X119Y121_B5 = CLBLM_L_X76Y122_SLICE_X117Y122_AQ;
  assign CLBLM_L_X74Y103_SLICE_X112Y103_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y103_SLICE_X112Y103_A5 = CLBLL_R_X73Y102_SLICE_X111Y102_AQ;
  assign CLBLM_L_X74Y103_SLICE_X112Y103_A6 = CLBLL_R_X73Y104_SLICE_X110Y104_DO6;
  assign CLBLL_R_X73Y109_SLICE_X110Y109_C2 = 1'b1;
  assign CLBLL_R_X77Y121_SLICE_X119Y121_B6 = 1'b1;
  assign CLBLM_L_X74Y103_SLICE_X112Y103_B1 = CLBLL_R_X73Y104_SLICE_X110Y104_DO6;
  assign CLBLL_R_X77Y104_SLICE_X118Y104_A1 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X110Y109_C3 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X118Y104_A2 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X118Y104_A3 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X118Y104_A4 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X118Y104_A5 = 1'b1;
  assign CLBLL_R_X73Y109_SLICE_X110Y109_C4 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X118Y104_A6 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X118Y104_AX = CLBLL_R_X77Y104_SLICE_X118Y104_BQ;
  assign CLBLM_L_X74Y103_SLICE_X112Y103_B5 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLL_R_X77Y104_SLICE_X118Y104_B1 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X118Y104_B2 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X111Y131_A1 = CLBLM_L_X70Y136_SLICE_X105Y136_A5Q;
  assign CLBLL_R_X73Y131_SLICE_X111Y131_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y104_SLICE_X118Y104_B5 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X111Y131_A3 = CLBLL_R_X73Y131_SLICE_X111Y131_AQ;
  assign CLBLL_R_X77Y104_SLICE_X118Y104_B6 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X111Y131_A4 = CLBLM_L_X60Y94_SLICE_X90Y94_AQ;
  assign CLBLL_R_X73Y131_SLICE_X111Y131_A5 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X118Y104_BX = CLBLL_R_X77Y104_SLICE_X118Y104_CQ;
  assign CLBLL_R_X77Y104_SLICE_X118Y104_C1 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X118Y104_C2 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X118Y104_C3 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X111Y131_A6 = CLBLM_L_X74Y132_SLICE_X112Y132_CQ;
  assign CLBLL_R_X83Y94_SLICE_X130Y94_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X83Y94_SLICE_X130Y94_A2 = CLBLL_R_X83Y94_SLICE_X130Y94_BQ;
  assign CLBLL_R_X83Y94_SLICE_X130Y94_A3 = 1'b1;
  assign CLBLL_R_X83Y94_SLICE_X130Y94_A4 = CLBLM_L_X82Y98_SLICE_X128Y98_A5Q;
  assign CLBLL_R_X83Y94_SLICE_X130Y94_A5 = CLBLL_R_X83Y94_SLICE_X130Y94_A5Q;
  assign CLBLL_R_X83Y94_SLICE_X130Y94_A6 = 1'b1;
  assign CLBLL_R_X77Y121_SLICE_X119Y121_C1 = CLBLM_L_X78Y123_SLICE_X121Y123_CO6;
  assign CLBLL_R_X77Y104_SLICE_X118Y104_C4 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X118Y104_CX = CLBLL_R_X77Y104_SLICE_X119Y104_AQ;
  assign CLBLL_R_X83Y94_SLICE_X130Y94_B1 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X118Y104_D1 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X118Y104_D2 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X118Y104_D3 = 1'b1;
  assign CLBLL_R_X83Y94_SLICE_X130Y94_B2 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X118Y104_D5 = 1'b1;
  assign CLBLL_R_X83Y94_SLICE_X130Y94_B3 = 1'b1;
  assign CLBLL_R_X83Y94_SLICE_X130Y94_B4 = 1'b1;
  assign CLBLL_R_X83Y94_SLICE_X130Y94_B5 = 1'b1;
  assign CLBLL_R_X83Y94_SLICE_X130Y94_B6 = 1'b1;
  assign CLBLL_R_X83Y94_SLICE_X130Y94_BX = CLBLL_R_X83Y94_SLICE_X130Y94_A5Q;
  assign CLBLL_R_X83Y94_SLICE_X130Y94_C1 = 1'b1;
  assign CLBLL_R_X83Y94_SLICE_X130Y94_C2 = 1'b1;
  assign CLBLL_R_X83Y94_SLICE_X130Y94_C3 = 1'b1;
  assign CLBLL_R_X83Y94_SLICE_X130Y94_C4 = 1'b1;
  assign CLBLL_R_X83Y94_SLICE_X130Y94_C5 = 1'b1;
  assign CLBLL_R_X83Y94_SLICE_X130Y94_C6 = 1'b1;
  assign CLBLL_R_X77Y121_SLICE_X119Y121_C5 = CLBLM_L_X78Y122_SLICE_X120Y122_DO6;
  assign CLBLL_R_X83Y94_SLICE_X130Y94_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLL_R_X77Y104_SLICE_X118Y104_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X73Y131_SLICE_X111Y131_D1 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X111Y131_D2 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X111Y131_D3 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X111Y131_D4 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X111Y131_D5 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X111Y131_D6 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X111Y131_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X83Y94_SLICE_X130Y94_D1 = 1'b1;
  assign CLBLL_R_X83Y94_SLICE_X130Y94_D2 = 1'b1;
  assign CLBLL_R_X83Y94_SLICE_X130Y94_D3 = 1'b1;
  assign CLBLL_R_X83Y94_SLICE_X130Y94_D4 = 1'b1;
  assign CLBLL_R_X83Y94_SLICE_X130Y94_D5 = 1'b1;
  assign CLBLL_R_X83Y94_SLICE_X130Y94_D6 = 1'b1;
  assign CLBLL_R_X83Y94_SLICE_X130Y94_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X77Y104_SLICE_X119Y104_A1 = CLBLM_L_X64Y106_SLICE_X97Y106_AQ;
  assign CLBLL_R_X77Y104_SLICE_X119Y104_A2 = CLBLL_R_X79Y104_SLICE_X122Y104_BQ;
  assign CLBLL_R_X77Y104_SLICE_X119Y104_A3 = CLBLL_R_X77Y104_SLICE_X119Y104_AQ;
  assign CLBLL_R_X77Y104_SLICE_X119Y104_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y104_SLICE_X119Y104_A5 = CLBLM_L_X78Y104_SLICE_X120Y104_BQ;
  assign CLBLL_R_X77Y104_SLICE_X119Y104_A6 = 1'b1;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_A1 = CLBLM_L_X64Y105_SLICE_X96Y105_C5Q;
  assign CLBLL_R_X77Y104_SLICE_X119Y104_B1 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X119Y104_B2 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X119Y104_B3 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X119Y104_B4 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X119Y104_B5 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X119Y104_B6 = 1'b1;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_B1 = 1'b1;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_B2 = CLBLM_L_X64Y102_SLICE_X96Y102_A5Q;
  assign CLBLL_R_X77Y104_SLICE_X119Y104_C1 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X119Y104_C2 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X119Y104_C3 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X119Y104_C4 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X119Y104_C5 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X119Y104_C6 = 1'b1;
  assign CLBLL_R_X83Y94_SLICE_X131Y94_A1 = 1'b1;
  assign CLBLL_R_X83Y94_SLICE_X131Y94_A2 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X119Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X83Y94_SLICE_X131Y94_A3 = 1'b1;
  assign CLBLL_R_X83Y94_SLICE_X131Y94_A4 = 1'b1;
  assign CLBLL_R_X83Y94_SLICE_X131Y94_A5 = 1'b1;
  assign CLBLL_R_X83Y94_SLICE_X131Y94_A6 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X119Y104_D1 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X119Y104_D2 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X119Y104_D3 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X119Y104_D4 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X119Y104_D5 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X119Y104_D6 = 1'b1;
  assign CLBLL_R_X83Y94_SLICE_X131Y94_B1 = 1'b1;
  assign CLBLL_R_X83Y94_SLICE_X131Y94_B2 = 1'b1;
  assign CLBLL_R_X77Y104_SLICE_X119Y104_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X83Y94_SLICE_X131Y94_B3 = 1'b1;
  assign CLBLL_R_X83Y94_SLICE_X131Y94_B4 = 1'b1;
  assign CLBLL_R_X83Y94_SLICE_X131Y94_B5 = 1'b1;
  assign CLBLL_R_X83Y94_SLICE_X131Y94_B6 = 1'b1;
  assign CLBLL_R_X83Y94_SLICE_X131Y94_C1 = 1'b1;
  assign CLBLL_R_X83Y94_SLICE_X131Y94_C2 = 1'b1;
  assign CLBLL_R_X83Y94_SLICE_X131Y94_C3 = 1'b1;
  assign CLBLL_R_X77Y121_SLICE_X119Y121_D6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X83Y94_SLICE_X131Y94_C4 = 1'b1;
  assign CLBLL_R_X83Y94_SLICE_X131Y94_C5 = 1'b1;
  assign CLBLL_R_X83Y94_SLICE_X131Y94_C6 = 1'b1;
  assign CLBLM_L_X74Y133_SLICE_X112Y133_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X83Y94_SLICE_X131Y94_D1 = 1'b1;
  assign CLBLL_R_X83Y94_SLICE_X131Y94_D2 = 1'b1;
  assign CLBLL_R_X83Y94_SLICE_X131Y94_D3 = 1'b1;
  assign CLBLL_R_X83Y94_SLICE_X131Y94_D4 = 1'b1;
  assign CLBLL_R_X83Y94_SLICE_X131Y94_D5 = 1'b1;
  assign CLBLL_R_X83Y94_SLICE_X131Y94_D6 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_C3 = 1'b1;
  assign CLBLM_L_X76Y119_SLICE_X116Y119_D6 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_C4 = 1'b1;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_B1 = CLBLM_R_X63Y103_SLICE_X95Y103_AQ;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_B2 = CLBLM_L_X64Y101_SLICE_X96Y101_BQ;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_B3 = CLBLM_R_X63Y103_SLICE_X94Y103_AQ;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_B4 = CLBLM_L_X64Y101_SLICE_X96Y101_B5Q;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_B5 = CLBLM_R_X63Y101_SLICE_X94Y101_AQ;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_B6 = CLBLM_L_X62Y103_SLICE_X93Y103_DQ;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_C1 = CLBLM_L_X62Y103_SLICE_X92Y103_B5Q;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_C2 = CLBLM_L_X62Y100_SLICE_X92Y100_AQ;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_C3 = CLBLM_L_X62Y101_SLICE_X92Y101_AQ;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_C4 = CLBLM_L_X62Y103_SLICE_X92Y103_BQ;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_C5 = CLBLM_L_X62Y103_SLICE_X93Y103_CQ;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_C6 = CLBLM_L_X64Y101_SLICE_X96Y101_A5Q;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y133_SLICE_X112Y133_C1 = CLBLM_L_X74Y132_SLICE_X112Y132_AQ;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_D1 = CLBLM_L_X62Y102_SLICE_X92Y102_DO6;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_D2 = CLBLM_R_X63Y103_SLICE_X95Y103_CO6;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_D3 = CLBLM_R_X63Y102_SLICE_X94Y102_CO6;
  assign CLBLM_L_X74Y133_SLICE_X112Y133_C2 = CLBLM_L_X74Y134_SLICE_X113Y134_BQ;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_D4 = CLBLM_R_X63Y101_SLICE_X94Y101_CO6;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_D5 = CLBLM_L_X62Y103_SLICE_X92Y103_CO6;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_D6 = CLBLM_R_X63Y103_SLICE_X94Y103_BO6;
  assign CLBLM_L_X74Y133_SLICE_X112Y133_C3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y133_SLICE_X112Y133_C4 = CLBLM_L_X74Y133_SLICE_X112Y133_BQ;
  assign CLBLM_L_X74Y133_SLICE_X112Y133_C5 = CLBLM_L_X74Y133_SLICE_X112Y133_DO6;
  assign CLBLM_L_X74Y133_SLICE_X112Y133_C6 = CLBLM_L_X74Y133_SLICE_X112Y133_CQ;
  assign CLBLM_L_X80Y132_SLICE_X125Y132_A1 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X125Y132_A2 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X125Y132_A3 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X125Y132_A4 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X125Y132_A5 = 1'b1;
  assign CLBLM_L_X74Y133_SLICE_X112Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X80Y132_SLICE_X125Y132_A6 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X125Y132_B1 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X125Y132_B2 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X125Y132_B3 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X125Y132_B4 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X125Y132_B5 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X125Y132_B6 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X125Y132_C1 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X125Y132_C2 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X125Y132_C3 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X125Y132_C4 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X125Y132_C5 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X125Y132_C6 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_D6 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X125Y132_D1 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X125Y132_D2 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X125Y132_D3 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X125Y132_D4 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X125Y132_D5 = 1'b1;
  assign CLBLM_L_X74Y133_SLICE_X112Y133_D1 = CLBLM_L_X74Y129_SLICE_X112Y129_BQ;
  assign CLBLM_L_X80Y132_SLICE_X125Y132_D6 = 1'b1;
  assign CLBLM_L_X74Y133_SLICE_X112Y133_D2 = CLBLM_L_X74Y134_SLICE_X113Y134_A5Q;
  assign CLBLM_L_X80Y132_SLICE_X124Y132_A1 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X124Y132_A2 = 1'b1;
  assign CLBLM_L_X74Y133_SLICE_X112Y133_D3 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X124Y132_A3 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X124Y132_A4 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X124Y132_A5 = 1'b1;
  assign CLBLM_L_X80Y132_SLICE_X124Y132_A6 = 1'b1;
  assign CLBLM_L_X74Y133_SLICE_X112Y133_D4 = CLBLM_L_X74Y134_SLICE_X113Y134_CQ;
  assign CLBLL_R_X73Y132_SLICE_X110Y132_A1 = CLBLM_L_X74Y132_SLICE_X112Y132_CQ;
  assign CLBLL_R_X73Y132_SLICE_X110Y132_A2 = 1'b1;
  assign CLBLL_R_X73Y132_SLICE_X110Y132_A3 = CLBLM_L_X74Y132_SLICE_X113Y132_BQ;
  assign CLBLL_R_X73Y132_SLICE_X110Y132_A4 = CLBLL_R_X73Y132_SLICE_X111Y132_AO5;
  assign CLBLL_R_X73Y132_SLICE_X110Y132_A5 = CLBLL_R_X73Y131_SLICE_X110Y131_AQ;
  assign CLBLL_R_X73Y132_SLICE_X110Y132_A6 = 1'b1;
  assign CLBLM_L_X74Y104_SLICE_X113Y104_A1 = 1'b1;
  assign CLBLM_L_X74Y104_SLICE_X113Y104_A2 = 1'b1;
  assign CLBLM_L_X74Y104_SLICE_X113Y104_A3 = 1'b1;
  assign CLBLL_R_X73Y132_SLICE_X110Y132_B1 = CLBLL_R_X73Y133_SLICE_X110Y133_A5Q;
  assign CLBLL_R_X73Y132_SLICE_X110Y132_B2 = CLBLM_L_X70Y136_SLICE_X105Y136_CO6;
  assign CLBLL_R_X73Y132_SLICE_X110Y132_B3 = CLBLL_R_X73Y132_SLICE_X111Y132_CO6;
  assign CLBLL_R_X73Y132_SLICE_X110Y132_B4 = CLBLM_L_X74Y134_SLICE_X113Y134_CQ;
  assign CLBLL_R_X73Y132_SLICE_X110Y132_B5 = CLBLM_L_X74Y134_SLICE_X113Y134_A5Q;
  assign CLBLL_R_X73Y132_SLICE_X110Y132_B6 = CLBLL_R_X73Y133_SLICE_X111Y133_A5Q;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_A2 = 1'b1;
  assign CLBLM_L_X74Y104_SLICE_X113Y104_B1 = 1'b1;
  assign CLBLL_R_X73Y132_SLICE_X110Y132_C1 = 1'b1;
  assign CLBLL_R_X73Y132_SLICE_X110Y132_C2 = 1'b1;
  assign CLBLL_R_X73Y132_SLICE_X110Y132_C3 = 1'b1;
  assign CLBLL_R_X73Y132_SLICE_X110Y132_C4 = 1'b1;
  assign CLBLL_R_X73Y132_SLICE_X110Y132_C5 = 1'b1;
  assign CLBLL_R_X73Y132_SLICE_X110Y132_C6 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_A3 = CLBLM_L_X70Y125_SLICE_X104Y125_AQ;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_A4 = CLBLL_R_X71Y126_SLICE_X107Y126_BQ;
  assign CLBLM_L_X74Y104_SLICE_X113Y104_C1 = 1'b1;
  assign CLBLM_L_X74Y104_SLICE_X113Y104_C2 = 1'b1;
  assign CLBLM_L_X74Y104_SLICE_X113Y104_C3 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_A5 = 1'b1;
  assign CLBLM_L_X74Y104_SLICE_X113Y104_C4 = 1'b1;
  assign CLBLM_L_X74Y104_SLICE_X113Y104_C6 = 1'b1;
  assign CLBLL_R_X73Y132_SLICE_X110Y132_D1 = 1'b1;
  assign CLBLL_R_X73Y132_SLICE_X110Y132_D2 = 1'b1;
  assign CLBLL_R_X73Y132_SLICE_X110Y132_D3 = 1'b1;
  assign CLBLL_R_X73Y132_SLICE_X110Y132_D4 = 1'b1;
  assign CLBLL_R_X73Y132_SLICE_X110Y132_D5 = 1'b1;
  assign CLBLL_R_X73Y132_SLICE_X110Y132_D6 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_A6 = 1'b1;
  assign CLBLM_L_X74Y104_SLICE_X113Y104_D1 = 1'b1;
  assign CLBLM_L_X74Y104_SLICE_X113Y104_D2 = 1'b1;
  assign CLBLM_L_X74Y104_SLICE_X113Y104_D3 = 1'b1;
  assign CLBLM_L_X74Y104_SLICE_X113Y104_D4 = 1'b1;
  assign CLBLM_L_X74Y104_SLICE_X112Y104_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y104_SLICE_X112Y104_A2 = CLBLM_L_X72Y103_SLICE_X108Y103_BO6;
  assign CLBLM_L_X74Y104_SLICE_X112Y104_A3 = CLBLM_L_X74Y104_SLICE_X112Y104_AQ;
  assign CLBLM_L_X74Y104_SLICE_X112Y104_A4 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X74Y104_SLICE_X112Y104_A5 = CLBLM_L_X74Y103_SLICE_X112Y103_BQ;
  assign CLBLM_L_X74Y104_SLICE_X112Y104_A6 = CLBLL_R_X73Y104_SLICE_X110Y104_DO5;
  assign CLBLM_L_X74Y104_SLICE_X112Y104_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y104_SLICE_X112Y104_B2 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X74Y104_SLICE_X112Y104_B3 = CLBLM_L_X74Y104_SLICE_X112Y104_AQ;
  assign CLBLM_L_X74Y104_SLICE_X112Y104_B4 = CLBLM_L_X72Y103_SLICE_X108Y103_BO5;
  assign CLBLM_L_X74Y104_SLICE_X112Y104_B5 = CLBLL_R_X73Y104_SLICE_X110Y104_DO5;
  assign CLBLM_L_X74Y104_SLICE_X112Y104_B6 = CLBLM_L_X74Y104_SLICE_X112Y104_BQ;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y132_SLICE_X111Y132_A1 = CLBLM_L_X74Y135_SLICE_X113Y135_BQ;
  assign CLBLL_R_X73Y132_SLICE_X111Y132_A2 = CLBLM_L_X76Y133_SLICE_X116Y133_BQ;
  assign CLBLL_R_X73Y132_SLICE_X111Y132_A3 = CLBLM_L_X76Y130_SLICE_X116Y130_DQ;
  assign CLBLL_R_X73Y132_SLICE_X111Y132_A4 = CLBLM_L_X76Y125_SLICE_X117Y125_BQ;
  assign CLBLL_R_X73Y132_SLICE_X111Y132_A5 = CLBLL_R_X75Y133_SLICE_X115Y133_AQ;
  assign CLBLL_R_X73Y132_SLICE_X111Y132_A6 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_B2 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_B3 = CLBLM_L_X70Y123_SLICE_X104Y123_AQ;
  assign CLBLM_L_X74Y104_SLICE_X112Y104_C1 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLL_R_X73Y132_SLICE_X111Y132_B1 = CLBLL_R_X75Y133_SLICE_X115Y133_AQ;
  assign CLBLL_R_X73Y132_SLICE_X111Y132_B2 = CLBLM_L_X76Y125_SLICE_X117Y125_BQ;
  assign CLBLL_R_X73Y132_SLICE_X111Y132_B3 = CLBLM_L_X76Y130_SLICE_X116Y130_DQ;
  assign CLBLL_R_X73Y132_SLICE_X111Y132_B4 = CLBLM_L_X76Y133_SLICE_X116Y133_BQ;
  assign CLBLL_R_X73Y132_SLICE_X111Y132_B5 = CLBLM_L_X74Y133_SLICE_X112Y133_AQ;
  assign CLBLL_R_X73Y132_SLICE_X111Y132_B6 = CLBLM_L_X74Y135_SLICE_X113Y135_BQ;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_B4 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_B5 = 1'b1;
  assign CLBLL_R_X73Y132_SLICE_X111Y132_C1 = CLBLM_L_X74Y132_SLICE_X113Y132_BQ;
  assign CLBLL_R_X73Y132_SLICE_X111Y132_C2 = CLBLM_L_X76Y133_SLICE_X116Y133_BQ;
  assign CLBLL_R_X73Y132_SLICE_X111Y132_C3 = CLBLM_L_X76Y125_SLICE_X117Y125_BQ;
  assign CLBLL_R_X73Y132_SLICE_X111Y132_C4 = CLBLM_L_X74Y135_SLICE_X113Y135_BQ;
  assign CLBLL_R_X73Y132_SLICE_X111Y132_C5 = CLBLL_R_X75Y133_SLICE_X115Y133_AQ;
  assign CLBLL_R_X73Y132_SLICE_X111Y132_C6 = CLBLM_L_X76Y130_SLICE_X116Y130_DQ;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_B6 = 1'b1;
  assign CLBLM_L_X74Y104_SLICE_X112Y104_D3 = 1'b1;
  assign CLBLM_L_X74Y104_SLICE_X112Y104_D4 = 1'b1;
  assign CLBLM_L_X74Y104_SLICE_X112Y104_D5 = 1'b1;
  assign CLBLM_L_X74Y104_SLICE_X112Y104_D6 = 1'b1;
  assign CLBLM_L_X74Y104_SLICE_X112Y104_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X73Y132_SLICE_X111Y132_D1 = 1'b1;
  assign CLBLL_R_X73Y132_SLICE_X111Y132_D2 = 1'b1;
  assign CLBLL_R_X73Y132_SLICE_X111Y132_D3 = 1'b1;
  assign CLBLL_R_X73Y132_SLICE_X111Y132_D4 = 1'b1;
  assign CLBLL_R_X73Y132_SLICE_X111Y132_D5 = 1'b1;
  assign CLBLL_R_X73Y132_SLICE_X111Y132_D6 = 1'b1;
  assign CLBLM_R_X67Y116_SLICE_X101Y116_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y116_SLICE_X101Y116_A2 = CLBLM_R_X67Y115_SLICE_X100Y115_AQ;
  assign CLBLM_R_X67Y116_SLICE_X101Y116_A3 = CLBLM_R_X67Y116_SLICE_X101Y116_AQ;
  assign CLBLM_R_X67Y116_SLICE_X101Y116_A4 = CLBLM_R_X67Y115_SLICE_X100Y115_A5Q;
  assign CLBLM_R_X67Y116_SLICE_X101Y116_A5 = CLBLM_R_X67Y116_SLICE_X101Y116_A5Q;
  assign CLBLM_R_X67Y116_SLICE_X101Y116_A6 = 1'b1;
  assign CLBLM_R_X67Y116_SLICE_X101Y116_B1 = 1'b1;
  assign CLBLM_R_X67Y116_SLICE_X101Y116_B2 = CLBLM_R_X67Y115_SLICE_X100Y115_AQ;
  assign CLBLM_R_X67Y116_SLICE_X101Y116_B3 = CLBLM_R_X67Y116_SLICE_X101Y116_AQ;
  assign CLBLM_R_X67Y116_SLICE_X101Y116_B4 = 1'b1;
  assign CLBLM_R_X67Y116_SLICE_X101Y116_B5 = CLBLM_R_X67Y115_SLICE_X100Y115_A5Q;
  assign CLBLM_R_X67Y116_SLICE_X101Y116_B6 = 1'b1;
  assign CLBLM_R_X67Y116_SLICE_X101Y116_BX = CLBLM_R_X67Y116_SLICE_X100Y116_B5Q;
  assign CLBLM_R_X67Y116_SLICE_X101Y116_C1 = 1'b1;
  assign CLBLM_R_X67Y116_SLICE_X101Y116_C2 = 1'b1;
  assign CLBLM_R_X67Y116_SLICE_X101Y116_C3 = 1'b1;
  assign CLBLM_R_X67Y116_SLICE_X101Y116_C4 = 1'b1;
  assign CLBLM_R_X67Y116_SLICE_X101Y116_C5 = 1'b1;
  assign CLBLM_R_X67Y116_SLICE_X101Y116_C6 = 1'b1;
  assign CLBLM_R_X67Y116_SLICE_X101Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X67Y116_SLICE_X101Y116_D1 = 1'b1;
  assign CLBLM_R_X67Y116_SLICE_X101Y116_D2 = 1'b1;
  assign CLBLM_R_X67Y116_SLICE_X101Y116_D3 = 1'b1;
  assign CLBLM_R_X67Y116_SLICE_X101Y116_D4 = 1'b1;
  assign CLBLM_R_X67Y116_SLICE_X101Y116_D5 = 1'b1;
  assign CLBLM_R_X67Y116_SLICE_X101Y116_D6 = 1'b1;
  assign CLBLM_R_X67Y116_SLICE_X101Y116_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X67Y116_SLICE_X100Y116_A1 = CLBLM_R_X67Y118_SLICE_X100Y118_A5Q;
  assign CLBLM_R_X67Y116_SLICE_X100Y116_A2 = CLBLM_R_X67Y116_SLICE_X101Y116_BO6;
  assign CLBLM_R_X67Y116_SLICE_X100Y116_A3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y116_SLICE_X100Y116_A4 = CLBLM_R_X67Y116_SLICE_X101Y116_BQ;
  assign CLBLM_R_X67Y116_SLICE_X100Y116_A5 = CLBLM_R_X67Y116_SLICE_X100Y116_C5Q;
  assign CLBLM_R_X67Y116_SLICE_X100Y116_A6 = 1'b1;
  assign CLBLM_R_X67Y116_SLICE_X100Y116_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y116_SLICE_X100Y116_B2 = CLBLM_R_X67Y116_SLICE_X100Y116_BQ;
  assign CLBLM_R_X67Y116_SLICE_X100Y116_B3 = CLBLM_R_X67Y115_SLICE_X100Y115_A5Q;
  assign CLBLM_R_X67Y116_SLICE_X100Y116_B4 = CLBLM_R_X67Y115_SLICE_X100Y115_AQ;
  assign CLBLM_R_X67Y116_SLICE_X100Y116_B5 = CLBLM_R_X67Y116_SLICE_X101Y116_AQ;
  assign CLBLM_R_X67Y116_SLICE_X100Y116_B6 = 1'b1;
  assign CLBLM_R_X67Y116_SLICE_X100Y116_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y116_SLICE_X100Y116_C2 = CLBLM_R_X67Y116_SLICE_X100Y116_AQ;
  assign CLBLM_R_X67Y116_SLICE_X100Y116_C3 = CLBLM_R_X67Y116_SLICE_X100Y116_BQ;
  assign CLBLM_R_X67Y116_SLICE_X100Y116_C4 = CLBLM_R_X67Y116_SLICE_X101Y116_BQ;
  assign CLBLM_R_X67Y116_SLICE_X100Y116_C5 = CLBLM_R_X67Y116_SLICE_X100Y116_DO6;
  assign CLBLM_R_X67Y116_SLICE_X100Y116_C6 = 1'b1;
  assign CLBLM_R_X67Y116_SLICE_X100Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X67Y116_SLICE_X100Y116_D1 = CLBLM_R_X67Y116_SLICE_X101Y116_AQ;
  assign CLBLM_R_X67Y116_SLICE_X100Y116_D2 = CLBLM_R_X67Y116_SLICE_X101Y116_A5Q;
  assign CLBLM_R_X67Y116_SLICE_X100Y116_D3 = CLBLM_R_X67Y115_SLICE_X100Y115_AQ;
  assign CLBLM_R_X67Y116_SLICE_X100Y116_D4 = CLBLM_R_X67Y115_SLICE_X100Y115_A5Q;
  assign CLBLM_R_X67Y116_SLICE_X100Y116_D5 = CLBLM_R_X67Y116_SLICE_X100Y116_B5Q;
  assign CLBLM_R_X67Y116_SLICE_X100Y116_D6 = CLBLM_R_X67Y116_SLICE_X101Y116_BQ;
  assign CLBLM_R_X67Y116_SLICE_X100Y116_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_D6 = 1'b1;
  assign LIOI3_X0Y83_OLOGIC_X0Y84_D1 = CLBLM_L_X60Y99_SLICE_X90Y99_CQ;
  assign LIOI3_X0Y83_OLOGIC_X0Y84_T1 = 1'b1;
  assign RIOI3_X105Y127_OLOGIC_X1Y128_D1 = CLBLM_R_X65Y110_SLICE_X99Y110_CQ;
  assign LIOI3_X0Y83_OLOGIC_X0Y83_D1 = CLBLM_L_X70Y99_SLICE_X104Y99_AQ;
  assign RIOI3_X105Y127_OLOGIC_X1Y128_T1 = 1'b1;
  assign LIOI3_X0Y83_OLOGIC_X0Y83_T1 = 1'b1;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_D1 = CLBLM_L_X72Y107_SLICE_X108Y107_A5Q;
  assign CLBLM_R_X67Y103_SLICE_X101Y103_D4 = 1'b1;
  assign CLBLM_R_X67Y103_SLICE_X101Y103_D5 = 1'b1;
  assign CLBLM_R_X67Y103_SLICE_X101Y103_D6 = 1'b1;
  assign LIOB33_X0Y127_IOB_X0Y127_O = CLBLL_L_X34Y126_SLICE_X50Y126_AO6;
  assign LIOB33_X0Y127_IOB_X0Y128_O = CLBLL_R_X73Y131_SLICE_X110Y131_AQ;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_T1 = 1'b1;
  assign CLBLL_R_X73Y133_SLICE_X110Y133_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y133_SLICE_X110Y133_A2 = CLBLL_R_X75Y133_SLICE_X114Y133_CO5;
  assign CLBLL_R_X73Y133_SLICE_X110Y133_A3 = CLBLL_R_X73Y133_SLICE_X110Y133_AQ;
  assign CLBLL_R_X73Y133_SLICE_X110Y133_A4 = CLBLL_R_X75Y133_SLICE_X115Y133_BQ;
  assign CLBLL_R_X73Y133_SLICE_X110Y133_A5 = CLBLL_R_X73Y133_SLICE_X110Y133_A5Q;
  assign CLBLL_R_X73Y133_SLICE_X110Y133_A6 = 1'b1;
  assign CLBLL_R_X73Y133_SLICE_X110Y133_B1 = CLBLM_L_X72Y133_SLICE_X108Y133_A5Q;
  assign CLBLL_R_X73Y133_SLICE_X110Y133_B2 = CLBLL_R_X73Y133_SLICE_X110Y133_BQ;
  assign CLBLL_R_X73Y133_SLICE_X110Y133_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y133_SLICE_X110Y133_B4 = CLBLM_L_X72Y133_SLICE_X108Y133_AQ;
  assign CLBLL_R_X73Y133_SLICE_X110Y133_B5 = CLBLL_R_X73Y132_SLICE_X110Y132_BO6;
  assign CLBLL_R_X73Y133_SLICE_X110Y133_B6 = CLBLL_R_X73Y132_SLICE_X110Y132_AO5;
  assign CLBLM_R_X67Y103_SLICE_X101Y103_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X73Y133_SLICE_X110Y133_C1 = CLBLL_R_X73Y133_SLICE_X110Y133_A5Q;
  assign CLBLL_R_X73Y133_SLICE_X110Y133_C2 = CLBLL_R_X73Y133_SLICE_X110Y133_AQ;
  assign CLBLL_R_X73Y133_SLICE_X110Y133_C3 = CLBLL_R_X75Y133_SLICE_X114Y133_AQ;
  assign CLBLL_R_X73Y133_SLICE_X110Y133_C4 = CLBLM_L_X70Y136_SLICE_X105Y136_A5Q;
  assign CLBLL_R_X73Y133_SLICE_X110Y133_C5 = 1'b1;
  assign CLBLL_R_X73Y133_SLICE_X110Y133_C6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y133_SLICE_X110Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X73Y133_SLICE_X110Y133_D1 = CLBLM_L_X74Y135_SLICE_X113Y135_BQ;
  assign CLBLL_R_X73Y133_SLICE_X110Y133_D2 = CLBLL_R_X73Y133_SLICE_X110Y133_CQ;
  assign CLBLL_R_X73Y133_SLICE_X110Y133_D3 = CLBLL_R_X75Y133_SLICE_X115Y133_AQ;
  assign CLBLL_R_X73Y133_SLICE_X110Y133_D4 = 1'b1;
  assign CLBLL_R_X73Y133_SLICE_X110Y133_D5 = CLBLM_L_X74Y134_SLICE_X113Y134_AQ;
  assign CLBLL_R_X73Y133_SLICE_X110Y133_D6 = CLBLM_L_X76Y133_SLICE_X116Y133_BQ;
  assign CLBLL_R_X73Y133_SLICE_X110Y133_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X103Y76_SLICE_X162Y76_C4 = 1'b1;
  assign LIOI3_X0Y55_OLOGIC_X0Y56_D1 = CLBLM_L_X62Y92_SLICE_X92Y92_BQ;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_T1 = 1'b1;
  assign CLBLL_R_X73Y133_SLICE_X111Y133_A1 = CLBLL_R_X73Y133_SLICE_X111Y133_DO6;
  assign CLBLL_R_X73Y133_SLICE_X111Y133_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y133_SLICE_X111Y133_A3 = CLBLL_R_X73Y133_SLICE_X111Y133_AQ;
  assign CLBLL_R_X73Y133_SLICE_X111Y133_A4 = CLBLM_L_X74Y132_SLICE_X112Y132_BO6;
  assign CLBLL_R_X73Y133_SLICE_X111Y133_A5 = CLBLM_L_X74Y134_SLICE_X113Y134_AQ;
  assign CLBLL_R_X73Y133_SLICE_X111Y133_A6 = CLBLM_L_X74Y134_SLICE_X112Y134_AO5;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_D3 = 1'b1;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_D4 = 1'b1;
  assign CLBLL_R_X73Y133_SLICE_X111Y133_AX = CLBLM_L_X60Y94_SLICE_X90Y94_AQ;
  assign LIOB33_X0Y123_IOB_X0Y123_O = CLBLM_R_X67Y108_SLICE_X100Y108_AO6;
  assign CLBLL_R_X73Y133_SLICE_X111Y133_B1 = CLBLL_R_X75Y133_SLICE_X115Y133_AQ;
  assign CLBLL_R_X73Y133_SLICE_X111Y133_B2 = CLBLM_L_X76Y130_SLICE_X116Y130_DQ;
  assign CLBLL_R_X73Y133_SLICE_X111Y133_B3 = CLBLM_L_X76Y125_SLICE_X117Y125_BQ;
  assign CLBLL_R_X73Y133_SLICE_X111Y133_B4 = CLBLM_L_X74Y134_SLICE_X113Y134_AQ;
  assign CLBLL_R_X73Y133_SLICE_X111Y133_B5 = CLBLM_L_X74Y135_SLICE_X113Y135_BQ;
  assign CLBLL_R_X73Y133_SLICE_X111Y133_B6 = CLBLM_L_X76Y133_SLICE_X116Y133_BQ;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_D5 = 1'b1;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_D6 = 1'b1;
  assign CLBLM_R_X103Y76_SLICE_X162Y76_C5 = 1'b1;
  assign CLBLL_R_X73Y133_SLICE_X111Y133_C1 = CLBLM_L_X76Y133_SLICE_X116Y133_BQ;
  assign CLBLL_R_X73Y133_SLICE_X111Y133_C2 = CLBLM_L_X74Y135_SLICE_X113Y135_BQ;
  assign CLBLL_R_X73Y133_SLICE_X111Y133_C3 = CLBLM_L_X74Y133_SLICE_X112Y133_CQ;
  assign CLBLL_R_X73Y133_SLICE_X111Y133_C4 = CLBLL_R_X75Y133_SLICE_X115Y133_AQ;
  assign CLBLL_R_X73Y133_SLICE_X111Y133_C5 = CLBLM_L_X76Y125_SLICE_X117Y125_BQ;
  assign CLBLL_R_X73Y133_SLICE_X111Y133_C6 = CLBLM_L_X76Y130_SLICE_X116Y130_DQ;
  assign CLBLL_R_X73Y133_SLICE_X111Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOB33_X105Y105_IOB_X1Y106_O = CLBLL_R_X75Y103_SLICE_X115Y103_AQ;
  assign CLBLL_R_X73Y133_SLICE_X111Y133_D1 = CLBLM_L_X74Y135_SLICE_X113Y135_BQ;
  assign CLBLL_R_X73Y133_SLICE_X111Y133_D2 = CLBLM_L_X76Y133_SLICE_X116Y133_BQ;
  assign CLBLL_R_X73Y133_SLICE_X111Y133_D3 = 1'b1;
  assign CLBLL_R_X73Y133_SLICE_X111Y133_D4 = CLBLL_R_X73Y133_SLICE_X110Y133_CQ;
  assign CLBLL_R_X73Y133_SLICE_X111Y133_D5 = CLBLL_R_X75Y133_SLICE_X115Y133_AQ;
  assign CLBLL_R_X73Y133_SLICE_X111Y133_D6 = CLBLM_L_X74Y133_SLICE_X112Y133_AQ;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X103Y76_SLICE_X162Y76_C6 = 1'b1;
  assign CLBLL_R_X73Y133_SLICE_X111Y133_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign LIOI3_X0Y55_OLOGIC_X0Y56_T1 = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_D1 = CLBLM_R_X65Y106_SLICE_X99Y106_DQ;
  assign CLBLM_L_X68Y108_SLICE_X103Y108_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y108_SLICE_X103Y108_A6 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_A1 = CLBLM_L_X64Y106_SLICE_X96Y106_BQ;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_A2 = CLBLM_L_X62Y107_SLICE_X93Y107_CO6;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_A3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_A4 = CLBLM_R_X67Y103_SLICE_X100Y103_BQ;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_A5 = CLBLM_R_X63Y105_SLICE_X95Y105_A5Q;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_A6 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_B1 = CLBLM_R_X63Y107_SLICE_X95Y107_DQ;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_B2 = CLBLM_R_X63Y105_SLICE_X95Y105_BQ;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_B3 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_B4 = CLBLM_L_X64Y106_SLICE_X96Y106_DO5;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_B6 = CLBLM_L_X64Y105_SLICE_X96Y105_BO6;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_C1 = CLBLM_R_X63Y105_SLICE_X95Y105_C5Q;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_C2 = CLBLM_R_X63Y105_SLICE_X95Y105_CQ;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_C3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_C4 = CLBLM_R_X63Y105_SLICE_X95Y105_A5Q;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_C5 = CLBLM_L_X62Y107_SLICE_X93Y107_CO6;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_C6 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_D1 = CLBLM_L_X64Y105_SLICE_X97Y105_BQ;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_D2 = CLBLM_R_X63Y105_SLICE_X95Y105_CQ;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_D3 = CLBLM_L_X64Y105_SLICE_X97Y105_DO6;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_D4 = CLBLM_R_X63Y105_SLICE_X94Y105_CQ;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_D5 = CLBLM_R_X63Y105_SLICE_X95Y105_C5Q;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_D6 = CLBLM_R_X63Y105_SLICE_X94Y105_C5Q;
  assign LIOI3_X0Y55_OLOGIC_X0Y55_D1 = CLBLM_L_X60Y97_SLICE_X91Y97_AQ;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_T1 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_A1 = CLBLM_L_X64Y105_SLICE_X96Y105_AO6;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_A2 = CLBLM_L_X62Y105_SLICE_X93Y105_BQ;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_A3 = CLBLM_R_X63Y105_SLICE_X94Y105_AQ;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_A5 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_A6 = CLBLM_L_X64Y106_SLICE_X96Y106_DO5;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_B1 = CLBLM_L_X64Y106_SLICE_X97Y106_AO6;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_B2 = CLBLM_R_X63Y105_SLICE_X94Y105_BQ;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_B3 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_B4 = CLBLM_R_X63Y105_SLICE_X95Y105_BQ;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_B5 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_B5 = CLBLL_R_X71Y119_SLICE_X106Y119_A5Q;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_B6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X68Y108_SLICE_X103Y108_C1 = CLBLM_L_X68Y106_SLICE_X103Y106_BQ;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_B6 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_C1 = CLBLM_R_X63Y105_SLICE_X94Y105_C5Q;
  assign CLBLM_L_X68Y108_SLICE_X103Y108_C2 = CLBLM_L_X68Y106_SLICE_X103Y106_B5Q;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_C2 = CLBLM_R_X63Y105_SLICE_X94Y105_CQ;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_C3 = CLBLM_R_X63Y105_SLICE_X95Y105_C5Q;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_C4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_C5 = CLBLM_L_X64Y105_SLICE_X97Y105_DO6;
  assign CLBLM_L_X68Y108_SLICE_X103Y108_C3 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_C6 = 1'b1;
  assign CLBLM_R_X103Y76_SLICE_X162Y76_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X68Y108_SLICE_X103Y108_C4 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_D1 = CLBLM_R_X63Y105_SLICE_X94Y105_C5Q;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_D2 = CLBLM_R_X63Y105_SLICE_X94Y105_CQ;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_D3 = CLBLM_L_X62Y107_SLICE_X93Y107_A5Q;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_D4 = CLBLM_L_X62Y105_SLICE_X93Y105_BQ;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_D5 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_D6 = CLBLM_R_X63Y105_SLICE_X94Y105_AQ;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign LIOI3_X0Y55_OLOGIC_X0Y55_T1 = 1'b1;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_C3 = CLBLM_L_X74Y119_SLICE_X112Y119_AQ;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_C5 = CLBLM_L_X72Y118_SLICE_X108Y118_B5Q;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_C6 = 1'b1;
  assign LIOB33_X0Y129_IOB_X0Y130_O = 1'b1;
  assign LIOB33_X0Y129_IOB_X0Y129_O = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X73Y134_SLICE_X110Y134_A1 = CLBLM_L_X74Y134_SLICE_X113Y134_CQ;
  assign CLBLL_R_X73Y134_SLICE_X110Y134_A2 = CLBLM_L_X70Y136_SLICE_X105Y136_CO6;
  assign CLBLL_R_X73Y134_SLICE_X110Y134_A3 = CLBLL_R_X73Y133_SLICE_X110Y133_A5Q;
  assign CLBLL_R_X73Y134_SLICE_X110Y134_A4 = CLBLM_L_X74Y134_SLICE_X113Y134_A5Q;
  assign CLBLL_R_X73Y134_SLICE_X110Y134_A5 = CLBLL_R_X71Y134_SLICE_X106Y134_AQ;
  assign CLBLL_R_X73Y134_SLICE_X110Y134_A6 = 1'b1;
  assign CLBLL_R_X73Y134_SLICE_X110Y134_B1 = 1'b1;
  assign CLBLL_R_X73Y134_SLICE_X110Y134_B2 = 1'b1;
  assign CLBLL_R_X73Y134_SLICE_X110Y134_B3 = 1'b1;
  assign CLBLL_R_X73Y134_SLICE_X110Y134_B4 = 1'b1;
  assign CLBLL_R_X73Y134_SLICE_X110Y134_B5 = 1'b1;
  assign CLBLL_R_X73Y134_SLICE_X110Y134_B6 = 1'b1;
  assign CLBLL_R_X73Y134_SLICE_X110Y134_C1 = 1'b1;
  assign CLBLL_R_X73Y134_SLICE_X110Y134_C2 = 1'b1;
  assign CLBLL_R_X73Y134_SLICE_X110Y134_C3 = 1'b1;
  assign CLBLL_R_X73Y134_SLICE_X110Y134_C4 = 1'b1;
  assign CLBLL_R_X73Y134_SLICE_X110Y134_C5 = 1'b1;
  assign CLBLL_R_X73Y134_SLICE_X110Y134_C6 = 1'b1;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_D4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_D5 = CLBLM_L_X72Y117_SLICE_X108Y117_AQ;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_A4 = CLBLM_L_X74Y126_SLICE_X112Y126_BO6;
  assign CLBLL_R_X73Y134_SLICE_X110Y134_D1 = 1'b1;
  assign CLBLL_R_X73Y134_SLICE_X110Y134_D2 = 1'b1;
  assign CLBLL_R_X73Y134_SLICE_X110Y134_D3 = 1'b1;
  assign CLBLL_R_X73Y134_SLICE_X110Y134_D4 = 1'b1;
  assign CLBLL_R_X73Y134_SLICE_X110Y134_D5 = 1'b1;
  assign CLBLL_R_X73Y134_SLICE_X110Y134_D6 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y134_SLICE_X111Y134_A1 = CLBLM_L_X74Y132_SLICE_X112Y132_A5Q;
  assign CLBLL_R_X73Y134_SLICE_X111Y134_A2 = CLBLL_R_X73Y133_SLICE_X110Y133_DO6;
  assign CLBLL_R_X73Y134_SLICE_X111Y134_A3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X73Y134_SLICE_X111Y134_A4 = CLBLM_L_X74Y132_SLICE_X112Y132_AQ;
  assign CLBLL_R_X73Y134_SLICE_X111Y134_A5 = CLBLM_L_X74Y134_SLICE_X112Y134_AO6;
  assign CLBLL_R_X73Y134_SLICE_X111Y134_A6 = CLBLL_R_X73Y134_SLICE_X111Y134_AQ;
  assign CLBLL_R_X73Y134_SLICE_X111Y134_B1 = 1'b1;
  assign CLBLL_R_X73Y134_SLICE_X111Y134_B2 = 1'b1;
  assign CLBLL_R_X73Y134_SLICE_X111Y134_B3 = 1'b1;
  assign CLBLL_R_X73Y134_SLICE_X111Y134_B4 = 1'b1;
  assign CLBLL_R_X73Y134_SLICE_X111Y134_B5 = 1'b1;
  assign CLBLL_R_X73Y134_SLICE_X111Y134_B6 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_A6 = CLBLL_R_X73Y126_SLICE_X111Y126_AQ;
  assign CLBLL_R_X73Y134_SLICE_X111Y134_C1 = 1'b1;
  assign CLBLL_R_X73Y134_SLICE_X111Y134_C2 = 1'b1;
  assign CLBLL_R_X73Y134_SLICE_X111Y134_C3 = 1'b1;
  assign CLBLL_R_X73Y134_SLICE_X111Y134_C4 = 1'b1;
  assign CLBLL_R_X73Y134_SLICE_X111Y134_C5 = 1'b1;
  assign CLBLL_R_X73Y134_SLICE_X111Y134_C6 = 1'b1;
  assign CLBLL_R_X73Y134_SLICE_X111Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X73Y134_SLICE_X111Y134_D1 = 1'b1;
  assign CLBLL_R_X73Y134_SLICE_X111Y134_D2 = 1'b1;
  assign CLBLL_R_X73Y134_SLICE_X111Y134_D3 = 1'b1;
  assign CLBLL_R_X73Y134_SLICE_X111Y134_D4 = 1'b1;
  assign CLBLL_R_X73Y134_SLICE_X111Y134_D5 = 1'b1;
  assign CLBLL_R_X73Y134_SLICE_X111Y134_D6 = 1'b1;
  assign CLBLL_R_X73Y134_SLICE_X111Y134_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X67Y118_SLICE_X101Y118_A1 = 1'b1;
  assign CLBLM_R_X67Y118_SLICE_X101Y118_A2 = CLBLM_R_X67Y118_SLICE_X101Y118_BQ;
  assign CLBLM_R_X67Y118_SLICE_X101Y118_A3 = CLBLM_R_X67Y118_SLICE_X101Y118_AQ;
  assign CLBLM_R_X67Y118_SLICE_X101Y118_A4 = CLBLM_R_X67Y116_SLICE_X100Y116_CQ;
  assign CLBLM_R_X67Y118_SLICE_X101Y118_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y118_SLICE_X101Y118_A6 = 1'b1;
  assign CLBLM_R_X67Y118_SLICE_X101Y118_B1 = 1'b1;
  assign CLBLM_R_X67Y118_SLICE_X101Y118_B2 = 1'b1;
  assign CLBLM_R_X67Y118_SLICE_X101Y118_B3 = 1'b1;
  assign CLBLM_R_X67Y118_SLICE_X101Y118_B4 = 1'b1;
  assign CLBLM_R_X67Y118_SLICE_X101Y118_B5 = 1'b1;
  assign CLBLM_R_X67Y118_SLICE_X101Y118_B6 = 1'b1;
  assign CLBLM_R_X67Y118_SLICE_X101Y118_BX = CLBLM_R_X67Y118_SLICE_X101Y118_AQ;
  assign CLBLM_R_X67Y118_SLICE_X101Y118_C1 = 1'b1;
  assign CLBLM_R_X67Y118_SLICE_X101Y118_C2 = 1'b1;
  assign CLBLM_R_X67Y118_SLICE_X101Y118_C3 = 1'b1;
  assign CLBLM_R_X67Y118_SLICE_X101Y118_C4 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_A1 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_A2 = CLBLM_R_X63Y105_SLICE_X94Y105_BQ;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_A3 = CLBLM_R_X63Y106_SLICE_X95Y106_AQ;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_A5 = CLBLM_L_X64Y105_SLICE_X97Y105_DO6;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_A6 = CLBLM_L_X62Y106_SLICE_X93Y106_DO6;
  assign CLBLM_R_X67Y118_SLICE_X101Y118_C5 = 1'b1;
  assign CLBLM_R_X67Y118_SLICE_X101Y118_C6 = 1'b1;
  assign CLBLM_R_X67Y118_SLICE_X101Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_B1 = CLBLM_L_X64Y105_SLICE_X96Y105_AO6;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_B2 = CLBLM_R_X63Y106_SLICE_X95Y106_BQ;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_B3 = CLBLM_L_X62Y106_SLICE_X93Y106_BQ;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_B5 = CLBLM_L_X64Y106_SLICE_X96Y106_BO6;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_B6 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X67Y118_SLICE_X101Y118_D1 = 1'b1;
  assign CLBLM_L_X68Y108_SLICE_X102Y108_C4 = CLBLM_L_X68Y108_SLICE_X102Y108_A5Q;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_C2 = CLBLM_R_X63Y106_SLICE_X95Y106_CQ;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_C3 = CLBLM_L_X64Y106_SLICE_X97Y106_C5Q;
  assign CLBLM_L_X68Y108_SLICE_X102Y108_C5 = CLBLM_L_X68Y108_SLICE_X102Y108_B5Q;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_C4 = CLBLM_L_X64Y105_SLICE_X96Y105_AO5;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_C5 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_C6 = CLBLM_R_X63Y107_SLICE_X94Y107_BQ;
  assign CLBLM_R_X67Y118_SLICE_X100Y118_A1 = CLBLM_R_X67Y118_SLICE_X101Y118_A5Q;
  assign CLBLM_L_X68Y108_SLICE_X102Y108_C6 = CLBLM_L_X68Y108_SLICE_X103Y108_BQ;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X67Y118_SLICE_X100Y118_A2 = CLBLM_R_X67Y116_SLICE_X100Y116_CQ;
  assign CLBLM_R_X67Y118_SLICE_X100Y118_A3 = CLBLM_R_X67Y118_SLICE_X100Y118_AQ;
  assign CLBLM_R_X67Y118_SLICE_X100Y118_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X67Y118_SLICE_X100Y118_A5 = CLBLM_R_X67Y118_SLICE_X100Y118_A5Q;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_D1 = CLBLM_R_X63Y107_SLICE_X95Y107_AQ;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_D2 = CLBLM_R_X63Y106_SLICE_X95Y106_CQ;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_D3 = CLBLM_L_X62Y106_SLICE_X93Y106_AQ;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_D4 = CLBLM_L_X64Y106_SLICE_X96Y106_BQ;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_D5 = CLBLM_R_X63Y105_SLICE_X94Y105_CQ;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_AX = CLBLM_L_X74Y126_SLICE_X112Y126_CO5;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_D6 = CLBLM_R_X63Y105_SLICE_X94Y105_C5Q;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X67Y118_SLICE_X100Y118_B2 = 1'b1;
  assign CLBLM_R_X67Y118_SLICE_X100Y118_B3 = 1'b1;
  assign CLBLM_R_X67Y118_SLICE_X100Y118_B4 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_A1 = CLBLM_R_X63Y105_SLICE_X94Y105_CQ;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_A2 = CLBLM_R_X63Y105_SLICE_X94Y105_C5Q;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_A3 = CLBLM_R_X63Y105_SLICE_X95Y105_A5Q;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_A4 = CLBLM_L_X60Y101_SLICE_X90Y101_BQ;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_A5 = CLBLM_L_X64Y105_SLICE_X97Y105_DO6;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_A6 = 1'b1;
  assign CLBLM_R_X67Y118_SLICE_X100Y118_C1 = 1'b1;
  assign CLBLM_R_X67Y118_SLICE_X100Y118_C2 = 1'b1;
  assign CLBLM_R_X67Y118_SLICE_X100Y118_C3 = 1'b1;
  assign CLBLM_R_X67Y118_SLICE_X100Y118_C4 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_B1 = CLBLM_L_X64Y106_SLICE_X97Y106_C5Q;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_B2 = CLBLM_R_X63Y106_SLICE_X94Y106_BQ;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_B3 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_B5 = CLBLM_R_X63Y105_SLICE_X94Y105_AQ;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_B6 = CLBLM_L_X64Y105_SLICE_X96Y105_AO6;
  assign CLBLM_R_X67Y118_SLICE_X100Y118_D1 = 1'b1;
  assign CLBLM_R_X67Y118_SLICE_X100Y118_D2 = 1'b1;
  assign CLBLM_R_X67Y118_SLICE_X100Y118_D3 = 1'b1;
  assign CLBLM_R_X67Y118_SLICE_X100Y118_D4 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_C1 = CLBLM_R_X63Y106_SLICE_X94Y106_BQ;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_C2 = CLBLM_L_X60Y101_SLICE_X90Y101_BQ;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_C3 = CLBLM_L_X64Y106_SLICE_X96Y106_A5Q;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_C4 = CLBLM_R_X63Y105_SLICE_X94Y105_CQ;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_C5 = CLBLM_R_X63Y105_SLICE_X94Y105_C5Q;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_C6 = CLBLM_R_X63Y107_SLICE_X94Y107_BQ;
  assign CLBLM_R_X67Y118_SLICE_X100Y118_D6 = 1'b1;
  assign CLBLM_R_X67Y118_SLICE_X100Y118_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_D1 = CLBLM_L_X62Y106_SLICE_X93Y106_BQ;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_D2 = CLBLM_R_X63Y105_SLICE_X94Y105_BQ;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_D3 = CLBLM_R_X63Y105_SLICE_X95Y105_A5Q;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_D4 = CLBLM_R_X63Y106_SLICE_X94Y106_AO5;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_B1 = CLBLM_L_X74Y126_SLICE_X113Y126_A5Q;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_D5 = CLBLM_L_X62Y106_SLICE_X93Y106_AO6;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_D6 = CLBLM_L_X64Y106_SLICE_X96Y106_BQ;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign LIOB33_X0Y131_IOB_X0Y132_O = CLBLM_L_X70Y134_SLICE_X104Y134_CO5;
  assign LIOB33_X0Y131_IOB_X0Y131_O = CLBLM_L_X62Y107_SLICE_X92Y107_AO5;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_B2 = CLBLM_L_X74Y126_SLICE_X112Y126_A5Q;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_B3 = 1'b1;
  assign CLBLM_R_X103Y69_SLICE_X163Y69_C5 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_B4 = CLBLL_R_X75Y128_SLICE_X115Y128_AO6;
  assign CLBLM_L_X74Y107_SLICE_X113Y107_A1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y107_SLICE_X113Y107_A2 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X74Y107_SLICE_X113Y107_A3 = CLBLM_L_X74Y107_SLICE_X113Y107_AQ;
  assign CLBLM_L_X74Y107_SLICE_X113Y107_A4 = CLBLM_L_X72Y108_SLICE_X109Y108_CO6;
  assign CLBLM_L_X74Y107_SLICE_X113Y107_A5 = CLBLM_L_X72Y108_SLICE_X108Y108_BO5;
  assign CLBLM_L_X74Y107_SLICE_X113Y107_A6 = CLBLM_L_X74Y107_SLICE_X112Y107_CQ;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_B5 = 1'b1;
  assign CLBLM_L_X74Y107_SLICE_X113Y107_B1 = 1'b1;
  assign CLBLM_L_X74Y107_SLICE_X113Y107_B2 = 1'b1;
  assign CLBLM_L_X74Y107_SLICE_X113Y107_B3 = 1'b1;
  assign CLBLM_L_X74Y107_SLICE_X113Y107_B4 = 1'b1;
  assign CLBLM_L_X74Y107_SLICE_X113Y107_B5 = 1'b1;
  assign CLBLM_L_X74Y107_SLICE_X113Y107_B6 = 1'b1;
  assign CLBLM_L_X74Y107_SLICE_X113Y107_C1 = 1'b1;
  assign CLBLM_L_X74Y107_SLICE_X113Y107_C2 = 1'b1;
  assign CLBLM_L_X74Y107_SLICE_X113Y107_C3 = 1'b1;
  assign CLBLM_L_X74Y107_SLICE_X113Y107_C4 = 1'b1;
  assign CLBLM_L_X74Y107_SLICE_X113Y107_C5 = 1'b1;
  assign CLBLM_L_X74Y107_SLICE_X113Y107_C6 = 1'b1;
  assign CLBLM_L_X74Y107_SLICE_X113Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_B6 = 1'b1;
  assign CLBLM_L_X74Y107_SLICE_X113Y107_D1 = 1'b1;
  assign CLBLM_L_X74Y107_SLICE_X113Y107_D2 = 1'b1;
  assign CLBLM_L_X74Y107_SLICE_X113Y107_D3 = 1'b1;
  assign CLBLM_L_X74Y107_SLICE_X113Y107_D4 = 1'b1;
  assign CLBLM_L_X74Y107_SLICE_X113Y107_D5 = 1'b1;
  assign CLBLM_L_X74Y107_SLICE_X113Y107_D6 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X118Y108_A1 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X118Y108_A2 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X118Y108_A3 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X118Y108_A4 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X118Y108_A5 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X118Y108_A6 = 1'b1;
  assign CLBLM_L_X74Y107_SLICE_X112Y107_A1 = CLBLM_L_X72Y109_SLICE_X108Y109_BO6;
  assign CLBLM_L_X74Y107_SLICE_X112Y107_A2 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLL_R_X77Y108_SLICE_X118Y108_AX = CLBLL_R_X71Y100_SLICE_X106Y100_BQ;
  assign CLBLM_L_X74Y107_SLICE_X112Y107_A3 = CLBLM_L_X74Y107_SLICE_X112Y107_AQ;
  assign CLBLL_R_X77Y108_SLICE_X118Y108_B1 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X118Y108_B2 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X118Y108_B3 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X118Y108_B4 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X118Y108_B5 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X118Y108_B6 = 1'b1;
  assign CLBLM_L_X74Y107_SLICE_X112Y107_A4 = CLBLL_R_X73Y107_SLICE_X111Y107_CQ;
  assign CLBLM_L_X74Y107_SLICE_X112Y107_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y107_SLICE_X112Y107_A6 = CLBLM_L_X72Y108_SLICE_X109Y108_CO5;
  assign CLBLL_R_X77Y108_SLICE_X118Y108_C1 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X118Y108_C2 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X118Y108_C3 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X118Y108_C4 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X118Y108_C5 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X118Y108_C6 = 1'b1;
  assign CLBLM_L_X74Y107_SLICE_X112Y107_B2 = CLBLM_L_X74Y107_SLICE_X112Y107_BQ;
  assign CLBLM_L_X74Y107_SLICE_X112Y107_B3 = CLBLM_L_X72Y108_SLICE_X109Y108_BO5;
  assign CLBLL_R_X77Y108_SLICE_X118Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y107_SLICE_X112Y107_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y107_SLICE_X112Y107_B6 = CLBLL_R_X73Y107_SLICE_X110Y107_AQ;
  assign CLBLM_L_X74Y107_SLICE_X112Y107_C1 = CLBLM_L_X72Y108_SLICE_X108Y108_BO5;
  assign CLBLM_L_X74Y107_SLICE_X112Y107_C2 = CLBLM_L_X74Y107_SLICE_X112Y107_CQ;
  assign CLBLL_R_X77Y108_SLICE_X118Y108_D1 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X118Y108_D2 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X118Y108_D3 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X118Y108_D4 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X118Y108_D5 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X118Y108_D6 = 1'b1;
  assign CLBLM_L_X74Y107_SLICE_X112Y107_C6 = CLBLM_L_X72Y108_SLICE_X109Y108_BO5;
  assign CLBLM_L_X74Y107_SLICE_X112Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X77Y108_SLICE_X118Y108_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y107_SLICE_X112Y107_D1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y107_SLICE_X112Y107_D2 = CLBLM_L_X72Y108_SLICE_X108Y108_BO6;
  assign CLBLM_L_X74Y107_SLICE_X112Y107_D3 = CLBLM_L_X74Y107_SLICE_X112Y107_DQ;
  assign CLBLM_L_X74Y107_SLICE_X112Y107_D4 = CLBLM_L_X74Y107_SLICE_X112Y107_BQ;
  assign CLBLM_L_X74Y107_SLICE_X112Y107_D5 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X74Y107_SLICE_X112Y107_D6 = CLBLM_L_X72Y108_SLICE_X109Y108_CO6;
  assign CLBLM_L_X74Y107_SLICE_X112Y107_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_D1 = CLBLM_L_X78Y106_SLICE_X120Y106_AQ;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_T1 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X119Y108_A1 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X119Y108_A2 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X119Y108_A3 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X119Y108_A4 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X119Y108_A5 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X119Y108_A6 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X119Y108_B1 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X119Y108_B2 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X119Y108_B3 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X119Y108_B4 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X119Y108_B5 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X119Y108_B6 = 1'b1;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_D2 = 1'b1;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_D3 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X119Y108_C1 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X119Y108_C2 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X119Y108_C3 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X119Y108_C4 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X119Y108_C5 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X119Y108_C6 = 1'b1;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_D4 = 1'b1;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_D5 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_A4 = CLBLM_L_X64Y106_SLICE_X96Y106_BO6;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_A5 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_A6 = CLBLM_R_X63Y106_SLICE_X94Y106_BQ;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_B1 = CLBLM_L_X64Y105_SLICE_X96Y105_AO5;
  assign CLBLL_R_X77Y108_SLICE_X119Y108_D1 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X119Y108_D2 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X119Y108_D3 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X119Y108_D4 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X119Y108_D5 = 1'b1;
  assign CLBLL_R_X77Y108_SLICE_X119Y108_D6 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_B2 = CLBLM_R_X63Y107_SLICE_X95Y107_BQ;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_B3 = CLBLM_R_X63Y107_SLICE_X95Y107_AQ;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_B5 = CLBLM_L_X64Y106_SLICE_X96Y106_BO5;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_B6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_C1 = CLBLM_L_X64Y106_SLICE_X96Y106_BO5;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_C2 = CLBLM_L_X64Y106_SLICE_X96Y106_CQ;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_C3 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_C4 = CLBLM_L_X64Y105_SLICE_X96Y105_BO6;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_C5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_C6 = CLBLM_R_X63Y107_SLICE_X95Y107_CQ;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_D1 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_D2 = CLBLM_L_X64Y105_SLICE_X96Y105_BO6;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_D3 = CLBLM_R_X63Y107_SLICE_X95Y107_DQ;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_D4 = CLBLM_L_X64Y106_SLICE_X96Y106_DO6;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_D5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_D6 = CLBLM_R_X63Y107_SLICE_X95Y107_CQ;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_A1 = CLBLM_L_X64Y105_SLICE_X96Y105_AO5;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_A3 = CLBLM_R_X63Y107_SLICE_X94Y107_AQ;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_A4 = CLBLM_R_X63Y107_SLICE_X95Y107_BQ;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_A5 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_A6 = CLBLM_L_X64Y106_SLICE_X96Y106_DO6;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_B1 = CLBLM_L_X64Y105_SLICE_X96Y105_AO5;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_B2 = CLBLM_R_X63Y107_SLICE_X94Y107_BQ;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_B3 = CLBLM_R_X63Y107_SLICE_X94Y107_AQ;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_B5 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_B6 = CLBLM_L_X64Y106_SLICE_X96Y106_DO5;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_C1 = CLBLL_R_X75Y107_SLICE_X114Y107_AQ;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_C2 = CLBLM_R_X63Y105_SLICE_X94Y105_DO6;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_C3 = CLBLM_L_X62Y106_SLICE_X93Y106_AO6;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_C4 = CLBLM_R_X63Y107_SLICE_X95Y107_CQ;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_C5 = CLBLM_R_X63Y107_SLICE_X94Y107_DO6;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_C2 = CLBLM_L_X74Y126_SLICE_X113Y126_AQ;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_C6 = CLBLM_L_X62Y107_SLICE_X93Y107_CO5;
  assign LIOB33_X0Y133_IOB_X0Y133_O = CLBLM_R_X63Y105_SLICE_X95Y105_A5Q;
  assign LIOB33_X0Y133_IOB_X0Y134_O = CLBLM_L_X70Y135_SLICE_X104Y135_CO6;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_D1 = CLBLM_R_X63Y105_SLICE_X94Y105_CQ;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_D2 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_D3 = CLBLM_L_X62Y107_SLICE_X93Y107_A5Q;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_D4 = CLBLM_R_X63Y105_SLICE_X94Y105_C5Q;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_D5 = CLBLM_R_X63Y107_SLICE_X95Y107_DQ;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_D6 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y134_SLICE_X113Y134_AX = CLBLM_L_X74Y134_SLICE_X113Y134_DO6;
  assign CLBLM_L_X74Y134_SLICE_X113Y134_B2 = CLBLM_L_X74Y134_SLICE_X113Y134_BQ;
  assign CLBLM_L_X74Y134_SLICE_X113Y134_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y134_SLICE_X113Y134_B6 = CLBLM_L_X74Y132_SLICE_X112Y132_A5Q;
  assign RIOI3_X105Y83_OLOGIC_X1Y84_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_T1 = 1'b1;
  assign CLBLM_L_X74Y134_SLICE_X112Y134_A3 = 1'b1;
  assign CLBLM_L_X74Y134_SLICE_X112Y134_A4 = CLBLM_L_X74Y129_SLICE_X112Y129_BQ;
  assign CLBLM_L_X74Y134_SLICE_X112Y134_A5 = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_T1 = 1'b1;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_B6 = CLBLM_L_X70Y123_SLICE_X104Y123_A5Q;
  assign CLBLM_L_X74Y134_SLICE_X112Y134_B2 = CLBLM_L_X74Y134_SLICE_X112Y134_BQ;
  assign LIOB33_X0Y135_IOB_X0Y135_O = 1'b1;
  assign LIOB33_X0Y135_IOB_X0Y136_O = 1'b1;
  assign CLBLM_L_X74Y134_SLICE_X112Y134_B3 = CLBLM_L_X74Y134_SLICE_X113Y134_A5Q;
  assign CLBLM_L_X74Y134_SLICE_X112Y134_B4 = CLBLL_R_X75Y133_SLICE_X114Y133_BQ;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_C4 = CLBLM_L_X70Y123_SLICE_X104Y123_A5Q;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_C5 = CLBLM_L_X70Y123_SLICE_X104Y123_AQ;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_C6 = CLBLL_R_X71Y126_SLICE_X107Y126_BQ;
  assign CLBLM_L_X74Y134_SLICE_X112Y134_C3 = CLBLM_L_X74Y134_SLICE_X112Y134_DQ;
  assign CLBLM_L_X74Y134_SLICE_X112Y134_C4 = CLBLL_R_X75Y133_SLICE_X114Y133_BQ;
  assign CLBLM_L_X74Y134_SLICE_X112Y134_C5 = CLBLM_L_X74Y134_SLICE_X112Y134_BQ;
  assign CLBLM_L_X74Y134_SLICE_X112Y134_C6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y134_SLICE_X112Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y109_SLICE_X113Y109_A1 = CLBLM_L_X72Y109_SLICE_X109Y109_DQ;
  assign CLBLM_L_X74Y109_SLICE_X113Y109_A2 = CLBLL_R_X73Y109_SLICE_X110Y109_AQ;
  assign CLBLM_L_X74Y109_SLICE_X113Y109_A3 = CLBLM_L_X74Y109_SLICE_X113Y109_AQ;
  assign CLBLM_L_X74Y109_SLICE_X113Y109_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y109_SLICE_X113Y109_A5 = CLBLL_R_X75Y113_SLICE_X114Y113_AQ;
  assign CLBLM_L_X74Y109_SLICE_X113Y109_A6 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X113Y109_B1 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X111Y131_B1 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X113Y109_B2 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X113Y109_B3 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X113Y109_B4 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X113Y109_B5 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X111Y131_B2 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X113Y109_B6 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X113Y109_C1 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X111Y131_B3 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X113Y109_C2 = 1'b1;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_D5 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X113Y109_C3 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X113Y109_C4 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X111Y131_B4 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X113Y109_C5 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X113Y109_C6 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X113Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOB33_X105Y91_IOB_X1Y91_O = CLBLM_L_X68Y98_SLICE_X103Y98_AQ;
  assign CLBLL_R_X73Y131_SLICE_X111Y131_B5 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X113Y109_D1 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X111Y131_B6 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X113Y109_D2 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X113Y109_D3 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X113Y109_D4 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X113Y109_D5 = 1'b1;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_A5 = CLBLL_R_X73Y124_SLICE_X110Y124_AQ;
  assign CLBLM_L_X74Y109_SLICE_X113Y109_D6 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X113Y109_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign RIOI3_X105Y83_OLOGIC_X1Y83_D1 = CLBLM_R_X63Y105_SLICE_X95Y105_AQ;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_A6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_D6 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X112Y109_A1 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X112Y109_A2 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X112Y109_A3 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X112Y109_A4 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X112Y109_A5 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X112Y109_A6 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X112Y109_B1 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X112Y109_B2 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X111Y131_C1 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X112Y109_B3 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X112Y109_B4 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X112Y109_B5 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X112Y109_B6 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X111Y131_C2 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X112Y109_C1 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X111Y131_C3 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X112Y109_C2 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X112Y109_C3 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X112Y109_C4 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X112Y109_C5 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X111Y131_C4 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X112Y109_C6 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X111Y131_C5 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X111Y131_C6 = 1'b1;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_B3 = CLBLM_L_X70Y124_SLICE_X104Y124_AQ;
  assign CLBLM_L_X74Y109_SLICE_X112Y109_D1 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X112Y109_D2 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X112Y109_D3 = 1'b1;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_B4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y109_SLICE_X112Y109_D4 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X112Y109_D5 = 1'b1;
  assign CLBLM_L_X74Y109_SLICE_X112Y109_D6 = 1'b1;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_B5 = 1'b1;
  assign CLBLL_R_X73Y131_SLICE_X111Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_B6 = CLBLM_L_X70Y126_SLICE_X104Y126_CQ;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_T1 = 1'b1;
  assign LIOB33_X0Y77_IOB_X0Y78_O = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_C3 = CLBLM_L_X70Y124_SLICE_X104Y124_AQ;
  assign LIOB33_X0Y77_IOB_X0Y77_O = CLBLM_L_X60Y97_SLICE_X90Y97_BQ;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_C4 = CLBLM_L_X72Y122_SLICE_X109Y122_BQ;
  assign LIOB33_X0Y137_IOB_X0Y137_O = 1'b1;
  assign LIOB33_X0Y137_IOB_X0Y138_O = 1'b1;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_C5 = CLBLM_L_X70Y125_SLICE_X105Y125_AO5;
  assign LIOI3_X0Y89_OLOGIC_X0Y90_D1 = CLBLM_R_X63Y103_SLICE_X94Y103_AQ;
  assign LIOI3_X0Y89_OLOGIC_X0Y90_T1 = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_D1 = CLBLL_R_X83Y130_SLICE_X130Y130_BQ;
  assign LIOI3_X0Y89_OLOGIC_X0Y89_D1 = CLBLM_R_X63Y98_SLICE_X94Y98_BQ;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_T1 = 1'b1;
  assign LIOI3_X0Y89_OLOGIC_X0Y89_T1 = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_D1 = CLBLL_R_X83Y130_SLICE_X130Y130_AQ;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_T1 = 1'b1;
  assign LIOB33_X0Y125_IOB_X0Y126_O = CLBLL_L_X2Y131_SLICE_X0Y131_AO6;
  assign LIOB33_X0Y125_IOB_X0Y125_O = 1'b1;
  assign RIOB33_X105Y107_IOB_X1Y108_O = CLBLL_R_X77Y113_SLICE_X118Y113_AQ;
  assign RIOB33_X105Y107_IOB_X1Y107_O = CLBLM_R_X103Y69_SLICE_X162Y69_AQ;
  assign CLBLM_L_X76Y118_SLICE_X117Y118_A1 = CLBLM_L_X76Y123_SLICE_X117Y123_DO6;
  assign CLBLM_L_X76Y118_SLICE_X117Y118_A2 = CLBLM_L_X76Y118_SLICE_X117Y118_BQ;
  assign CLBLM_L_X76Y118_SLICE_X117Y118_A3 = CLBLM_L_X76Y118_SLICE_X117Y118_AQ;
  assign CLBLM_L_X76Y118_SLICE_X117Y118_A4 = 1'b1;
  assign CLBLM_L_X76Y118_SLICE_X117Y118_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X76Y118_SLICE_X117Y118_A6 = CLBLM_L_X76Y118_SLICE_X116Y118_CQ;
  assign CLBLM_L_X76Y118_SLICE_X117Y118_B1 = CLBLM_L_X76Y123_SLICE_X117Y123_DO6;
  assign CLBLM_L_X76Y118_SLICE_X117Y118_B2 = CLBLM_L_X76Y118_SLICE_X117Y118_BQ;
  assign CLBLM_L_X76Y118_SLICE_X117Y118_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X76Y118_SLICE_X117Y118_B4 = 1'b1;
  assign CLBLM_L_X76Y118_SLICE_X117Y118_B5 = CLBLM_L_X74Y123_SLICE_X113Y123_CO5;
  assign CLBLM_L_X76Y118_SLICE_X117Y118_B6 = CLBLM_L_X76Y118_SLICE_X116Y118_CQ;
  assign CLBLM_L_X76Y118_SLICE_X117Y118_C1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X76Y118_SLICE_X117Y118_C2 = CLBLM_L_X76Y118_SLICE_X116Y118_A5Q;
  assign CLBLM_L_X76Y118_SLICE_X117Y118_C3 = CLBLL_R_X77Y123_SLICE_X118Y123_DO6;
  assign CLBLM_L_X76Y118_SLICE_X117Y118_C4 = 1'b1;
  assign CLBLM_L_X76Y118_SLICE_X117Y118_C5 = CLBLM_L_X76Y118_SLICE_X117Y118_CQ;
  assign CLBLM_L_X76Y118_SLICE_X117Y118_C6 = CLBLM_L_X76Y118_SLICE_X116Y118_BQ;
  assign CLBLM_L_X76Y118_SLICE_X117Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X76Y118_SLICE_X117Y118_D1 = 1'b1;
  assign CLBLM_L_X76Y118_SLICE_X117Y118_D2 = 1'b1;
  assign CLBLM_L_X76Y118_SLICE_X117Y118_D3 = 1'b1;
  assign CLBLM_L_X76Y118_SLICE_X117Y118_D4 = 1'b1;
  assign CLBLM_L_X76Y118_SLICE_X117Y118_D5 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X105Y98_A1 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X105Y98_A2 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X105Y98_A3 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X105Y98_A4 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X105Y98_A5 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X105Y98_A6 = 1'b1;
  assign CLBLM_L_X76Y118_SLICE_X117Y118_D6 = 1'b1;
  assign CLBLM_L_X76Y118_SLICE_X116Y118_A1 = CLBLM_L_X76Y123_SLICE_X117Y123_DO6;
  assign CLBLM_L_X70Y98_SLICE_X105Y98_B1 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X105Y98_B2 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X105Y98_B3 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X105Y98_B4 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X105Y98_B5 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X105Y98_B6 = 1'b1;
  assign CLBLM_L_X76Y118_SLICE_X116Y118_A2 = 1'b1;
  assign CLBLM_L_X76Y118_SLICE_X116Y118_A3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X76Y118_SLICE_X116Y118_A4 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X105Y98_C1 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X105Y98_C2 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X105Y98_C3 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X105Y98_C4 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X105Y98_C5 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X105Y98_C6 = 1'b1;
  assign CLBLM_L_X76Y118_SLICE_X116Y118_AX = CLBLM_L_X76Y118_SLICE_X116Y118_BQ;
  assign CLBLM_L_X76Y118_SLICE_X116Y118_B1 = CLBLM_L_X76Y119_SLICE_X116Y119_A5Q;
  assign CLBLM_L_X76Y118_SLICE_X116Y118_B2 = CLBLM_L_X76Y118_SLICE_X116Y118_BQ;
  assign CLBLM_L_X76Y118_SLICE_X116Y118_B3 = CLBLM_L_X76Y118_SLICE_X116Y118_CQ;
  assign CLBLM_L_X76Y118_SLICE_X116Y118_B4 = CLBLM_L_X76Y118_SLICE_X117Y118_BQ;
  assign CLBLM_L_X76Y118_SLICE_X116Y118_B5 = CLBLM_L_X76Y118_SLICE_X117Y118_AQ;
  assign CLBLM_L_X76Y118_SLICE_X116Y118_B6 = CLBLM_L_X76Y118_SLICE_X116Y118_A5Q;
  assign CLBLM_L_X76Y118_SLICE_X116Y118_BX = CLBLM_L_X76Y118_SLICE_X116Y118_DQ;
  assign CLBLM_L_X70Y98_SLICE_X105Y98_D1 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X105Y98_D2 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X105Y98_D3 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X105Y98_D4 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X105Y98_D5 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X105Y98_D6 = 1'b1;
  assign CLBLM_L_X76Y118_SLICE_X116Y118_C3 = 1'b1;
  assign CLBLM_L_X76Y118_SLICE_X116Y118_C4 = 1'b1;
  assign CLBLM_L_X76Y118_SLICE_X116Y118_C6 = 1'b1;
  assign CLBLM_L_X76Y118_SLICE_X116Y118_CE = CLBLM_L_X76Y118_SLICE_X116Y118_AO6;
  assign CLBLM_L_X76Y118_SLICE_X116Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X76Y118_SLICE_X116Y118_CX = CLBLM_L_X76Y119_SLICE_X116Y119_A5Q;
  assign CLBLM_L_X70Y98_SLICE_X104Y98_A1 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X104Y98_A2 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X104Y98_A3 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X104Y98_A4 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X104Y98_A5 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X104Y98_A6 = 1'b1;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_D3 = 1'b1;
  assign CLBLM_L_X76Y118_SLICE_X116Y118_D1 = 1'b1;
  assign CLBLM_L_X76Y118_SLICE_X116Y118_D2 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X104Y98_AX = CLBLM_L_X70Y99_SLICE_X104Y99_AQ;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_D4 = CLBLL_R_X73Y119_SLICE_X110Y119_B5Q;
  assign CLBLM_L_X70Y98_SLICE_X104Y98_B1 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X104Y98_B2 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X104Y98_B3 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X104Y98_B4 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X104Y98_B5 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X104Y98_B6 = 1'b1;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_D5 = CLBLL_R_X73Y119_SLICE_X110Y119_CO6;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_D6 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X104Y98_C1 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X104Y98_C2 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X104Y98_C3 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X104Y98_C4 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X104Y98_C5 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X104Y98_C6 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X104Y98_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X70Y98_SLICE_X104Y98_D1 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X104Y98_D2 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X104Y98_D3 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X104Y98_D4 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X104Y98_D5 = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X104Y98_D6 = 1'b1;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign LIOB33_X0Y139_IOB_X0Y139_O = 1'b1;
  assign LIOB33_X0Y139_IOB_X0Y140_O = 1'b1;
  assign CLBLM_L_X70Y98_SLICE_X104Y98_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_A1 = CLBLM_L_X72Y119_SLICE_X108Y119_DO6;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_A2 = CLBLM_L_X72Y119_SLICE_X108Y119_BQ;
  assign RIOI3_X105Y145_OLOGIC_X1Y146_T1 = 1'b1;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_A3 = CLBLM_L_X72Y119_SLICE_X109Y119_A5Q;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_A4 = CLBLL_R_X71Y124_SLICE_X106Y124_BQ;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_A6 = 1'b1;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_B1 = 1'b1;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_B2 = CLBLM_L_X72Y119_SLICE_X109Y119_B5Q;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_B3 = CLBLM_L_X72Y119_SLICE_X109Y119_CO6;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_D1 = CLBLL_R_X75Y107_SLICE_X114Y107_AQ;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_B4 = CLBLL_R_X73Y118_SLICE_X111Y118_A5Q;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_B6 = CLBLM_L_X72Y119_SLICE_X108Y119_A5Q;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_C1 = CLBLM_L_X72Y119_SLICE_X109Y119_AQ;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_C2 = CLBLM_L_X70Y119_SLICE_X105Y119_A5Q;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_C3 = CLBLM_L_X68Y101_SLICE_X102Y101_BQ;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_C4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_T1 = 1'b1;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_T1 = 1'b1;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_C5 = CLBLM_L_X72Y119_SLICE_X108Y119_DO6;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_C6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1 = 1'b1;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X68Y109_SLICE_X103Y109_D3 = 1'b1;
  assign CLBLM_L_X76Y119_SLICE_X117Y119_A1 = 1'b1;
  assign CLBLM_L_X68Y109_SLICE_X103Y109_D4 = 1'b1;
  assign CLBLM_L_X76Y119_SLICE_X117Y119_A2 = 1'b1;
  assign CLBLM_L_X76Y119_SLICE_X117Y119_A3 = 1'b1;
  assign CLBLM_L_X76Y119_SLICE_X117Y119_A4 = 1'b1;
  assign CLBLM_L_X76Y119_SLICE_X117Y119_A5 = 1'b1;
  assign CLBLM_L_X68Y109_SLICE_X103Y109_D5 = 1'b1;
  assign CLBLM_L_X76Y119_SLICE_X117Y119_A6 = 1'b1;
  assign CLBLM_L_X76Y119_SLICE_X117Y119_B1 = 1'b1;
  assign CLBLM_L_X68Y109_SLICE_X103Y109_D6 = 1'b1;
  assign CLBLM_L_X76Y119_SLICE_X117Y119_B2 = 1'b1;
  assign CLBLM_L_X76Y119_SLICE_X117Y119_B3 = 1'b1;
  assign CLBLM_L_X76Y119_SLICE_X117Y119_B4 = 1'b1;
  assign CLBLM_L_X76Y119_SLICE_X117Y119_B5 = 1'b1;
  assign CLBLM_L_X76Y119_SLICE_X117Y119_B6 = 1'b1;
  assign CLBLM_L_X76Y119_SLICE_X117Y119_C1 = 1'b1;
  assign CLBLM_L_X76Y119_SLICE_X117Y119_C2 = 1'b1;
  assign CLBLM_L_X76Y119_SLICE_X117Y119_C3 = 1'b1;
  assign CLBLM_L_X76Y119_SLICE_X117Y119_C4 = 1'b1;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_D1 = CLBLM_L_X72Y119_SLICE_X109Y119_A5Q;
  assign CLBLM_L_X76Y119_SLICE_X117Y119_C5 = 1'b1;
  assign CLBLM_L_X76Y119_SLICE_X117Y119_C6 = 1'b1;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_D2 = CLBLM_L_X72Y119_SLICE_X108Y119_CQ;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_D3 = CLBLM_L_X72Y119_SLICE_X109Y119_B5Q;
  assign CLBLM_L_X76Y119_SLICE_X117Y119_D1 = 1'b1;
  assign CLBLM_L_X76Y119_SLICE_X117Y119_D2 = 1'b1;
  assign CLBLM_L_X76Y119_SLICE_X117Y119_D3 = 1'b1;
  assign CLBLM_L_X76Y119_SLICE_X117Y119_D4 = 1'b1;
  assign CLBLM_L_X70Y99_SLICE_X105Y99_A1 = CLBLM_L_X70Y100_SLICE_X105Y100_A5Q;
  assign CLBLM_L_X70Y99_SLICE_X105Y99_A2 = CLBLM_L_X70Y99_SLICE_X105Y99_BQ;
  assign CLBLM_L_X70Y99_SLICE_X105Y99_A3 = CLBLL_R_X71Y98_SLICE_X106Y98_A5Q;
  assign CLBLM_L_X70Y99_SLICE_X105Y99_A4 = CLBLM_L_X70Y101_SLICE_X105Y101_AQ;
  assign CLBLM_L_X70Y99_SLICE_X105Y99_A5 = CLBLM_L_X70Y100_SLICE_X105Y100_AQ;
  assign CLBLM_L_X70Y99_SLICE_X105Y99_A6 = 1'b1;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_D4 = CLBLM_L_X70Y119_SLICE_X105Y119_A5Q;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_D5 = CLBLM_L_X72Y119_SLICE_X109Y119_BQ;
  assign CLBLM_L_X76Y119_SLICE_X116Y119_A1 = CLBLM_L_X76Y123_SLICE_X117Y123_DO6;
  assign CLBLM_L_X70Y99_SLICE_X105Y99_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y99_SLICE_X105Y99_B2 = CLBLM_L_X70Y99_SLICE_X105Y99_BQ;
  assign CLBLM_L_X70Y99_SLICE_X105Y99_B3 = CLBLM_L_X70Y103_SLICE_X105Y103_CO6;
  assign CLBLM_L_X70Y99_SLICE_X105Y99_B4 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X70Y99_SLICE_X105Y99_B5 = CLBLM_L_X70Y103_SLICE_X105Y103_DO6;
  assign CLBLM_L_X70Y99_SLICE_X105Y99_B6 = CLBLM_L_X70Y100_SLICE_X104Y100_CQ;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_D6 = CLBLL_R_X73Y118_SLICE_X111Y118_A5Q;
  assign CLBLM_L_X76Y119_SLICE_X116Y119_A2 = CLBLM_L_X74Y117_SLICE_X112Y117_BQ;
  assign CLBLM_L_X76Y119_SLICE_X116Y119_A3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y99_SLICE_X105Y99_C1 = CLBLM_L_X70Y103_SLICE_X105Y103_CO6;
  assign CLBLM_L_X70Y99_SLICE_X105Y99_C2 = CLBLM_L_X70Y99_SLICE_X105Y99_CQ;
  assign CLBLM_L_X70Y99_SLICE_X105Y99_C3 = CLBLM_L_X70Y99_SLICE_X105Y99_BQ;
  assign CLBLM_L_X70Y99_SLICE_X105Y99_C4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y99_SLICE_X105Y99_C5 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X70Y99_SLICE_X105Y99_C6 = CLBLM_L_X70Y103_SLICE_X105Y103_DO5;
  assign CLBLM_L_X76Y119_SLICE_X116Y119_B1 = CLBLM_L_X76Y118_SLICE_X116Y118_AQ;
  assign CLBLM_L_X70Y99_SLICE_X105Y99_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X76Y119_SLICE_X116Y119_B2 = CLBLM_L_X76Y118_SLICE_X116Y118_BO6;
  assign CLBLM_L_X76Y119_SLICE_X116Y119_B4 = CLBLM_L_X76Y118_SLICE_X116Y118_DQ;
  assign CLBLM_L_X76Y119_SLICE_X116Y119_B5 = 1'b1;
  assign CLBLM_L_X70Y99_SLICE_X105Y99_D1 = 1'b1;
  assign CLBLM_L_X70Y99_SLICE_X105Y99_D2 = 1'b1;
  assign CLBLM_L_X68Y109_SLICE_X102Y109_A6 = 1'b1;
  assign CLBLM_L_X70Y99_SLICE_X105Y99_D3 = 1'b1;
  assign CLBLM_L_X70Y99_SLICE_X105Y99_D4 = 1'b1;
  assign CLBLM_L_X70Y99_SLICE_X105Y99_D5 = 1'b1;
  assign CLBLM_L_X70Y99_SLICE_X105Y99_D6 = 1'b1;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X70Y99_SLICE_X105Y99_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X76Y119_SLICE_X116Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X76Y119_SLICE_X116Y119_D1 = 1'b1;
  assign CLBLM_L_X70Y99_SLICE_X104Y99_A1 = CLBLM_L_X70Y101_SLICE_X104Y101_BQ;
  assign CLBLM_L_X70Y99_SLICE_X104Y99_A2 = CLBLM_L_X70Y100_SLICE_X105Y100_A5Q;
  assign CLBLM_L_X70Y99_SLICE_X104Y99_A3 = CLBLM_L_X70Y99_SLICE_X104Y99_AQ;
  assign CLBLM_L_X70Y99_SLICE_X104Y99_A4 = CLBLM_L_X60Y97_SLICE_X90Y97_BQ;
  assign CLBLM_L_X70Y99_SLICE_X104Y99_A5 = CLBLM_L_X70Y100_SLICE_X105Y100_AQ;
  assign CLBLM_L_X70Y99_SLICE_X104Y99_A6 = CLBLM_L_X70Y99_SLICE_X105Y99_CQ;
  assign CLBLM_L_X76Y119_SLICE_X116Y119_D2 = 1'b1;
  assign CLBLM_L_X76Y119_SLICE_X116Y119_D3 = 1'b1;
  assign CLBLM_L_X76Y119_SLICE_X116Y119_D4 = 1'b1;
  assign CLBLM_L_X70Y99_SLICE_X104Y99_AX = CLBLM_L_X70Y101_SLICE_X105Y101_AQ;
  assign CLBLL_R_X79Y104_SLICE_X122Y104_A3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y99_SLICE_X104Y99_B1 = CLBLM_L_X70Y100_SLICE_X104Y100_CQ;
  assign CLBLM_L_X70Y99_SLICE_X104Y99_B2 = CLBLM_L_X70Y101_SLICE_X104Y101_CQ;
  assign CLBLM_L_X70Y99_SLICE_X104Y99_B3 = CLBLM_L_X70Y101_SLICE_X104Y101_AQ;
  assign CLBLM_L_X70Y99_SLICE_X104Y99_B4 = CLBLL_R_X71Y100_SLICE_X106Y100_BQ;
  assign CLBLM_L_X70Y99_SLICE_X104Y99_B5 = CLBLM_L_X70Y100_SLICE_X105Y100_AQ;
  assign CLBLM_L_X70Y99_SLICE_X104Y99_B6 = CLBLM_L_X70Y100_SLICE_X105Y100_A5Q;
  assign CLBLM_L_X76Y119_SLICE_X116Y119_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_R_X67Y108_SLICE_X100Y108_A5 = CLBLM_R_X67Y108_SLICE_X100Y108_C5Q;
  assign LIOB33_X0Y141_IOB_X0Y141_O = 1'b1;
  assign LIOB33_X0Y141_IOB_X0Y142_O = 1'b1;
  assign CLBLM_L_X70Y99_SLICE_X104Y99_C1 = CLBLM_L_X70Y99_SLICE_X104Y99_AO6;
  assign CLBLM_L_X70Y99_SLICE_X104Y99_C2 = CLBLM_L_X70Y99_SLICE_X105Y99_AO6;
  assign CLBLM_L_X70Y99_SLICE_X104Y99_C3 = CLBLM_L_X70Y100_SLICE_X104Y100_DO6;
  assign CLBLM_L_X70Y99_SLICE_X104Y99_C4 = CLBLL_R_X71Y101_SLICE_X106Y101_DO6;
  assign CLBLM_L_X70Y99_SLICE_X104Y99_C5 = CLBLM_L_X70Y99_SLICE_X104Y99_DO6;
  assign CLBLM_L_X70Y99_SLICE_X104Y99_C6 = CLBLM_L_X70Y99_SLICE_X104Y99_BO6;
  assign CLBLM_L_X70Y99_SLICE_X104Y99_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X68Y109_SLICE_X102Y109_B4 = CLBLM_R_X65Y109_SLICE_X99Y109_A5Q;
  assign CLBLM_R_X67Y108_SLICE_X100Y108_A6 = 1'b1;
  assign CLBLM_L_X70Y99_SLICE_X104Y99_D1 = CLBLM_L_X70Y100_SLICE_X105Y100_AQ;
  assign CLBLM_L_X68Y109_SLICE_X102Y109_B5 = CLBLM_L_X68Y109_SLICE_X102Y109_A5Q;
  assign CLBLM_L_X70Y99_SLICE_X104Y99_D2 = 1'b1;
  assign CLBLM_L_X70Y99_SLICE_X104Y99_D3 = CLBLM_L_X70Y99_SLICE_X104Y99_AQ;
  assign CLBLM_L_X70Y99_SLICE_X104Y99_D4 = CLBLM_L_X70Y100_SLICE_X105Y100_A5Q;
  assign CLBLM_L_X70Y99_SLICE_X104Y99_D5 = CLBLM_L_X70Y102_SLICE_X105Y102_CQ;
  assign CLBLM_L_X68Y109_SLICE_X102Y109_B6 = 1'b1;
  assign CLBLM_L_X70Y99_SLICE_X104Y99_D6 = CLBLL_R_X71Y98_SLICE_X106Y98_A5Q;
  assign CLBLM_L_X70Y99_SLICE_X104Y99_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X79Y104_SLICE_X122Y104_B2 = CLBLL_R_X75Y124_SLICE_X115Y124_BQ;
  assign CLBLM_L_X78Y131_SLICE_X120Y131_C2 = 1'b1;
  assign CLBLM_L_X68Y109_SLICE_X102Y109_C6 = CLBLM_R_X67Y109_SLICE_X101Y109_DO6;
  assign CLBLL_R_X79Y104_SLICE_X122Y104_C2 = 1'b1;
  assign CLBLL_R_X79Y104_SLICE_X122Y104_C3 = 1'b1;
  assign CLBLM_L_X68Y109_SLICE_X102Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X68Y109_SLICE_X102Y109_D1 = CLBLM_R_X67Y110_SLICE_X101Y110_AQ;
  assign CLBLM_L_X68Y109_SLICE_X102Y109_D2 = CLBLM_L_X68Y109_SLICE_X102Y109_BO6;
  assign CLBLM_L_X68Y109_SLICE_X102Y109_D3 = CLBLM_R_X67Y110_SLICE_X101Y110_DQ;
  assign CLBLM_L_X82Y98_SLICE_X129Y98_A1 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X129Y98_A2 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X129Y98_A3 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X129Y98_A4 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X129Y98_A5 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X129Y98_A6 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X129Y98_B1 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X129Y98_B2 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X129Y98_B3 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X129Y98_B4 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X129Y98_B5 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X129Y98_B6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X129Y98_C1 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X129Y98_C2 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X129Y98_C3 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X129Y98_C4 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X129Y98_C5 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X129Y98_C6 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X129Y98_D1 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X129Y98_D2 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X129Y98_D3 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X129Y98_D4 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X129Y98_D5 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X129Y98_D6 = 1'b1;
  assign LIOI3_X0Y91_OLOGIC_X0Y92_D1 = CLBLM_L_X62Y95_SLICE_X92Y95_CQ;
  assign CLBLM_L_X82Y98_SLICE_X128Y98_A1 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X128Y98_A2 = CLBLM_L_X82Y98_SLICE_X128Y98_BQ;
  assign CLBLM_L_X82Y98_SLICE_X128Y98_A3 = CLBLM_L_X82Y98_SLICE_X128Y98_AQ;
  assign CLBLM_L_X82Y98_SLICE_X128Y98_A4 = CLBLL_R_X77Y104_SLICE_X118Y104_AQ;
  assign CLBLM_L_X82Y98_SLICE_X128Y98_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X82Y98_SLICE_X128Y98_A6 = 1'b1;
  assign LIOI3_X0Y91_OLOGIC_X0Y92_T1 = 1'b1;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_D1 = CLBLL_R_X83Y130_SLICE_X130Y130_DQ;
  assign CLBLM_L_X82Y98_SLICE_X128Y98_B1 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X128Y98_B2 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X128Y98_B3 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X128Y98_B4 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X128Y98_B5 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X128Y98_B6 = 1'b1;
  assign LIOI3_X0Y91_OLOGIC_X0Y91_D1 = CLBLM_L_X60Y99_SLICE_X90Y99_DQ;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_T1 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X128Y98_BX = CLBLM_L_X82Y98_SLICE_X128Y98_AQ;
  assign CLBLM_L_X82Y98_SLICE_X128Y98_C1 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X128Y98_C2 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X128Y98_C3 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X128Y98_C4 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X128Y98_C5 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X128Y98_C6 = 1'b1;
  assign LIOI3_X0Y91_OLOGIC_X0Y91_T1 = 1'b1;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_D1 = CLBLL_R_X83Y130_SLICE_X130Y130_CQ;
  assign CLBLM_L_X82Y98_SLICE_X128Y98_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X82Y98_SLICE_X128Y98_D1 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X128Y98_D2 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X128Y98_D3 = 1'b1;
  assign CLBLM_L_X82Y98_SLICE_X128Y98_D4 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_A1 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_A2 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_A3 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_A4 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_A5 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_A6 = 1'b1;
  assign CLBLM_L_X70Y100_SLICE_X105Y100_A1 = CLBLM_L_X70Y100_SLICE_X105Y100_B5Q;
  assign CLBLM_L_X70Y100_SLICE_X105Y100_A2 = CLBLM_R_X65Y103_SLICE_X99Y103_DO6;
  assign CLBLM_L_X70Y100_SLICE_X105Y100_A3 = CLBLM_L_X70Y100_SLICE_X105Y100_AQ;
  assign CLBLM_L_X70Y100_SLICE_X105Y100_A4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y100_SLICE_X105Y100_A5 = CLBLM_L_X70Y100_SLICE_X105Y100_A5Q;
  assign CLBLM_L_X70Y100_SLICE_X105Y100_A6 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_AX = CLBLM_L_X72Y111_SLICE_X108Y111_C5Q;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_B1 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_B5 = 1'b1;
  assign CLBLM_L_X70Y100_SLICE_X105Y100_B1 = CLBLM_L_X70Y100_SLICE_X105Y100_B5Q;
  assign CLBLM_L_X70Y100_SLICE_X105Y100_B2 = CLBLM_L_X70Y100_SLICE_X105Y100_BQ;
  assign CLBLM_L_X70Y100_SLICE_X105Y100_B3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y100_SLICE_X105Y100_B4 = CLBLL_R_X71Y100_SLICE_X106Y100_AO5;
  assign CLBLM_L_X70Y100_SLICE_X105Y100_B5 = CLBLL_R_X71Y98_SLICE_X106Y98_A5Q;
  assign CLBLM_L_X70Y100_SLICE_X105Y100_B6 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_B6 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_C1 = 1'b1;
  assign CLBLM_L_X70Y100_SLICE_X105Y100_C1 = CLBLM_L_X60Y99_SLICE_X90Y99_AQ;
  assign CLBLM_L_X70Y100_SLICE_X105Y100_C2 = CLBLL_R_X77Y108_SLICE_X118Y108_AQ;
  assign CLBLM_L_X70Y100_SLICE_X105Y100_C3 = CLBLL_R_X71Y101_SLICE_X106Y101_AQ;
  assign CLBLM_L_X70Y100_SLICE_X105Y100_C4 = CLBLM_L_X70Y100_SLICE_X105Y100_A5Q;
  assign CLBLM_L_X70Y100_SLICE_X105Y100_C5 = CLBLM_L_X70Y101_SLICE_X105Y101_BQ;
  assign CLBLM_L_X70Y100_SLICE_X105Y100_C6 = CLBLM_L_X70Y100_SLICE_X105Y100_AQ;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_C4 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_C5 = 1'b1;
  assign CLBLM_L_X70Y100_SLICE_X105Y100_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_D1 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_D2 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_D3 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_D4 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_D5 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_D6 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X70Y100_SLICE_X105Y100_CX = CLBLL_R_X77Y108_SLICE_X118Y108_AQ;
  assign CLBLM_L_X70Y100_SLICE_X105Y100_D1 = CLBLM_L_X70Y101_SLICE_X104Y101_AO6;
  assign CLBLM_L_X70Y100_SLICE_X105Y100_D2 = CLBLM_L_X70Y100_SLICE_X105Y100_CQ;
  assign CLBLM_L_X70Y100_SLICE_X105Y100_D3 = CLBLL_R_X71Y100_SLICE_X106Y100_AO6;
  assign CLBLM_L_X70Y100_SLICE_X105Y100_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X70Y100_SLICE_X105Y100_D4 = CLBLM_L_X70Y100_SLICE_X105Y100_CO6;
  assign CLBLM_L_X70Y100_SLICE_X105Y100_D5 = CLBLL_R_X71Y100_SLICE_X106Y100_CO6;
  assign CLBLM_L_X70Y100_SLICE_X105Y100_D6 = CLBLL_R_X71Y101_SLICE_X107Y101_AQ;
  assign CLBLM_L_X70Y100_SLICE_X104Y100_A1 = CLBLM_L_X70Y103_SLICE_X105Y103_CO6;
  assign CLBLM_L_X70Y100_SLICE_X104Y100_A2 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y100_SLICE_X104Y100_A3 = CLBLM_L_X70Y100_SLICE_X104Y100_AQ;
  assign CLBLM_L_X70Y100_SLICE_X104Y100_A4 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X70Y100_SLICE_X104Y100_A5 = CLBLM_L_X70Y101_SLICE_X104Y101_BQ;
  assign CLBLM_L_X70Y100_SLICE_X104Y100_A6 = CLBLM_L_X70Y103_SLICE_X104Y103_DO6;
  assign CLBLM_L_X70Y100_SLICE_X104Y100_AX = CLBLM_L_X60Y97_SLICE_X90Y97_BQ;
  assign CLBLM_L_X70Y100_SLICE_X104Y100_B1 = CLBLM_L_X70Y103_SLICE_X105Y103_CO6;
  assign CLBLM_L_X70Y100_SLICE_X104Y100_B2 = CLBLM_L_X70Y100_SLICE_X104Y100_BQ;
  assign CLBLM_L_X70Y100_SLICE_X104Y100_B3 = CLBLM_L_X70Y103_SLICE_X104Y103_C5Q;
  assign CLBLM_L_X70Y100_SLICE_X104Y100_B4 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X70Y100_SLICE_X104Y100_B5 = CLBLM_L_X70Y99_SLICE_X105Y99_CQ;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_A1 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_A2 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_A3 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_A4 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_A5 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_A6 = 1'b1;
  assign CLBLM_L_X70Y100_SLICE_X104Y100_B6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y100_SLICE_X104Y100_C2 = CLBLM_L_X70Y100_SLICE_X104Y100_CQ;
  assign CLBLM_L_X70Y100_SLICE_X104Y100_C3 = CLBLM_L_X70Y100_SLICE_X104Y100_AQ;
  assign CLBLM_L_X70Y100_SLICE_X104Y100_C4 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y100_SLICE_X104Y100_C6 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X70Y100_SLICE_X104Y100_C1 = CLBLM_L_X70Y103_SLICE_X104Y103_DO5;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_B1 = 1'b1;
  assign CLBLM_L_X70Y100_SLICE_X104Y100_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_B2 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_B3 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_B4 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_B5 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_B6 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_C1 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_C2 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_C3 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_C4 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_C5 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_C6 = 1'b1;
  assign CLBLM_L_X70Y100_SLICE_X104Y100_D1 = CLBLM_L_X70Y100_SLICE_X104Y100_BQ;
  assign CLBLM_L_X70Y100_SLICE_X104Y100_D2 = CLBLM_L_X70Y100_SLICE_X104Y100_AQ;
  assign CLBLM_L_X70Y100_SLICE_X104Y100_D3 = CLBLM_L_X70Y98_SLICE_X104Y98_AQ;
  assign CLBLM_L_X70Y100_SLICE_X104Y100_D4 = CLBLM_L_X70Y100_SLICE_X104Y100_A5Q;
  assign CLBLM_L_X70Y100_SLICE_X104Y100_D5 = CLBLM_L_X70Y100_SLICE_X105Y100_AQ;
  assign CLBLM_L_X70Y100_SLICE_X104Y100_D6 = CLBLM_L_X70Y100_SLICE_X105Y100_A5Q;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_D1 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_D2 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_D3 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_D4 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_D5 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_D6 = 1'b1;
  assign CLBLM_L_X74Y135_SLICE_X113Y135_B6 = CLBLM_L_X74Y135_SLICE_X113Y135_BQ;
  assign CLBLM_L_X74Y135_SLICE_X113Y135_C1 = CLBLM_L_X74Y134_SLICE_X113Y134_A5Q;
  assign LIOB33_X0Y145_IOB_X0Y146_O = CLBLM_L_X72Y123_SLICE_X108Y123_BO6;
  assign CLBLM_L_X70Y101_SLICE_X105Y101_A1 = CLBLM_L_X70Y100_SLICE_X105Y100_A5Q;
  assign CLBLM_L_X70Y101_SLICE_X105Y101_A2 = CLBLL_R_X71Y98_SLICE_X106Y98_A5Q;
  assign CLBLM_L_X70Y101_SLICE_X105Y101_A3 = CLBLM_L_X70Y102_SLICE_X105Y102_AQ;
  assign CLBLM_L_X70Y101_SLICE_X105Y101_A4 = CLBLL_R_X71Y100_SLICE_X106Y100_BQ;
  assign CLBLM_L_X70Y101_SLICE_X105Y101_A5 = CLBLM_L_X70Y100_SLICE_X105Y100_AQ;
  assign CLBLM_L_X70Y101_SLICE_X105Y101_A6 = 1'b1;
  assign LIOB33_X0Y145_IOB_X0Y145_O = CLBLL_R_X71Y130_SLICE_X106Y130_DO6;
  assign CLBLM_L_X70Y101_SLICE_X105Y101_AX = CLBLM_L_X70Y101_SLICE_X104Y101_AQ;
  assign CLBLM_L_X70Y101_SLICE_X105Y101_B1 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X70Y101_SLICE_X105Y101_B2 = CLBLM_L_X70Y101_SLICE_X105Y101_BQ;
  assign CLBLM_L_X70Y101_SLICE_X105Y101_B3 = CLBLM_L_X70Y103_SLICE_X105Y103_CO5;
  assign CLBLM_L_X70Y101_SLICE_X105Y101_B4 = CLBLM_L_X70Y103_SLICE_X105Y103_DO5;
  assign CLBLM_L_X70Y101_SLICE_X105Y101_B5 = CLBLL_R_X71Y101_SLICE_X107Y101_AQ;
  assign CLBLM_L_X70Y101_SLICE_X105Y101_B6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y101_SLICE_X105Y101_C1 = CLBLM_L_X70Y100_SLICE_X105Y100_DO6;
  assign CLBLM_L_X70Y101_SLICE_X105Y101_C2 = CLBLM_L_X70Y99_SLICE_X104Y99_CO6;
  assign CLBLM_L_X70Y101_SLICE_X105Y101_C3 = CLBLL_R_X71Y102_SLICE_X106Y102_DO6;
  assign CLBLM_L_X70Y101_SLICE_X105Y101_C4 = CLBLM_L_X70Y99_SLICE_X105Y99_AO5;
  assign CLBLM_L_X70Y101_SLICE_X105Y101_C5 = CLBLM_L_X70Y101_SLICE_X105Y101_DO6;
  assign CLBLM_L_X70Y101_SLICE_X105Y101_C6 = CLBLM_R_X65Y103_SLICE_X99Y103_DO6;
  assign CLBLM_L_X70Y101_SLICE_X105Y101_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_D1 = 1'b1;
  assign CLBLM_L_X70Y101_SLICE_X105Y101_D1 = CLBLM_L_X70Y101_SLICE_X105Y101_AO6;
  assign CLBLM_L_X70Y101_SLICE_X105Y101_D2 = CLBLL_R_X71Y98_SLICE_X106Y98_A5Q;
  assign CLBLM_L_X70Y101_SLICE_X105Y101_D3 = CLBLM_L_X70Y98_SLICE_X104Y98_AQ;
  assign CLBLM_L_X70Y101_SLICE_X105Y101_D4 = CLBLM_L_X70Y101_SLICE_X105Y101_AO5;
  assign CLBLM_L_X70Y101_SLICE_X105Y101_D5 = CLBLM_L_X70Y102_SLICE_X105Y102_BQ;
  assign CLBLM_L_X70Y101_SLICE_X105Y101_D6 = CLBLM_L_X70Y102_SLICE_X104Y102_BO6;
  assign CLBLM_L_X74Y135_SLICE_X113Y135_D1 = CLBLM_L_X74Y134_SLICE_X113Y134_A5Q;
  assign CLBLM_L_X70Y101_SLICE_X105Y101_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y135_SLICE_X113Y135_D2 = CLBLL_R_X75Y134_SLICE_X115Y134_CO6;
  assign CLBLM_L_X70Y101_SLICE_X104Y101_A1 = CLBLM_L_X70Y100_SLICE_X105Y100_A5Q;
  assign CLBLM_L_X70Y101_SLICE_X104Y101_A2 = CLBLM_R_X65Y103_SLICE_X99Y103_DO6;
  assign CLBLM_L_X70Y101_SLICE_X104Y101_A3 = CLBLL_R_X71Y98_SLICE_X106Y98_A5Q;
  assign CLBLM_L_X70Y101_SLICE_X104Y101_A4 = CLBLM_L_X60Y97_SLICE_X90Y97_BQ;
  assign CLBLM_L_X70Y101_SLICE_X104Y101_A5 = CLBLM_L_X70Y100_SLICE_X105Y100_AQ;
  assign CLBLM_L_X70Y101_SLICE_X104Y101_A6 = 1'b1;
  assign CLBLM_L_X74Y135_SLICE_X113Y135_D3 = CLBLM_L_X74Y135_SLICE_X113Y135_BQ;
  assign CLBLM_L_X74Y135_SLICE_X113Y135_D4 = 1'b1;
  assign CLBLM_L_X70Y101_SLICE_X104Y101_AX = CLBLM_L_X70Y100_SLICE_X104Y100_A5Q;
  assign CLBLM_L_X74Y135_SLICE_X113Y135_D5 = CLBLM_L_X74Y134_SLICE_X113Y134_CQ;
  assign CLBLM_L_X70Y101_SLICE_X104Y101_B1 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y101_SLICE_X104Y101_B2 = CLBLM_L_X70Y101_SLICE_X104Y101_BQ;
  assign CLBLM_L_X70Y101_SLICE_X104Y101_B3 = CLBLM_L_X70Y103_SLICE_X104Y103_C5Q;
  assign CLBLM_L_X70Y101_SLICE_X104Y101_B4 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X70Y101_SLICE_X104Y101_B5 = CLBLL_R_X71Y103_SLICE_X106Y103_BO6;
  assign CLBLM_L_X70Y101_SLICE_X104Y101_B6 = CLBLL_R_X71Y101_SLICE_X106Y101_CQ;
  assign CLBLM_L_X74Y135_SLICE_X113Y135_D6 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y101_SLICE_X104Y101_C1 = CLBLM_L_X70Y103_SLICE_X105Y103_CO5;
  assign CLBLM_L_X70Y101_SLICE_X104Y101_C2 = CLBLM_L_X70Y101_SLICE_X104Y101_CQ;
  assign CLBLM_L_X70Y101_SLICE_X104Y101_C3 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X70Y101_SLICE_X104Y101_C4 = CLBLL_R_X79Y96_SLICE_X122Y96_AO6;
  assign CLBLM_L_X70Y101_SLICE_X104Y101_C5 = CLBLM_L_X70Y103_SLICE_X104Y103_DO6;
  assign CLBLM_L_X70Y101_SLICE_X104Y101_C6 = CLBLM_L_X70Y100_SLICE_X104Y100_BQ;
  assign CLBLM_L_X70Y101_SLICE_X104Y101_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y135_SLICE_X113Y135_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X70Y101_SLICE_X104Y101_D1 = CLBLM_L_X70Y100_SLICE_X105Y100_BQ;
  assign CLBLM_L_X70Y101_SLICE_X104Y101_D2 = CLBLM_L_X70Y100_SLICE_X105Y100_A5Q;
  assign CLBLM_L_X70Y101_SLICE_X104Y101_D3 = CLBLM_R_X65Y102_SLICE_X99Y102_AQ;
  assign CLBLM_L_X70Y101_SLICE_X104Y101_D4 = CLBLM_L_X70Y100_SLICE_X105Y100_B5Q;
  assign CLBLM_L_X70Y101_SLICE_X104Y101_D5 = CLBLM_L_X70Y100_SLICE_X105Y100_AQ;
  assign CLBLM_L_X70Y101_SLICE_X104Y101_D6 = CLBLM_R_X65Y103_SLICE_X99Y103_DO6;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_T1 = 1'b1;
  assign CLBLM_L_X70Y101_SLICE_X104Y101_SR = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLM_L_X74Y135_SLICE_X112Y135_A1 = CLBLM_L_X74Y135_SLICE_X113Y135_CO6;
  assign CLBLM_L_X74Y135_SLICE_X112Y135_A2 = CLBLM_L_X74Y135_SLICE_X113Y135_DO6;
  assign CLBLM_L_X74Y135_SLICE_X112Y135_A3 = CLBLM_L_X74Y135_SLICE_X112Y135_AQ;
  assign CLBLM_L_X74Y135_SLICE_X112Y135_A4 = CLBLM_L_X74Y135_SLICE_X113Y135_BQ;
  assign CLBLM_L_X74Y135_SLICE_X112Y135_A5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X74Y135_SLICE_X112Y135_A6 = 1'b1;
  assign RIOB33_SING_X105Y100_IOB_X1Y100_O = CLBLM_L_X78Y104_SLICE_X120Y104_A5Q;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_D1 = 1'b1;
  assign CLBLM_L_X74Y135_SLICE_X112Y135_B1 = CLBLM_L_X74Y132_SLICE_X112Y132_C5Q;
  assign CLBLM_L_X74Y135_SLICE_X112Y135_B2 = CLBLM_L_X74Y134_SLICE_X112Y134_CQ;
  assign CLBLM_L_X74Y135_SLICE_X112Y135_B3 = CLBLM_L_X74Y135_SLICE_X112Y135_AQ;
  assign CLBLM_L_X74Y135_SLICE_X112Y135_B4 = CLBLM_L_X74Y134_SLICE_X112Y134_BQ;
  assign CLBLM_L_X74Y135_SLICE_X112Y135_B5 = CLBLL_R_X73Y134_SLICE_X110Y134_AO6;
  assign CLBLM_L_X74Y135_SLICE_X112Y135_B6 = CLBLL_R_X75Y133_SLICE_X114Y133_BQ;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_T1 = 1'b1;
  assign CLBLM_L_X74Y135_SLICE_X112Y135_C1 = 1'b1;
  assign CLBLM_L_X74Y135_SLICE_X112Y135_C2 = 1'b1;
  assign CLBLM_L_X74Y135_SLICE_X112Y135_C3 = 1'b1;
  assign CLBLM_L_X74Y135_SLICE_X112Y135_C4 = 1'b1;
  assign CLBLM_L_X74Y135_SLICE_X112Y135_C5 = 1'b1;
  assign CLBLM_L_X74Y135_SLICE_X112Y135_C6 = 1'b1;
  assign CLBLM_R_X65Y110_SLICE_X98Y110_A5 = CLBLM_R_X67Y111_SLICE_X101Y111_B5Q;
  assign CLBLM_R_X65Y110_SLICE_X98Y110_A6 = CLBLM_R_X65Y110_SLICE_X99Y110_AO6;
  assign CLBLM_L_X74Y135_SLICE_X112Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
endmodule
