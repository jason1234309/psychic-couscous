
module b15_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24;
  wire   [8:2] carry;

  FADDX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FADDX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  FADDX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n23), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .IN1(B[28]), .IN2(n20), .Q(SUM[28]) );
  XOR2X1 U2 ( .IN1(B[27]), .IN2(n19), .Q(SUM[27]) );
  XOR2X1 U3 ( .IN1(B[26]), .IN2(n18), .Q(SUM[26]) );
  XOR2X1 U4 ( .IN1(B[25]), .IN2(n17), .Q(SUM[25]) );
  XOR2X1 U5 ( .IN1(B[24]), .IN2(n16), .Q(SUM[24]) );
  XOR2X1 U6 ( .IN1(B[23]), .IN2(n15), .Q(SUM[23]) );
  XOR2X1 U7 ( .IN1(B[22]), .IN2(n14), .Q(SUM[22]) );
  XOR2X1 U8 ( .IN1(B[21]), .IN2(n13), .Q(SUM[21]) );
  XOR2X1 U9 ( .IN1(B[20]), .IN2(n6), .Q(SUM[20]) );
  XOR2X1 U10 ( .IN1(B[29]), .IN2(n21), .Q(SUM[29]) );
  XOR2X1 U11 ( .IN1(B[30]), .IN2(n22), .Q(SUM[30]) );
  XNOR2X1 U12 ( .IN1(B[31]), .IN2(n24), .Q(SUM[31]) );
  NAND2X0 U13 ( .IN1(B[30]), .IN2(n22), .QN(n24) );
  AND2X1 U14 ( .IN1(B[10]), .IN2(n8), .Q(n1) );
  AND2X1 U15 ( .IN1(B[11]), .IN2(n1), .Q(n2) );
  AND2X1 U16 ( .IN1(B[14]), .IN2(n10), .Q(n3) );
  AND2X1 U17 ( .IN1(B[15]), .IN2(n3), .Q(n4) );
  AND2X1 U18 ( .IN1(B[18]), .IN2(n12), .Q(n5) );
  AND2X1 U19 ( .IN1(B[19]), .IN2(n5), .Q(n6) );
  XOR2X1 U20 ( .IN1(B[19]), .IN2(n5), .Q(SUM[19]) );
  XOR2X1 U21 ( .IN1(B[18]), .IN2(n12), .Q(SUM[18]) );
  AND2X1 U22 ( .IN1(B[8]), .IN2(carry[8]), .Q(n7) );
  AND2X1 U23 ( .IN1(B[9]), .IN2(n7), .Q(n8) );
  AND2X1 U24 ( .IN1(B[12]), .IN2(n2), .Q(n9) );
  AND2X1 U25 ( .IN1(B[13]), .IN2(n9), .Q(n10) );
  AND2X1 U26 ( .IN1(B[16]), .IN2(n4), .Q(n11) );
  AND2X1 U27 ( .IN1(B[17]), .IN2(n11), .Q(n12) );
  AND2X1 U28 ( .IN1(B[20]), .IN2(n6), .Q(n13) );
  AND2X1 U29 ( .IN1(B[21]), .IN2(n13), .Q(n14) );
  AND2X1 U30 ( .IN1(B[22]), .IN2(n14), .Q(n15) );
  AND2X1 U31 ( .IN1(B[23]), .IN2(n15), .Q(n16) );
  AND2X1 U32 ( .IN1(B[24]), .IN2(n16), .Q(n17) );
  AND2X1 U33 ( .IN1(B[25]), .IN2(n17), .Q(n18) );
  AND2X1 U34 ( .IN1(B[26]), .IN2(n18), .Q(n19) );
  AND2X1 U35 ( .IN1(B[27]), .IN2(n19), .Q(n20) );
  AND2X1 U36 ( .IN1(B[28]), .IN2(n20), .Q(n21) );
  AND2X1 U37 ( .IN1(B[29]), .IN2(n21), .Q(n22) );
  XOR2X1 U38 ( .IN1(B[17]), .IN2(n11), .Q(SUM[17]) );
  XOR2X1 U39 ( .IN1(B[16]), .IN2(n4), .Q(SUM[16]) );
  XOR2X1 U40 ( .IN1(B[15]), .IN2(n3), .Q(SUM[15]) );
  XOR2X1 U41 ( .IN1(B[14]), .IN2(n10), .Q(SUM[14]) );
  XOR2X1 U42 ( .IN1(B[13]), .IN2(n9), .Q(SUM[13]) );
  XOR2X1 U43 ( .IN1(B[12]), .IN2(n2), .Q(SUM[12]) );
  XOR2X1 U44 ( .IN1(B[11]), .IN2(n1), .Q(SUM[11]) );
  XOR2X1 U45 ( .IN1(B[10]), .IN2(n8), .Q(SUM[10]) );
  XOR2X1 U46 ( .IN1(B[9]), .IN2(n7), .Q(SUM[9]) );
  XOR2X1 U47 ( .IN1(B[8]), .IN2(carry[8]), .Q(SUM[8]) );
  AND2X1 U48 ( .IN1(B[0]), .IN2(A[0]), .Q(n23) );
  XOR2X1 U49 ( .IN1(B[0]), .IN2(A[0]), .Q(SUM[0]) );
endmodule


module b15_DW01_add_2 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24;
  wire   [8:2] carry;

  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FADDX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  FADDX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n7), .CO(carry[2]), .S(SUM[1]) );
  AND2X1 U1 ( .IN1(B[10]), .IN2(n9), .Q(n1) );
  AND2X1 U2 ( .IN1(B[11]), .IN2(n1), .Q(n2) );
  AND2X1 U3 ( .IN1(B[14]), .IN2(n11), .Q(n3) );
  AND2X1 U4 ( .IN1(B[15]), .IN2(n3), .Q(n4) );
  AND2X1 U5 ( .IN1(B[18]), .IN2(n13), .Q(n5) );
  AND2X1 U6 ( .IN1(B[19]), .IN2(n5), .Q(n6) );
  AND2X1 U7 ( .IN1(B[0]), .IN2(A[0]), .Q(n7) );
  XNOR2X1 U8 ( .IN1(B[31]), .IN2(n24), .Q(SUM[31]) );
  NAND2X0 U9 ( .IN1(B[30]), .IN2(n23), .QN(n24) );
  XOR2X1 U10 ( .IN1(B[29]), .IN2(n22), .Q(SUM[29]) );
  XOR2X1 U11 ( .IN1(B[28]), .IN2(n21), .Q(SUM[28]) );
  XOR2X1 U12 ( .IN1(B[27]), .IN2(n20), .Q(SUM[27]) );
  XOR2X1 U13 ( .IN1(B[26]), .IN2(n19), .Q(SUM[26]) );
  XOR2X1 U14 ( .IN1(B[25]), .IN2(n18), .Q(SUM[25]) );
  XOR2X1 U15 ( .IN1(B[24]), .IN2(n17), .Q(SUM[24]) );
  XOR2X1 U16 ( .IN1(B[23]), .IN2(n16), .Q(SUM[23]) );
  XOR2X1 U17 ( .IN1(B[22]), .IN2(n15), .Q(SUM[22]) );
  XOR2X1 U18 ( .IN1(B[21]), .IN2(n14), .Q(SUM[21]) );
  XOR2X1 U19 ( .IN1(B[20]), .IN2(n6), .Q(SUM[20]) );
  XOR2X1 U20 ( .IN1(B[19]), .IN2(n5), .Q(SUM[19]) );
  XOR2X1 U21 ( .IN1(B[18]), .IN2(n13), .Q(SUM[18]) );
  XOR2X1 U22 ( .IN1(B[30]), .IN2(n23), .Q(SUM[30]) );
  AND2X1 U23 ( .IN1(B[8]), .IN2(carry[8]), .Q(n8) );
  AND2X1 U24 ( .IN1(B[9]), .IN2(n8), .Q(n9) );
  AND2X1 U25 ( .IN1(B[12]), .IN2(n2), .Q(n10) );
  AND2X1 U26 ( .IN1(B[13]), .IN2(n10), .Q(n11) );
  AND2X1 U27 ( .IN1(B[16]), .IN2(n4), .Q(n12) );
  AND2X1 U28 ( .IN1(B[17]), .IN2(n12), .Q(n13) );
  AND2X1 U29 ( .IN1(B[20]), .IN2(n6), .Q(n14) );
  AND2X1 U30 ( .IN1(B[21]), .IN2(n14), .Q(n15) );
  AND2X1 U31 ( .IN1(B[22]), .IN2(n15), .Q(n16) );
  AND2X1 U32 ( .IN1(B[23]), .IN2(n16), .Q(n17) );
  AND2X1 U33 ( .IN1(B[24]), .IN2(n17), .Q(n18) );
  AND2X1 U34 ( .IN1(B[25]), .IN2(n18), .Q(n19) );
  AND2X1 U35 ( .IN1(B[26]), .IN2(n19), .Q(n20) );
  AND2X1 U36 ( .IN1(B[27]), .IN2(n20), .Q(n21) );
  AND2X1 U37 ( .IN1(B[28]), .IN2(n21), .Q(n22) );
  AND2X1 U38 ( .IN1(B[29]), .IN2(n22), .Q(n23) );
  XOR2X1 U39 ( .IN1(B[17]), .IN2(n12), .Q(SUM[17]) );
  XOR2X1 U40 ( .IN1(B[16]), .IN2(n4), .Q(SUM[16]) );
  XOR2X1 U41 ( .IN1(B[15]), .IN2(n3), .Q(SUM[15]) );
  XOR2X1 U42 ( .IN1(B[14]), .IN2(n11), .Q(SUM[14]) );
  XOR2X1 U43 ( .IN1(B[13]), .IN2(n10), .Q(SUM[13]) );
  XOR2X1 U44 ( .IN1(B[12]), .IN2(n2), .Q(SUM[12]) );
  XOR2X1 U45 ( .IN1(B[11]), .IN2(n1), .Q(SUM[11]) );
  XOR2X1 U46 ( .IN1(B[10]), .IN2(n9), .Q(SUM[10]) );
  XOR2X1 U47 ( .IN1(B[8]), .IN2(carry[8]), .Q(SUM[8]) );
  XOR2X1 U48 ( .IN1(B[9]), .IN2(n8), .Q(SUM[9]) );
  XOR2X1 U49 ( .IN1(B[0]), .IN2(A[0]), .Q(SUM[0]) );
endmodule


module b15_DW01_sub_2 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61;
  assign DIFF[0] = B[0];

  XOR2X1 U1 ( .IN1(n60), .IN2(n25), .Q(DIFF[29]) );
  XOR2X1 U2 ( .IN1(n59), .IN2(n24), .Q(DIFF[28]) );
  XOR2X1 U3 ( .IN1(n58), .IN2(n23), .Q(DIFF[27]) );
  XOR2X1 U4 ( .IN1(n57), .IN2(n22), .Q(DIFF[26]) );
  XOR2X1 U5 ( .IN1(n56), .IN2(n21), .Q(DIFF[25]) );
  XOR2X1 U6 ( .IN1(n55), .IN2(n20), .Q(DIFF[24]) );
  XOR2X1 U7 ( .IN1(n54), .IN2(n19), .Q(DIFF[23]) );
  XOR2X1 U8 ( .IN1(n53), .IN2(n18), .Q(DIFF[22]) );
  XOR2X1 U9 ( .IN1(n52), .IN2(n17), .Q(DIFF[21]) );
  XOR2X1 U10 ( .IN1(n51), .IN2(n16), .Q(DIFF[20]) );
  XOR2X1 U11 ( .IN1(n61), .IN2(n26), .Q(DIFF[30]) );
  AND2X1 U12 ( .IN1(n32), .IN2(n31), .Q(n1) );
  NAND2X0 U13 ( .IN1(n61), .IN2(n26), .QN(n30) );
  XOR2X1 U14 ( .IN1(n50), .IN2(n15), .Q(DIFF[19]) );
  XOR2X1 U15 ( .IN1(n49), .IN2(n14), .Q(DIFF[18]) );
  XOR2X1 U16 ( .IN1(n48), .IN2(n13), .Q(DIFF[17]) );
  AND2X1 U17 ( .IN1(n36), .IN2(n29), .Q(n2) );
  AND2X1 U18 ( .IN1(n37), .IN2(n2), .Q(n3) );
  AND2X1 U19 ( .IN1(n38), .IN2(n3), .Q(n4) );
  AND2X1 U20 ( .IN1(n39), .IN2(n4), .Q(n5) );
  AND2X1 U21 ( .IN1(n40), .IN2(n5), .Q(n6) );
  AND2X1 U22 ( .IN1(n41), .IN2(n6), .Q(n7) );
  AND2X1 U23 ( .IN1(n42), .IN2(n7), .Q(n8) );
  AND2X1 U24 ( .IN1(n43), .IN2(n8), .Q(n9) );
  AND2X1 U25 ( .IN1(n44), .IN2(n9), .Q(n10) );
  AND2X1 U26 ( .IN1(n45), .IN2(n10), .Q(n11) );
  AND2X1 U27 ( .IN1(n46), .IN2(n11), .Q(n12) );
  AND2X1 U28 ( .IN1(n47), .IN2(n12), .Q(n13) );
  AND2X1 U29 ( .IN1(n48), .IN2(n13), .Q(n14) );
  AND2X1 U30 ( .IN1(n49), .IN2(n14), .Q(n15) );
  AND2X1 U31 ( .IN1(n50), .IN2(n15), .Q(n16) );
  AND2X1 U32 ( .IN1(n51), .IN2(n16), .Q(n17) );
  AND2X1 U33 ( .IN1(n52), .IN2(n17), .Q(n18) );
  AND2X1 U34 ( .IN1(n53), .IN2(n18), .Q(n19) );
  AND2X1 U35 ( .IN1(n54), .IN2(n19), .Q(n20) );
  AND2X1 U36 ( .IN1(n55), .IN2(n20), .Q(n21) );
  AND2X1 U37 ( .IN1(n56), .IN2(n21), .Q(n22) );
  AND2X1 U38 ( .IN1(n57), .IN2(n22), .Q(n23) );
  AND2X1 U39 ( .IN1(n58), .IN2(n23), .Q(n24) );
  AND2X1 U40 ( .IN1(n59), .IN2(n24), .Q(n25) );
  AND2X1 U41 ( .IN1(n60), .IN2(n25), .Q(n26) );
  AND2X1 U42 ( .IN1(n34), .IN2(n28), .Q(n27) );
  AND2X1 U43 ( .IN1(n33), .IN2(n1), .Q(n28) );
  AND2X1 U44 ( .IN1(n35), .IN2(n27), .Q(n29) );
  XOR2X1 U45 ( .IN1(n47), .IN2(n12), .Q(DIFF[16]) );
  XOR2X1 U46 ( .IN1(n46), .IN2(n11), .Q(DIFF[15]) );
  XOR2X1 U47 ( .IN1(n45), .IN2(n10), .Q(DIFF[14]) );
  XOR2X1 U48 ( .IN1(n44), .IN2(n9), .Q(DIFF[13]) );
  XOR2X1 U49 ( .IN1(n43), .IN2(n8), .Q(DIFF[12]) );
  XOR2X1 U50 ( .IN1(n42), .IN2(n7), .Q(DIFF[11]) );
  XOR2X1 U51 ( .IN1(n41), .IN2(n6), .Q(DIFF[10]) );
  XOR2X1 U52 ( .IN1(n40), .IN2(n5), .Q(DIFF[9]) );
  XOR2X1 U53 ( .IN1(n39), .IN2(n4), .Q(DIFF[8]) );
  XOR2X1 U54 ( .IN1(n38), .IN2(n3), .Q(DIFF[7]) );
  XOR2X1 U55 ( .IN1(n37), .IN2(n2), .Q(DIFF[6]) );
  XOR2X1 U56 ( .IN1(n36), .IN2(n29), .Q(DIFF[5]) );
  XOR2X1 U57 ( .IN1(n34), .IN2(n28), .Q(DIFF[3]) );
  XOR2X1 U58 ( .IN1(n33), .IN2(n1), .Q(DIFF[2]) );
  XOR2X1 U59 ( .IN1(n32), .IN2(n31), .Q(DIFF[1]) );
  XOR2X1 U60 ( .IN1(B[31]), .IN2(n30), .Q(DIFF[31]) );
  XOR2X1 U61 ( .IN1(n35), .IN2(n27), .Q(DIFF[4]) );
  INVX0 U62 ( .IN(B[0]), .QN(n31) );
  INVX0 U63 ( .IN(B[6]), .QN(n37) );
  INVX0 U64 ( .IN(B[7]), .QN(n38) );
  INVX0 U65 ( .IN(B[8]), .QN(n39) );
  INVX0 U66 ( .IN(B[9]), .QN(n40) );
  INVX0 U67 ( .IN(B[10]), .QN(n41) );
  INVX0 U68 ( .IN(B[11]), .QN(n42) );
  INVX0 U69 ( .IN(B[12]), .QN(n43) );
  INVX0 U70 ( .IN(B[13]), .QN(n44) );
  INVX0 U71 ( .IN(B[14]), .QN(n45) );
  INVX0 U72 ( .IN(B[15]), .QN(n46) );
  INVX0 U73 ( .IN(B[4]), .QN(n35) );
  INVX0 U74 ( .IN(B[3]), .QN(n34) );
  INVX0 U75 ( .IN(B[2]), .QN(n33) );
  INVX0 U76 ( .IN(B[1]), .QN(n32) );
  INVX0 U77 ( .IN(B[5]), .QN(n36) );
  INVX0 U78 ( .IN(B[16]), .QN(n47) );
  INVX0 U79 ( .IN(B[17]), .QN(n48) );
  INVX0 U80 ( .IN(B[18]), .QN(n49) );
  INVX0 U81 ( .IN(B[19]), .QN(n50) );
  INVX0 U82 ( .IN(B[20]), .QN(n51) );
  INVX0 U83 ( .IN(B[21]), .QN(n52) );
  INVX0 U84 ( .IN(B[22]), .QN(n53) );
  INVX0 U85 ( .IN(B[23]), .QN(n54) );
  INVX0 U86 ( .IN(B[24]), .QN(n55) );
  INVX0 U87 ( .IN(B[25]), .QN(n56) );
  INVX0 U88 ( .IN(B[26]), .QN(n57) );
  INVX0 U89 ( .IN(B[27]), .QN(n58) );
  INVX0 U90 ( .IN(B[28]), .QN(n59) );
  INVX0 U91 ( .IN(B[29]), .QN(n60) );
  INVX0 U92 ( .IN(B[30]), .QN(n61) );
endmodule


module b15_DW01_inc_0 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;

  wire   [31:2] carry;

  HADDX1 U1_1_30 ( .A0(A[30]), .B0(carry[30]), .C1(carry[31]), .SO(SUM[30]) );
  HADDX1 U1_1_29 ( .A0(A[29]), .B0(carry[29]), .C1(carry[30]), .SO(SUM[29]) );
  HADDX1 U1_1_28 ( .A0(A[28]), .B0(carry[28]), .C1(carry[29]), .SO(SUM[28]) );
  HADDX1 U1_1_27 ( .A0(A[27]), .B0(carry[27]), .C1(carry[28]), .SO(SUM[27]) );
  HADDX1 U1_1_26 ( .A0(A[26]), .B0(carry[26]), .C1(carry[27]), .SO(SUM[26]) );
  HADDX1 U1_1_25 ( .A0(A[25]), .B0(carry[25]), .C1(carry[26]), .SO(SUM[25]) );
  HADDX1 U1_1_24 ( .A0(A[24]), .B0(carry[24]), .C1(carry[25]), .SO(SUM[24]) );
  HADDX1 U1_1_23 ( .A0(A[23]), .B0(carry[23]), .C1(carry[24]), .SO(SUM[23]) );
  HADDX1 U1_1_22 ( .A0(A[22]), .B0(carry[22]), .C1(carry[23]), .SO(SUM[22]) );
  HADDX1 U1_1_21 ( .A0(A[21]), .B0(carry[21]), .C1(carry[22]), .SO(SUM[21]) );
  HADDX1 U1_1_20 ( .A0(A[20]), .B0(carry[20]), .C1(carry[21]), .SO(SUM[20]) );
  HADDX1 U1_1_19 ( .A0(A[19]), .B0(carry[19]), .C1(carry[20]), .SO(SUM[19]) );
  HADDX1 U1_1_18 ( .A0(A[18]), .B0(carry[18]), .C1(carry[19]), .SO(SUM[18]) );
  HADDX1 U1_1_17 ( .A0(A[17]), .B0(carry[17]), .C1(carry[18]), .SO(SUM[17]) );
  HADDX1 U1_1_16 ( .A0(A[16]), .B0(carry[16]), .C1(carry[17]), .SO(SUM[16]) );
  HADDX1 U1_1_15 ( .A0(A[15]), .B0(carry[15]), .C1(carry[16]), .SO(SUM[15]) );
  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .IN(A[0]), .QN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[31]), .IN2(A[31]), .Q(SUM[31]) );
endmodule


module b15_DW01_inc_1 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;

  wire   [31:2] carry;

  HADDX1 U1_1_30 ( .A0(A[30]), .B0(carry[30]), .C1(carry[31]), .SO(SUM[30]) );
  HADDX1 U1_1_29 ( .A0(A[29]), .B0(carry[29]), .C1(carry[30]), .SO(SUM[29]) );
  HADDX1 U1_1_28 ( .A0(A[28]), .B0(carry[28]), .C1(carry[29]), .SO(SUM[28]) );
  HADDX1 U1_1_27 ( .A0(A[27]), .B0(carry[27]), .C1(carry[28]), .SO(SUM[27]) );
  HADDX1 U1_1_26 ( .A0(A[26]), .B0(carry[26]), .C1(carry[27]), .SO(SUM[26]) );
  HADDX1 U1_1_25 ( .A0(A[25]), .B0(carry[25]), .C1(carry[26]), .SO(SUM[25]) );
  HADDX1 U1_1_24 ( .A0(A[24]), .B0(carry[24]), .C1(carry[25]), .SO(SUM[24]) );
  HADDX1 U1_1_23 ( .A0(A[23]), .B0(carry[23]), .C1(carry[24]), .SO(SUM[23]) );
  HADDX1 U1_1_22 ( .A0(A[22]), .B0(carry[22]), .C1(carry[23]), .SO(SUM[22]) );
  HADDX1 U1_1_21 ( .A0(A[21]), .B0(carry[21]), .C1(carry[22]), .SO(SUM[21]) );
  HADDX1 U1_1_20 ( .A0(A[20]), .B0(carry[20]), .C1(carry[21]), .SO(SUM[20]) );
  HADDX1 U1_1_19 ( .A0(A[19]), .B0(carry[19]), .C1(carry[20]), .SO(SUM[19]) );
  HADDX1 U1_1_18 ( .A0(A[18]), .B0(carry[18]), .C1(carry[19]), .SO(SUM[18]) );
  HADDX1 U1_1_17 ( .A0(A[17]), .B0(carry[17]), .C1(carry[18]), .SO(SUM[17]) );
  HADDX1 U1_1_16 ( .A0(A[16]), .B0(carry[16]), .C1(carry[17]), .SO(SUM[16]) );
  HADDX1 U1_1_15 ( .A0(A[15]), .B0(carry[15]), .C1(carry[16]), .SO(SUM[15]) );
  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .IN(A[0]), .QN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[31]), .IN2(A[31]), .Q(SUM[31]) );
endmodule


module b15_DW01_sub_3 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61;
  assign DIFF[0] = B[0];

  AND2X1 U1 ( .IN1(n59), .IN2(n29), .Q(n1) );
  AND2X1 U2 ( .IN1(n58), .IN2(n1), .Q(n2) );
  AND2X1 U3 ( .IN1(n55), .IN2(n16), .Q(n3) );
  AND2X1 U4 ( .IN1(n54), .IN2(n3), .Q(n4) );
  AND2X1 U5 ( .IN1(n52), .IN2(n17), .Q(n5) );
  AND2X1 U6 ( .IN1(n51), .IN2(n5), .Q(n6) );
  AND2X1 U7 ( .IN1(n50), .IN2(n6), .Q(n7) );
  AND2X1 U8 ( .IN1(n49), .IN2(n7), .Q(n8) );
  AND2X1 U9 ( .IN1(n48), .IN2(n8), .Q(n9) );
  AND2X1 U10 ( .IN1(n47), .IN2(n9), .Q(n10) );
  AND2X1 U11 ( .IN1(n46), .IN2(n10), .Q(n11) );
  AND2X1 U12 ( .IN1(n44), .IN2(n18), .Q(n12) );
  AND2X1 U13 ( .IN1(n43), .IN2(n12), .Q(n13) );
  AND2X1 U14 ( .IN1(n42), .IN2(n13), .Q(n14) );
  XOR2X1 U15 ( .IN1(n31), .IN2(n28), .Q(DIFF[30]) );
  AND2X1 U16 ( .IN1(n57), .IN2(n2), .Q(n15) );
  AND2X1 U17 ( .IN1(n56), .IN2(n15), .Q(n16) );
  AND2X1 U18 ( .IN1(n53), .IN2(n4), .Q(n17) );
  AND2X1 U19 ( .IN1(n45), .IN2(n11), .Q(n18) );
  AND2X1 U20 ( .IN1(n41), .IN2(n14), .Q(n19) );
  AND2X1 U21 ( .IN1(n40), .IN2(n19), .Q(n20) );
  AND2X1 U22 ( .IN1(n39), .IN2(n20), .Q(n21) );
  AND2X1 U23 ( .IN1(n38), .IN2(n21), .Q(n22) );
  AND2X1 U24 ( .IN1(n37), .IN2(n22), .Q(n23) );
  AND2X1 U25 ( .IN1(n36), .IN2(n23), .Q(n24) );
  AND2X1 U26 ( .IN1(n35), .IN2(n24), .Q(n25) );
  AND2X1 U27 ( .IN1(n34), .IN2(n25), .Q(n26) );
  AND2X1 U28 ( .IN1(n33), .IN2(n26), .Q(n27) );
  AND2X1 U29 ( .IN1(n32), .IN2(n27), .Q(n28) );
  XOR2X1 U30 ( .IN1(n32), .IN2(n27), .Q(DIFF[29]) );
  XOR2X1 U31 ( .IN1(n33), .IN2(n26), .Q(DIFF[28]) );
  XOR2X1 U32 ( .IN1(n34), .IN2(n25), .Q(DIFF[27]) );
  XOR2X1 U33 ( .IN1(n35), .IN2(n24), .Q(DIFF[26]) );
  XOR2X1 U34 ( .IN1(n36), .IN2(n23), .Q(DIFF[25]) );
  XOR2X1 U35 ( .IN1(n37), .IN2(n22), .Q(DIFF[24]) );
  XOR2X1 U36 ( .IN1(n38), .IN2(n21), .Q(DIFF[23]) );
  XOR2X1 U37 ( .IN1(n39), .IN2(n20), .Q(DIFF[22]) );
  XOR2X1 U38 ( .IN1(n40), .IN2(n19), .Q(DIFF[21]) );
  XOR2X1 U39 ( .IN1(n41), .IN2(n14), .Q(DIFF[20]) );
  XOR2X1 U40 ( .IN1(n57), .IN2(n2), .Q(DIFF[4]) );
  XOR2X1 U41 ( .IN1(n58), .IN2(n1), .Q(DIFF[3]) );
  XOR2X1 U42 ( .IN1(n59), .IN2(n29), .Q(DIFF[2]) );
  XOR2X1 U43 ( .IN1(n56), .IN2(n15), .Q(DIFF[5]) );
  XOR2X1 U44 ( .IN1(n42), .IN2(n13), .Q(DIFF[19]) );
  XOR2X1 U45 ( .IN1(n43), .IN2(n12), .Q(DIFF[18]) );
  XOR2X1 U46 ( .IN1(n44), .IN2(n18), .Q(DIFF[17]) );
  XOR2X1 U47 ( .IN1(n45), .IN2(n11), .Q(DIFF[16]) );
  XOR2X1 U48 ( .IN1(n46), .IN2(n10), .Q(DIFF[15]) );
  XOR2X1 U49 ( .IN1(n47), .IN2(n9), .Q(DIFF[14]) );
  XOR2X1 U50 ( .IN1(n48), .IN2(n8), .Q(DIFF[13]) );
  XOR2X1 U51 ( .IN1(n49), .IN2(n7), .Q(DIFF[12]) );
  XOR2X1 U52 ( .IN1(n50), .IN2(n6), .Q(DIFF[11]) );
  XOR2X1 U53 ( .IN1(n51), .IN2(n5), .Q(DIFF[10]) );
  XOR2X1 U54 ( .IN1(n52), .IN2(n17), .Q(DIFF[9]) );
  XOR2X1 U55 ( .IN1(n53), .IN2(n4), .Q(DIFF[8]) );
  XOR2X1 U56 ( .IN1(n54), .IN2(n3), .Q(DIFF[7]) );
  XOR2X1 U57 ( .IN1(n55), .IN2(n16), .Q(DIFF[6]) );
  XOR2X1 U58 ( .IN1(B[31]), .IN2(n30), .Q(DIFF[31]) );
  NAND2X0 U59 ( .IN1(n31), .IN2(n28), .QN(n30) );
  INVX0 U60 ( .IN(B[2]), .QN(n59) );
  INVX0 U61 ( .IN(B[3]), .QN(n58) );
  INVX0 U62 ( .IN(B[4]), .QN(n57) );
  INVX0 U63 ( .IN(B[5]), .QN(n56) );
  INVX0 U64 ( .IN(B[6]), .QN(n55) );
  INVX0 U65 ( .IN(B[7]), .QN(n54) );
  INVX0 U66 ( .IN(B[8]), .QN(n53) );
  INVX0 U67 ( .IN(B[9]), .QN(n52) );
  INVX0 U68 ( .IN(B[10]), .QN(n51) );
  INVX0 U69 ( .IN(B[11]), .QN(n50) );
  INVX0 U70 ( .IN(B[12]), .QN(n49) );
  INVX0 U71 ( .IN(B[13]), .QN(n48) );
  INVX0 U72 ( .IN(B[14]), .QN(n47) );
  INVX0 U73 ( .IN(B[20]), .QN(n41) );
  INVX0 U74 ( .IN(B[21]), .QN(n40) );
  INVX0 U75 ( .IN(B[22]), .QN(n39) );
  INVX0 U76 ( .IN(B[23]), .QN(n38) );
  INVX0 U77 ( .IN(B[24]), .QN(n37) );
  INVX0 U78 ( .IN(B[25]), .QN(n36) );
  INVX0 U79 ( .IN(B[26]), .QN(n35) );
  INVX0 U80 ( .IN(B[27]), .QN(n34) );
  INVX0 U81 ( .IN(B[28]), .QN(n33) );
  INVX0 U82 ( .IN(B[29]), .QN(n32) );
  INVX0 U83 ( .IN(B[30]), .QN(n31) );
  INVX0 U84 ( .IN(B[15]), .QN(n46) );
  INVX0 U85 ( .IN(B[16]), .QN(n45) );
  INVX0 U86 ( .IN(B[17]), .QN(n44) );
  INVX0 U87 ( .IN(B[18]), .QN(n43) );
  INVX0 U88 ( .IN(B[19]), .QN(n42) );
  AND2X1 U89 ( .IN1(n60), .IN2(n61), .Q(n29) );
  INVX0 U90 ( .IN(B[1]), .QN(n60) );
  XOR2X1 U91 ( .IN1(n60), .IN2(n61), .Q(DIFF[1]) );
  INVX0 U92 ( .IN(B[0]), .QN(n61) );
endmodule


module b15_DW01_add_6 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28;
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  AND2X1 U1 ( .IN1(n23), .IN2(A[5]), .Q(n1) );
  AND2X1 U2 ( .IN1(n1), .IN2(A[6]), .Q(n2) );
  AND2X1 U3 ( .IN1(n2), .IN2(A[7]), .Q(n3) );
  AND2X1 U4 ( .IN1(n3), .IN2(A[8]), .Q(n4) );
  AND2X1 U5 ( .IN1(n4), .IN2(A[9]), .Q(n5) );
  AND2X1 U6 ( .IN1(n5), .IN2(A[10]), .Q(n6) );
  AND2X1 U7 ( .IN1(n24), .IN2(A[12]), .Q(n7) );
  AND2X1 U8 ( .IN1(n7), .IN2(A[13]), .Q(n8) );
  AND2X1 U9 ( .IN1(n8), .IN2(A[14]), .Q(n9) );
  AND2X1 U10 ( .IN1(n25), .IN2(A[16]), .Q(n10) );
  AND2X1 U11 ( .IN1(n10), .IN2(A[17]), .Q(n11) );
  AND2X1 U12 ( .IN1(n11), .IN2(A[18]), .Q(n12) );
  AND2X1 U13 ( .IN1(n26), .IN2(A[20]), .Q(n13) );
  AND2X1 U14 ( .IN1(n13), .IN2(A[21]), .Q(n14) );
  AND2X1 U15 ( .IN1(n14), .IN2(A[22]), .Q(n15) );
  AND2X1 U16 ( .IN1(n27), .IN2(A[24]), .Q(n16) );
  AND2X1 U17 ( .IN1(n16), .IN2(A[25]), .Q(n17) );
  AND2X1 U18 ( .IN1(n17), .IN2(A[26]), .Q(n18) );
  AND2X1 U19 ( .IN1(n18), .IN2(A[27]), .Q(n19) );
  AND2X1 U20 ( .IN1(n19), .IN2(A[28]), .Q(n20) );
  AND2X1 U21 ( .IN1(n20), .IN2(A[29]), .Q(n21) );
  XOR2X1 U22 ( .IN1(n19), .IN2(A[28]), .Q(SUM[28]) );
  XOR2X1 U23 ( .IN1(n18), .IN2(A[27]), .Q(SUM[27]) );
  XOR2X1 U24 ( .IN1(n17), .IN2(A[26]), .Q(SUM[26]) );
  XOR2X1 U25 ( .IN1(n16), .IN2(A[25]), .Q(SUM[25]) );
  XOR2X1 U26 ( .IN1(n27), .IN2(A[24]), .Q(SUM[24]) );
  XOR2X1 U27 ( .IN1(n15), .IN2(A[23]), .Q(SUM[23]) );
  XOR2X1 U28 ( .IN1(n14), .IN2(A[22]), .Q(SUM[22]) );
  XOR2X1 U29 ( .IN1(n20), .IN2(A[29]), .Q(SUM[29]) );
  XOR2X1 U30 ( .IN1(n21), .IN2(A[30]), .Q(SUM[30]) );
  AND2X1 U31 ( .IN1(A[2]), .IN2(A[3]), .Q(n22) );
  AND2X1 U32 ( .IN1(n22), .IN2(A[4]), .Q(n23) );
  AND2X1 U33 ( .IN1(n6), .IN2(A[11]), .Q(n24) );
  AND2X1 U34 ( .IN1(n9), .IN2(A[15]), .Q(n25) );
  AND2X1 U35 ( .IN1(n12), .IN2(A[19]), .Q(n26) );
  AND2X1 U36 ( .IN1(n15), .IN2(A[23]), .Q(n27) );
  XNOR2X1 U37 ( .IN1(n28), .IN2(A[31]), .Q(SUM[31]) );
  NAND2X0 U38 ( .IN1(n21), .IN2(A[30]), .QN(n28) );
  XOR2X1 U39 ( .IN1(n13), .IN2(A[21]), .Q(SUM[21]) );
  XOR2X1 U40 ( .IN1(n26), .IN2(A[20]), .Q(SUM[20]) );
  XOR2X1 U41 ( .IN1(n12), .IN2(A[19]), .Q(SUM[19]) );
  XOR2X1 U42 ( .IN1(n11), .IN2(A[18]), .Q(SUM[18]) );
  XOR2X1 U43 ( .IN1(n10), .IN2(A[17]), .Q(SUM[17]) );
  XOR2X1 U44 ( .IN1(n25), .IN2(A[16]), .Q(SUM[16]) );
  XOR2X1 U45 ( .IN1(n9), .IN2(A[15]), .Q(SUM[15]) );
  XOR2X1 U46 ( .IN1(n8), .IN2(A[14]), .Q(SUM[14]) );
  XOR2X1 U47 ( .IN1(n7), .IN2(A[13]), .Q(SUM[13]) );
  XOR2X1 U48 ( .IN1(n24), .IN2(A[12]), .Q(SUM[12]) );
  XOR2X1 U49 ( .IN1(n6), .IN2(A[11]), .Q(SUM[11]) );
  XOR2X1 U50 ( .IN1(n5), .IN2(A[10]), .Q(SUM[10]) );
  XOR2X1 U51 ( .IN1(n4), .IN2(A[9]), .Q(SUM[9]) );
  XOR2X1 U52 ( .IN1(n3), .IN2(A[8]), .Q(SUM[8]) );
  XOR2X1 U53 ( .IN1(n2), .IN2(A[7]), .Q(SUM[7]) );
  XOR2X1 U54 ( .IN1(n1), .IN2(A[6]), .Q(SUM[6]) );
  XOR2X1 U55 ( .IN1(n23), .IN2(A[5]), .Q(SUM[5]) );
  XOR2X1 U56 ( .IN1(A[2]), .IN2(A[3]), .Q(SUM[3]) );
  XOR2X1 U57 ( .IN1(n22), .IN2(A[4]), .Q(SUM[4]) );
  INVX0 U58 ( .IN(A[2]), .QN(SUM[2]) );
endmodule


module b15_DW01_add_9 ( A, B, CI, SUM, CO );
  input [29:0] A;
  input [29:0] B;
  output [29:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29;

  AND2X1 U1 ( .IN1(B[19]), .IN2(n29), .Q(n1) );
  AND2X1 U2 ( .IN1(B[20]), .IN2(n1), .Q(n2) );
  AND2X1 U3 ( .IN1(B[21]), .IN2(n2), .Q(n3) );
  AND2X1 U4 ( .IN1(B[22]), .IN2(n3), .Q(n4) );
  AND2X1 U5 ( .IN1(B[23]), .IN2(n4), .Q(n5) );
  AND2X1 U6 ( .IN1(B[24]), .IN2(n5), .Q(n6) );
  AND2X1 U7 ( .IN1(B[25]), .IN2(n6), .Q(n7) );
  AND2X1 U8 ( .IN1(B[26]), .IN2(n7), .Q(n8) );
  AND2X1 U9 ( .IN1(B[27]), .IN2(n8), .Q(n9) );
  AND2X1 U10 ( .IN1(B[28]), .IN2(n9), .Q(n10) );
  AND2X1 U11 ( .IN1(B[2]), .IN2(n13), .Q(n11) );
  XOR2X1 U12 ( .IN1(B[29]), .IN2(n10), .Q(SUM[29]) );
  XOR2X1 U13 ( .IN1(B[28]), .IN2(n9), .Q(SUM[28]) );
  AND2X1 U14 ( .IN1(B[0]), .IN2(A[0]), .Q(n12) );
  AND2X1 U15 ( .IN1(B[1]), .IN2(n12), .Q(n13) );
  AND2X1 U16 ( .IN1(B[3]), .IN2(n11), .Q(n14) );
  AND2X1 U17 ( .IN1(B[4]), .IN2(n14), .Q(n15) );
  AND2X1 U18 ( .IN1(B[5]), .IN2(n15), .Q(n16) );
  AND2X1 U19 ( .IN1(B[6]), .IN2(n16), .Q(n17) );
  AND2X1 U20 ( .IN1(B[7]), .IN2(n17), .Q(n18) );
  AND2X1 U21 ( .IN1(B[8]), .IN2(n18), .Q(n19) );
  AND2X1 U22 ( .IN1(B[9]), .IN2(n19), .Q(n20) );
  AND2X1 U23 ( .IN1(B[10]), .IN2(n20), .Q(n21) );
  AND2X1 U24 ( .IN1(B[11]), .IN2(n21), .Q(n22) );
  AND2X1 U25 ( .IN1(B[12]), .IN2(n22), .Q(n23) );
  AND2X1 U26 ( .IN1(B[13]), .IN2(n23), .Q(n24) );
  AND2X1 U27 ( .IN1(B[14]), .IN2(n24), .Q(n25) );
  AND2X1 U28 ( .IN1(B[15]), .IN2(n25), .Q(n26) );
  AND2X1 U29 ( .IN1(B[16]), .IN2(n26), .Q(n27) );
  AND2X1 U30 ( .IN1(B[17]), .IN2(n27), .Q(n28) );
  AND2X1 U31 ( .IN1(B[18]), .IN2(n28), .Q(n29) );
  XOR2X1 U32 ( .IN1(B[27]), .IN2(n8), .Q(SUM[27]) );
  XOR2X1 U33 ( .IN1(B[26]), .IN2(n7), .Q(SUM[26]) );
  XOR2X1 U34 ( .IN1(B[25]), .IN2(n6), .Q(SUM[25]) );
  XOR2X1 U35 ( .IN1(B[24]), .IN2(n5), .Q(SUM[24]) );
  XOR2X1 U36 ( .IN1(B[23]), .IN2(n4), .Q(SUM[23]) );
  XOR2X1 U37 ( .IN1(B[22]), .IN2(n3), .Q(SUM[22]) );
  XOR2X1 U38 ( .IN1(B[21]), .IN2(n2), .Q(SUM[21]) );
  XOR2X1 U39 ( .IN1(B[20]), .IN2(n1), .Q(SUM[20]) );
  XOR2X1 U40 ( .IN1(B[19]), .IN2(n29), .Q(SUM[19]) );
  XOR2X1 U41 ( .IN1(B[18]), .IN2(n28), .Q(SUM[18]) );
  XOR2X1 U42 ( .IN1(B[17]), .IN2(n27), .Q(SUM[17]) );
  XOR2X1 U43 ( .IN1(B[16]), .IN2(n26), .Q(SUM[16]) );
  XOR2X1 U44 ( .IN1(B[15]), .IN2(n25), .Q(SUM[15]) );
  XOR2X1 U45 ( .IN1(B[14]), .IN2(n24), .Q(SUM[14]) );
  XOR2X1 U46 ( .IN1(B[13]), .IN2(n23), .Q(SUM[13]) );
  XOR2X1 U47 ( .IN1(B[12]), .IN2(n22), .Q(SUM[12]) );
  XOR2X1 U48 ( .IN1(B[11]), .IN2(n21), .Q(SUM[11]) );
  XOR2X1 U49 ( .IN1(B[10]), .IN2(n20), .Q(SUM[10]) );
  XOR2X1 U50 ( .IN1(B[9]), .IN2(n19), .Q(SUM[9]) );
  XOR2X1 U51 ( .IN1(B[8]), .IN2(n18), .Q(SUM[8]) );
  XOR2X1 U52 ( .IN1(B[7]), .IN2(n17), .Q(SUM[7]) );
  XOR2X1 U53 ( .IN1(B[6]), .IN2(n16), .Q(SUM[6]) );
  XOR2X1 U54 ( .IN1(B[5]), .IN2(n15), .Q(SUM[5]) );
  XOR2X1 U55 ( .IN1(B[4]), .IN2(n14), .Q(SUM[4]) );
  XOR2X1 U56 ( .IN1(B[3]), .IN2(n11), .Q(SUM[3]) );
  XOR2X1 U57 ( .IN1(B[2]), .IN2(n13), .Q(SUM[2]) );
  XOR2X1 U58 ( .IN1(B[1]), .IN2(n12), .Q(SUM[1]) );
  XOR2X1 U59 ( .IN1(B[0]), .IN2(A[0]), .Q(SUM[0]) );
endmodule


module b15_DW01_add_10 ( A, B, CI, SUM, CO );
  input [29:0] A;
  input [29:0] B;
  output [29:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29;

  AND2X1 U1 ( .IN1(B[18]), .IN2(n29), .Q(n1) );
  AND2X1 U2 ( .IN1(B[19]), .IN2(n1), .Q(n2) );
  AND2X1 U3 ( .IN1(B[20]), .IN2(n2), .Q(n3) );
  AND2X1 U4 ( .IN1(B[21]), .IN2(n3), .Q(n4) );
  AND2X1 U5 ( .IN1(B[22]), .IN2(n4), .Q(n5) );
  AND2X1 U6 ( .IN1(B[23]), .IN2(n5), .Q(n6) );
  AND2X1 U7 ( .IN1(B[24]), .IN2(n6), .Q(n7) );
  AND2X1 U8 ( .IN1(B[25]), .IN2(n7), .Q(n8) );
  AND2X1 U9 ( .IN1(B[26]), .IN2(n8), .Q(n9) );
  AND2X1 U10 ( .IN1(B[27]), .IN2(n9), .Q(n10) );
  AND2X1 U11 ( .IN1(B[0]), .IN2(A[0]), .Q(n11) );
  AND2X1 U12 ( .IN1(B[28]), .IN2(n10), .Q(n12) );
  XOR2X1 U13 ( .IN1(B[29]), .IN2(n12), .Q(SUM[29]) );
  XOR2X1 U14 ( .IN1(B[28]), .IN2(n10), .Q(SUM[28]) );
  AND2X1 U15 ( .IN1(B[1]), .IN2(n11), .Q(n13) );
  AND2X1 U16 ( .IN1(B[2]), .IN2(n13), .Q(n14) );
  AND2X1 U17 ( .IN1(B[3]), .IN2(n14), .Q(n15) );
  AND2X1 U18 ( .IN1(B[4]), .IN2(n15), .Q(n16) );
  AND2X1 U19 ( .IN1(B[5]), .IN2(n16), .Q(n17) );
  AND2X1 U20 ( .IN1(B[6]), .IN2(n17), .Q(n18) );
  AND2X1 U21 ( .IN1(B[7]), .IN2(n18), .Q(n19) );
  AND2X1 U22 ( .IN1(B[8]), .IN2(n19), .Q(n20) );
  AND2X1 U23 ( .IN1(B[9]), .IN2(n20), .Q(n21) );
  AND2X1 U24 ( .IN1(B[10]), .IN2(n21), .Q(n22) );
  AND2X1 U25 ( .IN1(B[11]), .IN2(n22), .Q(n23) );
  AND2X1 U26 ( .IN1(B[12]), .IN2(n23), .Q(n24) );
  AND2X1 U27 ( .IN1(B[13]), .IN2(n24), .Q(n25) );
  AND2X1 U28 ( .IN1(B[14]), .IN2(n25), .Q(n26) );
  AND2X1 U29 ( .IN1(B[15]), .IN2(n26), .Q(n27) );
  AND2X1 U30 ( .IN1(B[16]), .IN2(n27), .Q(n28) );
  AND2X1 U31 ( .IN1(B[17]), .IN2(n28), .Q(n29) );
  XOR2X1 U32 ( .IN1(B[27]), .IN2(n9), .Q(SUM[27]) );
  XOR2X1 U33 ( .IN1(B[26]), .IN2(n8), .Q(SUM[26]) );
  XOR2X1 U34 ( .IN1(B[25]), .IN2(n7), .Q(SUM[25]) );
  XOR2X1 U35 ( .IN1(B[24]), .IN2(n6), .Q(SUM[24]) );
  XOR2X1 U36 ( .IN1(B[23]), .IN2(n5), .Q(SUM[23]) );
  XOR2X1 U37 ( .IN1(B[22]), .IN2(n4), .Q(SUM[22]) );
  XOR2X1 U38 ( .IN1(B[21]), .IN2(n3), .Q(SUM[21]) );
  XOR2X1 U39 ( .IN1(B[20]), .IN2(n2), .Q(SUM[20]) );
  XOR2X1 U40 ( .IN1(B[19]), .IN2(n1), .Q(SUM[19]) );
  XOR2X1 U41 ( .IN1(B[18]), .IN2(n29), .Q(SUM[18]) );
  XOR2X1 U42 ( .IN1(B[17]), .IN2(n28), .Q(SUM[17]) );
  XOR2X1 U43 ( .IN1(B[16]), .IN2(n27), .Q(SUM[16]) );
  XOR2X1 U44 ( .IN1(B[15]), .IN2(n26), .Q(SUM[15]) );
  XOR2X1 U45 ( .IN1(B[14]), .IN2(n25), .Q(SUM[14]) );
  XOR2X1 U46 ( .IN1(B[13]), .IN2(n24), .Q(SUM[13]) );
  XOR2X1 U47 ( .IN1(B[12]), .IN2(n23), .Q(SUM[12]) );
  XOR2X1 U48 ( .IN1(B[11]), .IN2(n22), .Q(SUM[11]) );
  XOR2X1 U49 ( .IN1(B[10]), .IN2(n21), .Q(SUM[10]) );
  XOR2X1 U50 ( .IN1(B[9]), .IN2(n20), .Q(SUM[9]) );
  XOR2X1 U51 ( .IN1(B[8]), .IN2(n19), .Q(SUM[8]) );
  XOR2X1 U52 ( .IN1(B[7]), .IN2(n18), .Q(SUM[7]) );
  XOR2X1 U53 ( .IN1(B[6]), .IN2(n17), .Q(SUM[6]) );
  XOR2X1 U54 ( .IN1(B[5]), .IN2(n16), .Q(SUM[5]) );
  XOR2X1 U55 ( .IN1(B[4]), .IN2(n15), .Q(SUM[4]) );
  XOR2X1 U56 ( .IN1(B[3]), .IN2(n14), .Q(SUM[3]) );
  XOR2X1 U57 ( .IN1(B[2]), .IN2(n13), .Q(SUM[2]) );
  XOR2X1 U58 ( .IN1(B[1]), .IN2(n11), .Q(SUM[1]) );
  XOR2X1 U59 ( .IN1(B[0]), .IN2(A[0]), .Q(SUM[0]) );
endmodule


module b15_DW01_add_11 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   carry_3_, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30;

  XOR2X1 U1 ( .IN1(n29), .IN2(n10), .Q(SUM[2]) );
  LSDNENX1 U2 ( .D(n10), .ENB(n29), .Q(carry_3_) );
  AND2X1 U3 ( .IN1(n28), .IN2(A[21]), .Q(n1) );
  AND2X1 U4 ( .IN1(n1), .IN2(A[22]), .Q(n2) );
  AND2X1 U5 ( .IN1(n2), .IN2(A[23]), .Q(n3) );
  AND2X1 U6 ( .IN1(n3), .IN2(A[24]), .Q(n4) );
  AND2X1 U7 ( .IN1(n4), .IN2(A[25]), .Q(n5) );
  AND2X1 U8 ( .IN1(n5), .IN2(A[26]), .Q(n6) );
  AND2X1 U9 ( .IN1(n6), .IN2(A[27]), .Q(n7) );
  AND2X1 U10 ( .IN1(n7), .IN2(A[28]), .Q(n8) );
  AND2X1 U11 ( .IN1(n8), .IN2(A[29]), .Q(n9) );
  XOR2X1 U12 ( .IN1(n8), .IN2(A[29]), .Q(SUM[29]) );
  XOR2X1 U13 ( .IN1(n7), .IN2(A[28]), .Q(SUM[28]) );
  XOR2X1 U14 ( .IN1(n6), .IN2(A[27]), .Q(SUM[27]) );
  XOR2X1 U15 ( .IN1(n5), .IN2(A[26]), .Q(SUM[26]) );
  XOR2X1 U16 ( .IN1(n4), .IN2(A[25]), .Q(SUM[25]) );
  XOR2X1 U17 ( .IN1(n3), .IN2(A[24]), .Q(SUM[24]) );
  XOR2X1 U18 ( .IN1(n2), .IN2(A[23]), .Q(SUM[23]) );
  XOR2X1 U19 ( .IN1(n1), .IN2(A[22]), .Q(SUM[22]) );
  XOR2X1 U20 ( .IN1(n28), .IN2(A[21]), .Q(SUM[21]) );
  XOR2X1 U21 ( .IN1(n27), .IN2(A[20]), .Q(SUM[20]) );
  XOR2X1 U22 ( .IN1(n26), .IN2(A[19]), .Q(SUM[19]) );
  XOR2X1 U23 ( .IN1(n25), .IN2(A[18]), .Q(SUM[18]) );
  XOR2X1 U24 ( .IN1(n24), .IN2(A[17]), .Q(SUM[17]) );
  XOR2X1 U25 ( .IN1(n23), .IN2(A[16]), .Q(SUM[16]) );
  XOR2X1 U26 ( .IN1(n22), .IN2(A[15]), .Q(SUM[15]) );
  XOR2X1 U27 ( .IN1(n21), .IN2(A[14]), .Q(SUM[14]) );
  XOR2X1 U28 ( .IN1(n20), .IN2(A[13]), .Q(SUM[13]) );
  XOR2X1 U29 ( .IN1(n19), .IN2(A[12]), .Q(SUM[12]) );
  XOR2X1 U30 ( .IN1(n18), .IN2(A[11]), .Q(SUM[11]) );
  XOR2X1 U31 ( .IN1(n17), .IN2(A[10]), .Q(SUM[10]) );
  XOR2X1 U32 ( .IN1(n16), .IN2(A[9]), .Q(SUM[9]) );
  XOR2X1 U33 ( .IN1(n15), .IN2(A[8]), .Q(SUM[8]) );
  XOR2X1 U34 ( .IN1(n9), .IN2(A[30]), .Q(SUM[30]) );
  INVX0 U35 ( .IN(A[0]), .QN(SUM[0]) );
  XOR2X1 U36 ( .IN1(A[0]), .IN2(A[1]), .Q(SUM[1]) );
  XOR2X1 U37 ( .IN1(n14), .IN2(A[7]), .Q(SUM[7]) );
  XOR2X1 U38 ( .IN1(n13), .IN2(A[6]), .Q(SUM[6]) );
  XOR2X1 U39 ( .IN1(n11), .IN2(A[4]), .Q(SUM[4]) );
  XOR2X1 U40 ( .IN1(carry_3_), .IN2(A[3]), .Q(SUM[3]) );
  XOR2X1 U41 ( .IN1(n12), .IN2(A[5]), .Q(SUM[5]) );
  INVX0 U42 ( .IN(A[2]), .QN(n29) );
  AND2X1 U43 ( .IN1(A[0]), .IN2(A[1]), .Q(n10) );
  AND2X1 U44 ( .IN1(carry_3_), .IN2(A[3]), .Q(n11) );
  AND2X1 U45 ( .IN1(n11), .IN2(A[4]), .Q(n12) );
  AND2X1 U46 ( .IN1(n12), .IN2(A[5]), .Q(n13) );
  AND2X1 U47 ( .IN1(n13), .IN2(A[6]), .Q(n14) );
  AND2X1 U48 ( .IN1(n14), .IN2(A[7]), .Q(n15) );
  AND2X1 U49 ( .IN1(n15), .IN2(A[8]), .Q(n16) );
  AND2X1 U50 ( .IN1(n16), .IN2(A[9]), .Q(n17) );
  AND2X1 U51 ( .IN1(n17), .IN2(A[10]), .Q(n18) );
  AND2X1 U52 ( .IN1(n18), .IN2(A[11]), .Q(n19) );
  AND2X1 U53 ( .IN1(n19), .IN2(A[12]), .Q(n20) );
  AND2X1 U54 ( .IN1(n20), .IN2(A[13]), .Q(n21) );
  AND2X1 U55 ( .IN1(n21), .IN2(A[14]), .Q(n22) );
  AND2X1 U56 ( .IN1(n22), .IN2(A[15]), .Q(n23) );
  AND2X1 U57 ( .IN1(n23), .IN2(A[16]), .Q(n24) );
  AND2X1 U58 ( .IN1(n24), .IN2(A[17]), .Q(n25) );
  AND2X1 U59 ( .IN1(n25), .IN2(A[18]), .Q(n26) );
  AND2X1 U60 ( .IN1(n26), .IN2(A[19]), .Q(n27) );
  AND2X1 U61 ( .IN1(n27), .IN2(A[20]), .Q(n28) );
  XNOR2X1 U62 ( .IN1(n30), .IN2(A[31]), .Q(SUM[31]) );
  NAND2X0 U63 ( .IN1(n9), .IN2(A[30]), .QN(n30) );
endmodule


module b15_DW01_add_12 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29;
  assign SUM[0] = A[0];

  XOR2X1 U1 ( .IN1(A[1]), .IN2(A[2]), .Q(SUM[2]) );
  XOR2X1 U2 ( .IN1(n1), .IN2(A[3]), .Q(SUM[3]) );
  XOR2X1 U3 ( .IN1(n2), .IN2(A[4]), .Q(SUM[4]) );
  XOR2X1 U4 ( .IN1(n3), .IN2(A[5]), .Q(SUM[5]) );
  XOR2X1 U5 ( .IN1(n4), .IN2(A[6]), .Q(SUM[6]) );
  XOR2X1 U6 ( .IN1(n5), .IN2(A[7]), .Q(SUM[7]) );
  INVX0 U7 ( .IN(A[1]), .QN(SUM[1]) );
  AND2X1 U8 ( .IN1(A[1]), .IN2(A[2]), .Q(n1) );
  AND2X1 U9 ( .IN1(n1), .IN2(A[3]), .Q(n2) );
  AND2X1 U10 ( .IN1(n2), .IN2(A[4]), .Q(n3) );
  AND2X1 U11 ( .IN1(n3), .IN2(A[5]), .Q(n4) );
  AND2X1 U12 ( .IN1(n4), .IN2(A[6]), .Q(n5) );
  AND2X1 U13 ( .IN1(n28), .IN2(A[14]), .Q(n6) );
  AND2X1 U14 ( .IN1(n6), .IN2(A[15]), .Q(n7) );
  AND2X1 U15 ( .IN1(n7), .IN2(A[16]), .Q(n8) );
  AND2X1 U16 ( .IN1(n8), .IN2(A[17]), .Q(n9) );
  AND2X1 U17 ( .IN1(n9), .IN2(A[18]), .Q(n10) );
  AND2X1 U18 ( .IN1(n10), .IN2(A[19]), .Q(n11) );
  AND2X1 U19 ( .IN1(n11), .IN2(A[20]), .Q(n12) );
  AND2X1 U20 ( .IN1(n12), .IN2(A[21]), .Q(n13) );
  AND2X1 U21 ( .IN1(n13), .IN2(A[22]), .Q(n14) );
  AND2X1 U22 ( .IN1(n14), .IN2(A[23]), .Q(n15) );
  AND2X1 U23 ( .IN1(n15), .IN2(A[24]), .Q(n16) );
  AND2X1 U24 ( .IN1(n16), .IN2(A[25]), .Q(n17) );
  AND2X1 U25 ( .IN1(n17), .IN2(A[26]), .Q(n18) );
  AND2X1 U26 ( .IN1(n18), .IN2(A[27]), .Q(n19) );
  AND2X1 U27 ( .IN1(n19), .IN2(A[28]), .Q(n20) );
  AND2X1 U28 ( .IN1(n20), .IN2(A[29]), .Q(n21) );
  XOR2X1 U29 ( .IN1(n22), .IN2(A[8]), .Q(SUM[8]) );
  XOR2X1 U30 ( .IN1(n23), .IN2(A[9]), .Q(SUM[9]) );
  XOR2X1 U31 ( .IN1(n24), .IN2(A[10]), .Q(SUM[10]) );
  XOR2X1 U32 ( .IN1(n25), .IN2(A[11]), .Q(SUM[11]) );
  XOR2X1 U33 ( .IN1(n26), .IN2(A[12]), .Q(SUM[12]) );
  XOR2X1 U34 ( .IN1(n27), .IN2(A[13]), .Q(SUM[13]) );
  XOR2X1 U35 ( .IN1(n28), .IN2(A[14]), .Q(SUM[14]) );
  XOR2X1 U36 ( .IN1(n6), .IN2(A[15]), .Q(SUM[15]) );
  XOR2X1 U37 ( .IN1(n7), .IN2(A[16]), .Q(SUM[16]) );
  XOR2X1 U38 ( .IN1(n20), .IN2(A[29]), .Q(SUM[29]) );
  XOR2X1 U39 ( .IN1(n19), .IN2(A[28]), .Q(SUM[28]) );
  XOR2X1 U40 ( .IN1(n18), .IN2(A[27]), .Q(SUM[27]) );
  XOR2X1 U41 ( .IN1(n17), .IN2(A[26]), .Q(SUM[26]) );
  XOR2X1 U42 ( .IN1(n16), .IN2(A[25]), .Q(SUM[25]) );
  XOR2X1 U43 ( .IN1(n15), .IN2(A[24]), .Q(SUM[24]) );
  XOR2X1 U44 ( .IN1(n14), .IN2(A[23]), .Q(SUM[23]) );
  XOR2X1 U45 ( .IN1(n13), .IN2(A[22]), .Q(SUM[22]) );
  XOR2X1 U46 ( .IN1(n12), .IN2(A[21]), .Q(SUM[21]) );
  XOR2X1 U47 ( .IN1(n11), .IN2(A[20]), .Q(SUM[20]) );
  XOR2X1 U48 ( .IN1(n10), .IN2(A[19]), .Q(SUM[19]) );
  XOR2X1 U49 ( .IN1(n9), .IN2(A[18]), .Q(SUM[18]) );
  XOR2X1 U50 ( .IN1(n8), .IN2(A[17]), .Q(SUM[17]) );
  XOR2X1 U51 ( .IN1(n21), .IN2(A[30]), .Q(SUM[30]) );
  XNOR2X1 U52 ( .IN1(n29), .IN2(A[31]), .Q(SUM[31]) );
  NAND2X0 U53 ( .IN1(n21), .IN2(A[30]), .QN(n29) );
  AND2X1 U54 ( .IN1(n5), .IN2(A[7]), .Q(n22) );
  AND2X1 U55 ( .IN1(n22), .IN2(A[8]), .Q(n23) );
  AND2X1 U56 ( .IN1(n23), .IN2(A[9]), .Q(n24) );
  AND2X1 U57 ( .IN1(n24), .IN2(A[10]), .Q(n25) );
  AND2X1 U58 ( .IN1(n25), .IN2(A[11]), .Q(n26) );
  AND2X1 U59 ( .IN1(n26), .IN2(A[12]), .Q(n27) );
  AND2X1 U60 ( .IN1(n27), .IN2(A[13]), .Q(n28) );
endmodule


module b15_DW01_add_13 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29;
  assign SUM[0] = A[0];

  XOR2X1 U1 ( .IN1(n18), .IN2(A[5]), .Q(SUM[5]) );
  XOR2X1 U2 ( .IN1(n19), .IN2(A[3]), .Q(SUM[3]) );
  XOR2X1 U3 ( .IN1(A[1]), .IN2(A[2]), .Q(SUM[2]) );
  INVX0 U4 ( .IN(A[1]), .QN(SUM[1]) );
  XOR2X1 U5 ( .IN1(n17), .IN2(A[4]), .Q(SUM[4]) );
  AND2X1 U6 ( .IN1(n22), .IN2(A[23]), .Q(n1) );
  AND2X1 U7 ( .IN1(n18), .IN2(A[5]), .Q(n2) );
  AND2X1 U8 ( .IN1(n2), .IN2(A[6]), .Q(n3) );
  AND2X1 U9 ( .IN1(n3), .IN2(A[7]), .Q(n4) );
  AND2X1 U10 ( .IN1(n4), .IN2(A[8]), .Q(n5) );
  AND2X1 U11 ( .IN1(n5), .IN2(A[9]), .Q(n6) );
  AND2X1 U12 ( .IN1(n6), .IN2(A[10]), .Q(n7) );
  AND2X1 U13 ( .IN1(n7), .IN2(A[11]), .Q(n8) );
  AND2X1 U14 ( .IN1(n8), .IN2(A[12]), .Q(n9) );
  AND2X1 U15 ( .IN1(n9), .IN2(A[13]), .Q(n10) );
  AND2X1 U16 ( .IN1(n10), .IN2(A[14]), .Q(n11) );
  AND2X1 U17 ( .IN1(n11), .IN2(A[15]), .Q(n12) );
  AND2X1 U18 ( .IN1(n12), .IN2(A[16]), .Q(n13) );
  AND2X1 U19 ( .IN1(n13), .IN2(A[17]), .Q(n14) );
  AND2X1 U20 ( .IN1(n14), .IN2(A[18]), .Q(n15) );
  AND2X1 U21 ( .IN1(n15), .IN2(A[19]), .Q(n16) );
  AND2X1 U22 ( .IN1(n19), .IN2(A[3]), .Q(n17) );
  AND2X1 U23 ( .IN1(n17), .IN2(A[4]), .Q(n18) );
  XOR2X1 U24 ( .IN1(n27), .IN2(A[29]), .Q(SUM[29]) );
  XOR2X1 U25 ( .IN1(n26), .IN2(A[28]), .Q(SUM[28]) );
  XOR2X1 U26 ( .IN1(n25), .IN2(A[27]), .Q(SUM[27]) );
  XOR2X1 U27 ( .IN1(n24), .IN2(A[26]), .Q(SUM[26]) );
  XOR2X1 U28 ( .IN1(n23), .IN2(A[25]), .Q(SUM[25]) );
  XOR2X1 U29 ( .IN1(n1), .IN2(A[24]), .Q(SUM[24]) );
  XOR2X1 U30 ( .IN1(n22), .IN2(A[23]), .Q(SUM[23]) );
  XOR2X1 U31 ( .IN1(n21), .IN2(A[22]), .Q(SUM[22]) );
  XOR2X1 U32 ( .IN1(n20), .IN2(A[21]), .Q(SUM[21]) );
  XOR2X1 U33 ( .IN1(n16), .IN2(A[20]), .Q(SUM[20]) );
  XOR2X1 U34 ( .IN1(n28), .IN2(A[30]), .Q(SUM[30]) );
  XNOR2X1 U35 ( .IN1(n29), .IN2(A[31]), .Q(SUM[31]) );
  NAND2X0 U36 ( .IN1(n28), .IN2(A[30]), .QN(n29) );
  XOR2X1 U37 ( .IN1(n15), .IN2(A[19]), .Q(SUM[19]) );
  AND2X1 U38 ( .IN1(A[1]), .IN2(A[2]), .Q(n19) );
  AND2X1 U39 ( .IN1(n16), .IN2(A[20]), .Q(n20) );
  AND2X1 U40 ( .IN1(n20), .IN2(A[21]), .Q(n21) );
  AND2X1 U41 ( .IN1(n21), .IN2(A[22]), .Q(n22) );
  AND2X1 U42 ( .IN1(n1), .IN2(A[24]), .Q(n23) );
  AND2X1 U43 ( .IN1(n23), .IN2(A[25]), .Q(n24) );
  AND2X1 U44 ( .IN1(n24), .IN2(A[26]), .Q(n25) );
  AND2X1 U45 ( .IN1(n25), .IN2(A[27]), .Q(n26) );
  AND2X1 U46 ( .IN1(n26), .IN2(A[28]), .Q(n27) );
  AND2X1 U47 ( .IN1(n27), .IN2(A[29]), .Q(n28) );
  XOR2X1 U48 ( .IN1(n14), .IN2(A[18]), .Q(SUM[18]) );
  XOR2X1 U49 ( .IN1(n13), .IN2(A[17]), .Q(SUM[17]) );
  XOR2X1 U50 ( .IN1(n12), .IN2(A[16]), .Q(SUM[16]) );
  XOR2X1 U51 ( .IN1(n11), .IN2(A[15]), .Q(SUM[15]) );
  XOR2X1 U52 ( .IN1(n10), .IN2(A[14]), .Q(SUM[14]) );
  XOR2X1 U53 ( .IN1(n9), .IN2(A[13]), .Q(SUM[13]) );
  XOR2X1 U54 ( .IN1(n8), .IN2(A[12]), .Q(SUM[12]) );
  XOR2X1 U55 ( .IN1(n7), .IN2(A[11]), .Q(SUM[11]) );
  XOR2X1 U56 ( .IN1(n6), .IN2(A[10]), .Q(SUM[10]) );
  XOR2X1 U57 ( .IN1(n5), .IN2(A[9]), .Q(SUM[9]) );
  XOR2X1 U58 ( .IN1(n4), .IN2(A[8]), .Q(SUM[8]) );
  XOR2X1 U59 ( .IN1(n3), .IN2(A[7]), .Q(SUM[7]) );
  XOR2X1 U60 ( .IN1(n2), .IN2(A[6]), .Q(SUM[6]) );
endmodule


module b15_DW01_inc_3 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;

  wire   [31:2] carry;

  HADDX1 U1_1_30 ( .A0(A[30]), .B0(carry[30]), .C1(carry[31]), .SO(SUM[30]) );
  HADDX1 U1_1_17 ( .A0(A[17]), .B0(carry[17]), .C1(carry[18]), .SO(SUM[17]) );
  HADDX1 U1_1_18 ( .A0(A[18]), .B0(carry[18]), .C1(carry[19]), .SO(SUM[18]) );
  HADDX1 U1_1_19 ( .A0(A[19]), .B0(carry[19]), .C1(carry[20]), .SO(SUM[19]) );
  HADDX1 U1_1_20 ( .A0(A[20]), .B0(carry[20]), .C1(carry[21]), .SO(SUM[20]) );
  HADDX1 U1_1_21 ( .A0(A[21]), .B0(carry[21]), .C1(carry[22]), .SO(SUM[21]) );
  HADDX1 U1_1_22 ( .A0(A[22]), .B0(carry[22]), .C1(carry[23]), .SO(SUM[22]) );
  HADDX1 U1_1_23 ( .A0(A[23]), .B0(carry[23]), .C1(carry[24]), .SO(SUM[23]) );
  HADDX1 U1_1_24 ( .A0(A[24]), .B0(carry[24]), .C1(carry[25]), .SO(SUM[24]) );
  HADDX1 U1_1_25 ( .A0(A[25]), .B0(carry[25]), .C1(carry[26]), .SO(SUM[25]) );
  HADDX1 U1_1_26 ( .A0(A[26]), .B0(carry[26]), .C1(carry[27]), .SO(SUM[26]) );
  HADDX1 U1_1_27 ( .A0(A[27]), .B0(carry[27]), .C1(carry[28]), .SO(SUM[27]) );
  HADDX1 U1_1_28 ( .A0(A[28]), .B0(carry[28]), .C1(carry[29]), .SO(SUM[28]) );
  HADDX1 U1_1_29 ( .A0(A[29]), .B0(carry[29]), .C1(carry[30]), .SO(SUM[29]) );
  HADDX1 U1_1_16 ( .A0(A[16]), .B0(carry[16]), .C1(carry[17]), .SO(SUM[16]) );
  HADDX1 U1_1_15 ( .A0(A[15]), .B0(carry[15]), .C1(carry[16]), .SO(SUM[15]) );
  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .IN(A[0]), .QN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[31]), .IN2(A[31]), .Q(SUM[31]) );
endmodule


module b15_DW01_add_14 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29;
  assign SUM[0] = A[0];

  XOR2X1 U1 ( .IN1(n15), .IN2(A[4]), .Q(SUM[4]) );
  XOR2X1 U2 ( .IN1(A[1]), .IN2(A[2]), .Q(SUM[2]) );
  XOR2X1 U3 ( .IN1(n16), .IN2(A[5]), .Q(SUM[5]) );
  XOR2X1 U4 ( .IN1(n14), .IN2(A[3]), .Q(SUM[3]) );
  XOR2X1 U5 ( .IN1(n25), .IN2(A[14]), .Q(SUM[14]) );
  XOR2X1 U6 ( .IN1(n24), .IN2(A[13]), .Q(SUM[13]) );
  XOR2X1 U7 ( .IN1(n23), .IN2(A[12]), .Q(SUM[12]) );
  XOR2X1 U8 ( .IN1(n22), .IN2(A[11]), .Q(SUM[11]) );
  XOR2X1 U9 ( .IN1(n21), .IN2(A[10]), .Q(SUM[10]) );
  XOR2X1 U10 ( .IN1(n20), .IN2(A[9]), .Q(SUM[9]) );
  XOR2X1 U11 ( .IN1(n19), .IN2(A[8]), .Q(SUM[8]) );
  XOR2X1 U12 ( .IN1(n18), .IN2(A[7]), .Q(SUM[7]) );
  XOR2X1 U13 ( .IN1(n17), .IN2(A[6]), .Q(SUM[6]) );
  AND2X1 U14 ( .IN1(n25), .IN2(A[14]), .Q(n1) );
  AND2X1 U15 ( .IN1(n1), .IN2(A[15]), .Q(n2) );
  AND2X1 U16 ( .IN1(n26), .IN2(A[17]), .Q(n3) );
  AND2X1 U17 ( .IN1(n3), .IN2(A[18]), .Q(n4) );
  AND2X1 U18 ( .IN1(n4), .IN2(A[19]), .Q(n5) );
  AND2X1 U19 ( .IN1(n27), .IN2(A[21]), .Q(n6) );
  AND2X1 U20 ( .IN1(n6), .IN2(A[22]), .Q(n7) );
  AND2X1 U21 ( .IN1(n7), .IN2(A[23]), .Q(n8) );
  AND2X1 U22 ( .IN1(n28), .IN2(A[25]), .Q(n9) );
  AND2X1 U23 ( .IN1(n9), .IN2(A[26]), .Q(n10) );
  AND2X1 U24 ( .IN1(n10), .IN2(A[27]), .Q(n11) );
  AND2X1 U25 ( .IN1(n11), .IN2(A[28]), .Q(n12) );
  AND2X1 U26 ( .IN1(n12), .IN2(A[29]), .Q(n13) );
  AND2X1 U27 ( .IN1(A[1]), .IN2(A[2]), .Q(n14) );
  AND2X1 U28 ( .IN1(n14), .IN2(A[3]), .Q(n15) );
  AND2X1 U29 ( .IN1(n15), .IN2(A[4]), .Q(n16) );
  AND2X1 U30 ( .IN1(n16), .IN2(A[5]), .Q(n17) );
  AND2X1 U31 ( .IN1(n17), .IN2(A[6]), .Q(n18) );
  AND2X1 U32 ( .IN1(n18), .IN2(A[7]), .Q(n19) );
  AND2X1 U33 ( .IN1(n19), .IN2(A[8]), .Q(n20) );
  AND2X1 U34 ( .IN1(n20), .IN2(A[9]), .Q(n21) );
  AND2X1 U35 ( .IN1(n21), .IN2(A[10]), .Q(n22) );
  AND2X1 U36 ( .IN1(n22), .IN2(A[11]), .Q(n23) );
  AND2X1 U37 ( .IN1(n23), .IN2(A[12]), .Q(n24) );
  AND2X1 U38 ( .IN1(n24), .IN2(A[13]), .Q(n25) );
  AND2X1 U39 ( .IN1(n2), .IN2(A[16]), .Q(n26) );
  AND2X1 U40 ( .IN1(n5), .IN2(A[20]), .Q(n27) );
  AND2X1 U41 ( .IN1(n8), .IN2(A[24]), .Q(n28) );
  XNOR2X1 U42 ( .IN1(n29), .IN2(A[31]), .Q(SUM[31]) );
  NAND2X0 U43 ( .IN1(n13), .IN2(A[30]), .QN(n29) );
  XOR2X1 U44 ( .IN1(n11), .IN2(A[28]), .Q(SUM[28]) );
  XOR2X1 U45 ( .IN1(n10), .IN2(A[27]), .Q(SUM[27]) );
  XOR2X1 U46 ( .IN1(n9), .IN2(A[26]), .Q(SUM[26]) );
  XOR2X1 U47 ( .IN1(n28), .IN2(A[25]), .Q(SUM[25]) );
  XOR2X1 U48 ( .IN1(n8), .IN2(A[24]), .Q(SUM[24]) );
  XOR2X1 U49 ( .IN1(n7), .IN2(A[23]), .Q(SUM[23]) );
  XOR2X1 U50 ( .IN1(n6), .IN2(A[22]), .Q(SUM[22]) );
  XOR2X1 U51 ( .IN1(n27), .IN2(A[21]), .Q(SUM[21]) );
  XOR2X1 U52 ( .IN1(n5), .IN2(A[20]), .Q(SUM[20]) );
  XOR2X1 U53 ( .IN1(n12), .IN2(A[29]), .Q(SUM[29]) );
  XOR2X1 U54 ( .IN1(n13), .IN2(A[30]), .Q(SUM[30]) );
  XOR2X1 U55 ( .IN1(n4), .IN2(A[19]), .Q(SUM[19]) );
  XOR2X1 U56 ( .IN1(n3), .IN2(A[18]), .Q(SUM[18]) );
  XOR2X1 U57 ( .IN1(n26), .IN2(A[17]), .Q(SUM[17]) );
  XOR2X1 U58 ( .IN1(n2), .IN2(A[16]), .Q(SUM[16]) );
  XOR2X1 U59 ( .IN1(n1), .IN2(A[15]), .Q(SUM[15]) );
  INVX0 U60 ( .IN(A[1]), .QN(SUM[1]) );
endmodule


module b15_DW01_add_21 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   carry_9_, carry_31_, carry_30_, carry_29_, carry_28_, carry_27_,
         carry_26_, carry_25_, carry_24_, carry_23_, carry_22_, carry_21_,
         carry_20_, carry_19_, carry_18_, carry_17_, carry_16_, carry_15_,
         carry_14_, carry_13_, carry_12_, carry_11_, carry_10_, n1;
  wire   [8:2] carry;

  XOR3X1 U1_31 ( .IN1(A[31]), .IN2(B[31]), .IN3(carry_31_), .Q(SUM[31]) );
  FADDX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  FADDX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry_29_), .CO(carry_30_), .S(
        SUM[29]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry_27_), .CO(carry_28_), .S(
        SUM[27]) );
  FADDX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry_25_), .CO(carry_26_), .S(
        SUM[25]) );
  FADDX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry_23_), .CO(carry_24_), .S(
        SUM[23]) );
  FADDX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry_22_), .CO(carry_23_), .S(
        SUM[22]) );
  FADDX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry_21_), .CO(carry_22_), .S(
        SUM[21]) );
  FADDX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry_20_), .CO(carry_21_), .S(
        SUM[20]) );
  FADDX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry_19_), .CO(carry_20_), .S(
        SUM[19]) );
  FADDX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry_18_), .CO(carry_19_), .S(
        SUM[18]) );
  FADDX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry_17_), .CO(carry_18_), .S(
        SUM[17]) );
  FADDX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry_16_), .CO(carry_17_), .S(
        SUM[16]) );
  FADDX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry_15_), .CO(carry_16_), .S(
        SUM[15]) );
  FADDX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry_14_), .CO(carry_15_), .S(
        SUM[14]) );
  FADDX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry_13_), .CO(carry_14_), .S(
        SUM[13]) );
  FADDX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry_12_), .CO(carry_13_), .S(
        SUM[12]) );
  FADDX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry_11_), .CO(carry_12_), .S(
        SUM[11]) );
  FADDX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry_10_), .CO(carry_11_), .S(
        SUM[10]) );
  FADDX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry_9_), .CO(carry_10_), .S(SUM[9])
         );
  FADDX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry_9_), .S(SUM[8])
         );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry_30_), .CO(carry_31_), .S(
        SUM[30]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry_28_), .CO(carry_29_), .S(
        SUM[28]) );
  FADDX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry_26_), .CO(carry_27_), .S(
        SUM[26]) );
  FADDX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry_24_), .CO(carry_25_), .S(
        SUM[24]) );
  FADDX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2X1 U1 ( .IN1(B[0]), .IN2(A[0]), .Q(n1) );
  XOR2X1 U2 ( .IN1(B[0]), .IN2(A[0]), .Q(SUM[0]) );
endmodule


module b15 ( BE_n, Address, W_R_n, D_C_n, M_IO_n, ADS_n, Datai, Datao, CLOCK, 
        NA_n, BS16_n, READY_n, HOLD, RESET, test_se, test_si1, test_so1, 
        test_si2, test_so2, test_si3, test_so3, test_si4, test_so4, test_si5, 
        test_so5, test_si6, test_so6, test_si7, test_so7, test_si8, test_so8, 
        test_si9, test_so9, test_si10, test_so10, test_si11, test_so11, 
        test_si12, test_so12, test_si13, test_so13, test_si14, test_so14, 
        test_si15, test_so15, test_si16, test_so16, test_si17, test_so17, 
        test_si18, test_so18, test_si19, test_so19, test_si20, test_so20 );
  output [3:0] BE_n;
  output [29:0] Address;
  input [31:0] Datai;
  output [31:0] Datao;
  input CLOCK, NA_n, BS16_n, READY_n, HOLD, RESET, test_se, test_si1, test_si2,
         test_si3, test_si4, test_si5, test_si6, test_si7, test_si8, test_si9,
         test_si10, test_si11, test_si12, test_si13, test_si14, test_si15,
         test_si16, test_si17, test_si18, test_si19, test_si20;
  output W_R_n, D_C_n, M_IO_n, ADS_n, test_so1, test_so2, test_so3, test_so4,
         test_so5, test_so6, test_so7, test_so8, test_so9, test_so10,
         test_so11, test_so12, test_so13, test_so14, test_so15, test_so16,
         test_so17, test_so18, test_so19, test_so20;
  wire   rEIP_31_, rEIP_30_, rEIP_29_, rEIP_28_, rEIP_27_, rEIP_25_, rEIP_24_,
         rEIP_23_, rEIP_22_, rEIP_21_, rEIP_20_, rEIP_19_, rEIP_18_, rEIP_17_,
         rEIP_16_, rEIP_15_, rEIP_14_, rEIP_13_, rEIP_12_, rEIP_11_, rEIP_10_,
         rEIP_9_, rEIP_8_, rEIP_7_, rEIP_5_, rEIP_4_, rEIP_3_, rEIP_2_,
         rEIP_1_, rEIP_0_, N425, N426, N427, N428, N429, N430, N431, N432,
         N433, N434, N435, N436, N437, N438, N439, N440, N441, N442, N443,
         N444, N445, N446, N447, N448, N449, N450, N451, N452, N453, N454,
         N455, N498, N499, N500, N501, N502, N503, N504, N505, N506, N507,
         N508, N509, N510, N511, N512, N513, N514, N515, N516, N517, N518,
         N519, N520, N521, N522, N523, N524, N525, N526, N527, N528,
         InstAddrPointer_30_, InstAddrPointer_29_, InstAddrPointer_27_,
         InstAddrPointer_26_, InstAddrPointer_25_, InstAddrPointer_24_,
         InstAddrPointer_23_, InstAddrPointer_22_, InstAddrPointer_21_,
         InstAddrPointer_20_, InstAddrPointer_19_, InstAddrPointer_18_,
         InstAddrPointer_17_, InstAddrPointer_16_, InstAddrPointer_15_,
         InstAddrPointer_14_, InstAddrPointer_13_, InstAddrPointer_12_,
         InstAddrPointer_11_, InstAddrPointer_10_, InstAddrPointer_9_,
         InstAddrPointer_8_, InstAddrPointer_6_, InstAddrPointer_5_,
         InstAddrPointer_4_, InstAddrPointer_3_, InstAddrPointer_2_,
         InstAddrPointer_1_, PhyAddrPointer_31_, PhyAddrPointer_30_,
         PhyAddrPointer_29_, PhyAddrPointer_28_, PhyAddrPointer_27_,
         PhyAddrPointer_26_, PhyAddrPointer_25_, PhyAddrPointer_23_,
         PhyAddrPointer_22_, PhyAddrPointer_21_, PhyAddrPointer_20_,
         PhyAddrPointer_19_, PhyAddrPointer_18_, PhyAddrPointer_17_,
         PhyAddrPointer_16_, PhyAddrPointer_15_, PhyAddrPointer_14_,
         PhyAddrPointer_13_, PhyAddrPointer_12_, PhyAddrPointer_11_,
         PhyAddrPointer_10_, PhyAddrPointer_9_, PhyAddrPointer_8_,
         PhyAddrPointer_7_, PhyAddrPointer_6_, PhyAddrPointer_5_,
         PhyAddrPointer_4_, PhyAddrPointer_2_, PhyAddrPointer_1_,
         PhyAddrPointer_0_, EAX_31_, EAX_29_, EAX_28_, EAX_27_, EAX_26_,
         EAX_25_, EAX_24_, EAX_23_, EAX_22_, EAX_21_, EAX_20_, EAX_19_,
         EAX_18_, EAX_17_, EAX_16_, EBX_30_, EBX_29_, EBX_28_, EBX_27_,
         EBX_26_, EBX_25_, EBX_24_, EBX_23_, EBX_22_, EBX_21_, EBX_20_,
         EBX_18_, EBX_17_, EBX_16_, EBX_15_, EBX_14_, EBX_13_, EBX_12_,
         EBX_11_, EBX_10_, EBX_9_, EBX_8_, EBX_7_, EBX_6_, EBX_5_, EBX_4_,
         EBX_3_, EBX_2_, EBX_1_, EBX_0_, N651, N652, N653, N654, N655, N656,
         N657, N811, N964, N965, N966, N967, N968, N969, N970, N971, N972,
         N973, N974, N975, N976, N977, N978, N979, N980, N981, N982, N983,
         N984, N985, N986, N987, N988, N989, N990, N991, N992, N993, N994,
         N995, N997, N998, N999, N1000, N1001, N1002, N1003, N1004, N1005,
         N1006, N1007, N1008, N1009, N1010, N1011, N1012, N1013, N1014, N1015,
         N1016, N1017, N1018, N1019, N1020, N1021, N1022, N1023, N1024, N1025,
         N1026, N1027, N1029, N1031, N1032, N1033, N1034, N1035, N1036, N1037,
         N1038, N1039, N1040, N1041, N1042, N1043, N1044, N1045, N1046, N1047,
         N1048, N1049, N1050, N1051, N1052, N1053, N1054, N1055, N1056, N1057,
         N1058, N1059, N1060, N1061, N1062, N1239, N1479, N1480, N1481, N1482,
         N1483, N1484, N1485, N1486, N1487, N1488, N1489, N1490, N1491, N1492,
         N1493, N1494, N1495, N1496, N1497, N1498, N1499, N1500, N1501, N1502,
         N1503, N1504, N1505, N1506, N1507, N1508, N1509, N1510, N1551, N1552,
         N1553, N1554, N1555, N1556, N1557, N1558, N1559, N1560, N1561, N1562,
         N1563, N1564, N1565, N1566, N1567, N1568, N1569, N1570, N1571, N1572,
         N1573, N1574, N1575, N1576, N1577, N1578, N1579, N1580, N1581, N1582,
         N1619, N1620, N1621, N1622, N1623, N1624, N1625, N1626, N1627, N1628,
         N1629, N1630, N1631, N1632, N1633, N1634, N1635, N1636, N1637, N1638,
         N1639, N1640, N1641, N1642, N1643, N1644, N1645, N1646, N1647, N1648,
         N1649, N1650, N1749, N1750, N1751, N1752, N1753, N1754, N1755, N1756,
         N1757, N1758, N1759, N1760, N1761, N1762, N1763, N1764, N1769, N1770,
         N1771, N1772, N1773, N1774, N1775, N1776, N1777, N1778, N1779, N1780,
         N1781, N1782, N1783, N1784, N1785, N1786, N1787, N1788, N1789, N1790,
         N1791, N1792, N1793, N1794, N1795, N1796, N1797, N1798, N1799, N1800,
         N1954, N1956, N1957, N1958, N1959, N1960, N1961, N1962, N1963, N1964,
         N1965, N1966, N1967, N1968, N1969, N1970, N1971, N1972, N1973, N1974,
         N1975, N1976, N1977, N1978, N1979, N1980, N1981, N1982, N1983, N1984,
         N1985, N1986, N1987, N2103, N2104, N2105, N2106, N2107, N2108, N2109,
         N2110, N2111, N2112, N2113, N2114, N2115, N2116, N2117, N2118, N2385,
         N2386, N2387, N2388, N2389, N2390, N2391, N2392, N2393, N2394, N2395,
         N2396, N2397, N2398, N2399, N2400, N2401, N2402, N2403, N2404, N2405,
         N2406, N2407, N2408, N2409, N2410, N2411, N2412, N2413, N2414, N2415,
         N2416, N2417, N2418, N2419, N2420, N2421, N2422, N2423, N2424, N2425,
         N2426, N2427, N2428, N2429, N2430, N2431, N2432, N2433, N2434, N2435,
         N2436, N2437, N2438, N2439, N2440, N2441, N2442, N2443, N2444, N2445,
         N2446, N2447, N2548, N2549, N2550, N2551, N2552, N2553, N2554, N2555,
         N2571, N2572, N2573, N2574, N2575, N2576, N2577, N2578, N2700, N2701,
         N2702, N2703, N2704, N2737, N2739, N2740, N2856, N2857, N2858, N2859,
         N2860, N2861, N2862, N2863, N2864, N2865, N2866, N2867, N2868, N2869,
         N2870, N2871, N2872, N2873, N2874, N2875, N2876, N2877, N2878, N2879,
         N2880, N2881, N2882, N2883, N2884, N2885, N2886, N2887, N2995, N2996,
         N2997, N2998, N2999, N3000, N3001, N3002, N3003, N3004, N3005, N3006,
         N3007, N3008, N3009, N3010, N3011, N3012, N3013, N3014, N3015, N3016,
         N3017, N3018, N3019, N3020, N3021, N3022, N3023, N3024, N3025, N3026,
         N3067, N3068, N3069, N3070, N3071, N3072, N3073, N3074, N3075, N3076,
         N3077, N3078, N3079, N3080, N3081, N3082, N3083, N3084, N3085, N3086,
         N3087, N3088, N3089, N3090, N3091, N3092, N3093, N3094, N3095, N3096,
         N3097, N3098, N3346, N3347, N3348, N3349, N3350, N3351, N3352, N3353,
         N3354, N3356, N3357, N3358, N3359, N3360, N3361, N3415, N3417, N3418,
         N3419, N3420, N3423, N3424, N3427, N3428, N3434, N3435, N3437, N3438,
         N3439, N3440, N3441, N3442, N3443, N3444, N3445, N3446, N3447, N3448,
         N3449, N3450, N3451, N3452, N3453, N3454, N3455, N3456, N3457, N3458,
         N3459, N3460, N3461, N3462, N3463, N3467, N3469, N3484, N3485, N3486,
         N3493, N3494, N3989, N3990, N3991, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n1415, n1416,
         n1434, n1435, n1436, n1472, n1490, n1491, n1492, n1548, n1550, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1595, n1596,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, r680_B_1_, r680_B_2_,
         r680_B_3_, r680_B_4_, gte_355_B_0_, add_div_311_A_0_,
         add_1_root_add_0_root_add_402_7_B_23_,
         add_1_root_add_0_root_add_402_7_B_24_,
         add_1_root_add_0_root_add_402_7_B_25_,
         add_1_root_add_0_root_add_402_7_B_26_,
         add_1_root_add_0_root_add_402_7_B_27_,
         add_1_root_add_0_root_add_402_7_B_28_,
         add_1_root_add_0_root_add_402_7_B_29_,
         add_1_root_add_0_root_add_402_7_B_30_,
         add_1_root_add_0_root_add_402_7_A_23_,
         add_2_root_sub_1_root_sub_357_2_SUM_2_,
         add_2_root_sub_1_root_sub_357_2_SUM_3_,
         add_2_root_sub_1_root_sub_357_2_SUM_4_,
         add_2_root_sub_1_root_sub_357_2_SUM_5_,
         add_2_root_sub_1_root_sub_357_2_SUM_6_,
         add_2_root_sub_1_root_sub_357_2_SUM_7_, mult_add_463_aco_A_0_, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2886, n2887, n2888, n2889, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5326;
  wire   [4:1] InstQueueRd_Addr;
  wire   [4:3] add_495_carry;
  wire   [14:1] add_div_457_carry;
  wire   [7:1] add_div_313_carry;
  wire   [6:1] add_div_311_carry;
  wire   [4:2] r698_carry;
  wire   [4:1] r679_carry;
  wire   [30:24] add_1_root_add_0_root_add_402_7_carry;
  wire   [30:24] add_1_root_add_0_root_add_391_7_carry;
  wire   [7:3] add_2_root_sub_1_root_sub_357_2_carry;
  assign test_so1 = Address[19];
  assign Datao[31] = 1'b0;
  assign test_so3 = Datao[19];

  b15_DW01_add_1 add_0_root_add_360_3 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N2392, N2391, N2390, N2389, N2388, 
        N2387, N2386, N2385}), .B({n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63, n64, n65}), .CI(1'b0), .SUM({N3098, 
        N3097, N3096, N3095, N3094, N3093, N3092, N3091, N3090, N3089, N3088, 
        N3087, N3086, N3085, N3084, N3083, N3082, N3081, N3080, N3079, N3078, 
        N3077, N3076, N3075, N3074, N3073, N3072, N3071, N3070, N3069, N3068, 
        N3067}), .CO() );
  b15_DW01_add_2 add_0_root_add_371_3 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N2392, N2391, N2390, N2389, N2388, 
        N2387, N2386, N2385}), .B({N2447, N2446, N2445, N2444, N2443, N2442, 
        N2441, N2440, N2439, N2438, N2437, N2436, N2435, N2434, N2433, N2432, 
        N2431, N2430, N2429, N2428, N2427, N2426, N2425, N2424, N2423, N2422, 
        N2421, N2420, N2419, N2418, N2417, N2416}), .CI(1'b0), .SUM({N2887, 
        N2886, N2885, N2884, N2883, N2882, N2881, N2880, N2879, N2878, N2877, 
        N2876, N2875, N2874, N2873, N2872, N2871, N2870, N2869, N2868, N2867, 
        N2866, N2865, N2864, N2863, N2862, N2861, N2860, N2859, N2858, N2857, 
        N2856}), .CO() );
  b15_DW01_sub_2 sub_414 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({N1954, EBX_30_, EBX_29_, EBX_28_, EBX_27_, EBX_26_, EBX_25_, EBX_24_, 
        EBX_23_, EBX_22_, EBX_21_, EBX_20_, test_so6, EBX_18_, EBX_17_, 
        EBX_16_, EBX_15_, EBX_14_, EBX_13_, EBX_12_, EBX_11_, EBX_10_, EBX_9_, 
        EBX_8_, EBX_7_, EBX_6_, EBX_5_, EBX_4_, EBX_3_, EBX_2_, EBX_1_, EBX_0_}), .CI(1'b0), .DIFF({N1987, N1986, N1985, N1984, N1983, N1982, N1981, N1980, 
        N1979, N1978, N1977, N1976, N1975, N1974, N1973, N1972, N1971, N1970, 
        N1969, N1968, N1967, N1966, N1965, N1964, N1963, N1962, N1961, N1960, 
        N1959, N1958, N1957, N1956}), .CO() );
  b15_DW01_inc_0 add_552 ( .A({N1954, EBX_30_, EBX_29_, EBX_28_, EBX_27_, 
        EBX_26_, EBX_25_, EBX_24_, EBX_23_, EBX_22_, EBX_21_, EBX_20_, 
        test_so6, EBX_18_, EBX_17_, EBX_16_, EBX_15_, EBX_14_, EBX_13_, 
        EBX_12_, EBX_11_, EBX_10_, EBX_9_, EBX_8_, EBX_7_, EBX_6_, EBX_5_, 
        EBX_4_, EBX_3_, EBX_2_, EBX_1_, EBX_0_}), .SUM({N1650, N1649, N1648, 
        N1647, N1646, N1645, N1644, N1643, N1642, N1641, N1640, N1639, N1638, 
        N1637, N1636, N1635, N1634, N1633, N1632, N1631, N1630, N1629, N1628, 
        N1627, N1626, N1625, N1624, N1623, N1622, N1621, N1620, N1619}) );
  b15_DW01_inc_1 add_546 ( .A({EAX_31_, test_so5, EAX_29_, EAX_28_, EAX_27_, 
        EAX_26_, EAX_25_, EAX_24_, EAX_23_, EAX_22_, EAX_21_, EAX_20_, EAX_19_, 
        EAX_18_, EAX_17_, EAX_16_, N3361, N3360, N3359, N3358, N3357, N3356, 
        test_so4, N3354, N3353, N3352, N3351, N3350, N3349, N3348, N3347, 
        N3346}), .SUM({N1582, N1581, N1580, N1579, N1578, N1577, N1576, N1575, 
        N1574, N1573, N1572, N1571, N1570, N1569, N1568, N1567, N1566, N1565, 
        N1564, N1563, N1562, N1561, N1560, N1559, N1558, N1557, N1556, N1555, 
        N1554, N1553, N1552, N1551}) );
  b15_DW01_sub_3 sub_320 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({N1029, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, 
        N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, 
        N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, 
        N998, N997}), .CI(1'b0), .DIFF({N1062, N1061, N1060, N1059, N1058, 
        N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, 
        N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, 
        N1037, N1036, N1035, N1034, N1033, N1032, N1031}), .CO() );
  b15_DW01_add_6 add_315 ( .A({PhyAddrPointer_31_, PhyAddrPointer_30_, 
        PhyAddrPointer_29_, PhyAddrPointer_28_, PhyAddrPointer_27_, 
        PhyAddrPointer_26_, PhyAddrPointer_25_, test_so16, PhyAddrPointer_23_, 
        PhyAddrPointer_22_, PhyAddrPointer_21_, PhyAddrPointer_20_, 
        PhyAddrPointer_19_, PhyAddrPointer_18_, PhyAddrPointer_17_, 
        PhyAddrPointer_16_, PhyAddrPointer_15_, PhyAddrPointer_14_, 
        PhyAddrPointer_13_, PhyAddrPointer_12_, PhyAddrPointer_11_, 
        PhyAddrPointer_10_, PhyAddrPointer_9_, PhyAddrPointer_8_, 
        PhyAddrPointer_7_, PhyAddrPointer_6_, PhyAddrPointer_5_, 
        PhyAddrPointer_4_, test_so15, PhyAddrPointer_2_, PhyAddrPointer_1_, 
        PhyAddrPointer_0_}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 
        1'b0}), .CI(1'b0), .SUM({N995, N994, N993, N992, N991, N990, N989, 
        N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, 
        N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, 
        N964}), .CO() );
  b15_DW01_add_9 add_div_197 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N498}), 
        .B({rEIP_30_, rEIP_29_, rEIP_28_, rEIP_27_, test_so19, rEIP_25_, 
        rEIP_24_, rEIP_23_, rEIP_22_, rEIP_21_, rEIP_20_, rEIP_19_, rEIP_18_, 
        rEIP_17_, rEIP_16_, rEIP_15_, rEIP_14_, rEIP_13_, rEIP_12_, rEIP_11_, 
        rEIP_10_, rEIP_9_, rEIP_8_, rEIP_7_, test_so18, rEIP_5_, rEIP_4_, 
        rEIP_3_, rEIP_2_, rEIP_1_}), .CI(1'b0), .SUM({N528, N527, N526, N525, 
        N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, 
        N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, 
        N500, N499}), .CO() );
  b15_DW01_add_10 add_div_125 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N425}), 
        .B({rEIP_31_, rEIP_30_, rEIP_29_, rEIP_28_, rEIP_27_, test_so19, 
        rEIP_25_, rEIP_24_, rEIP_23_, rEIP_22_, rEIP_21_, rEIP_20_, rEIP_19_, 
        rEIP_18_, rEIP_17_, rEIP_16_, rEIP_15_, rEIP_14_, rEIP_13_, rEIP_12_, 
        rEIP_11_, rEIP_10_, rEIP_9_, rEIP_8_, rEIP_7_, test_so18, rEIP_5_, 
        rEIP_4_, rEIP_3_, rEIP_2_}), .CI(1'b0), .SUM({N455, N454, N453, N452, 
        N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, 
        N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, 
        N427, N426}), .CO() );
  b15_DW01_add_11 r693 ( .A({N3467, InstAddrPointer_30_, InstAddrPointer_29_, 
        test_so8, InstAddrPointer_27_, InstAddrPointer_26_, 
        InstAddrPointer_25_, InstAddrPointer_24_, InstAddrPointer_23_, 
        InstAddrPointer_22_, InstAddrPointer_21_, InstAddrPointer_20_, 
        InstAddrPointer_19_, InstAddrPointer_18_, InstAddrPointer_17_, 
        InstAddrPointer_16_, InstAddrPointer_15_, InstAddrPointer_14_, 
        InstAddrPointer_13_, InstAddrPointer_12_, InstAddrPointer_11_, 
        InstAddrPointer_10_, InstAddrPointer_9_, InstAddrPointer_8_, test_so7, 
        InstAddrPointer_6_, InstAddrPointer_5_, InstAddrPointer_4_, 
        InstAddrPointer_3_, InstAddrPointer_2_, InstAddrPointer_1_, N3469}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1}), .CI(1'b0), 
        .SUM({N2447, N2446, N2445, N2444, N2443, N2442, N2441, N2440, N2439, 
        N2438, N2437, N2436, N2435, N2434, N2433, N2432, N2431, N2430, N2429, 
        N2428, N2427, N2426, N2425, N2424, N2423, N2422, N2421, N2420, N2419, 
        N2418, N2417, N2416}), .CO() );
  b15_DW01_add_12 r684 ( .A({N3467, InstAddrPointer_30_, InstAddrPointer_29_, 
        test_so8, InstAddrPointer_27_, InstAddrPointer_26_, 
        InstAddrPointer_25_, InstAddrPointer_24_, InstAddrPointer_23_, 
        InstAddrPointer_22_, InstAddrPointer_21_, InstAddrPointer_20_, 
        InstAddrPointer_19_, InstAddrPointer_18_, InstAddrPointer_17_, 
        InstAddrPointer_16_, InstAddrPointer_15_, InstAddrPointer_14_, 
        InstAddrPointer_13_, InstAddrPointer_12_, InstAddrPointer_11_, 
        InstAddrPointer_10_, InstAddrPointer_9_, InstAddrPointer_8_, test_so7, 
        InstAddrPointer_6_, InstAddrPointer_5_, InstAddrPointer_4_, 
        InstAddrPointer_3_, InstAddrPointer_2_, InstAddrPointer_1_, N3469}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0}), .CI(1'b0), 
        .SUM({n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, 
        n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, 
        n61, n62, n63, n64, n65}), .CO() );
  b15_DW01_add_13 r683 ( .A({rEIP_31_, rEIP_30_, rEIP_29_, rEIP_28_, rEIP_27_, 
        test_so19, rEIP_25_, rEIP_24_, rEIP_23_, rEIP_22_, rEIP_21_, rEIP_20_, 
        rEIP_19_, rEIP_18_, rEIP_17_, rEIP_16_, rEIP_15_, rEIP_14_, rEIP_13_, 
        rEIP_12_, rEIP_11_, rEIP_10_, rEIP_9_, rEIP_8_, rEIP_7_, test_so18, 
        rEIP_5_, rEIP_4_, rEIP_3_, rEIP_2_, rEIP_1_, rEIP_0_}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0}), .CI(1'b0), .SUM({N1800, N1799, 
        N1798, N1797, N1796, N1795, N1794, N1793, N1792, N1791, N1790, N1789, 
        N1788, N1787, N1786, N1785, N1784, N1783, N1782, N1781, N1780, N1779, 
        N1778, N1777, N1776, N1775, N1774, N1773, N1772, N1771, N1770, N1769}), 
        .CO() );
  b15_DW01_inc_3 r675 ( .A({N3467, InstAddrPointer_30_, InstAddrPointer_29_, 
        test_so8, InstAddrPointer_27_, InstAddrPointer_26_, 
        InstAddrPointer_25_, InstAddrPointer_24_, InstAddrPointer_23_, 
        InstAddrPointer_22_, InstAddrPointer_21_, InstAddrPointer_20_, 
        InstAddrPointer_19_, InstAddrPointer_18_, InstAddrPointer_17_, 
        InstAddrPointer_16_, InstAddrPointer_15_, InstAddrPointer_14_, 
        InstAddrPointer_13_, InstAddrPointer_12_, InstAddrPointer_11_, 
        InstAddrPointer_10_, InstAddrPointer_9_, InstAddrPointer_8_, test_so7, 
        InstAddrPointer_6_, InstAddrPointer_5_, InstAddrPointer_4_, 
        InstAddrPointer_3_, InstAddrPointer_2_, InstAddrPointer_1_, N3469}), 
        .SUM({N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, 
        N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, 
        N1491, N1490, N1489, N1488, N1487, N1486, N1485, N1484, N1483, N1482, 
        N1481, N1480, N1479}) );
  b15_DW01_add_14 r672 ( .A({PhyAddrPointer_31_, PhyAddrPointer_30_, 
        PhyAddrPointer_29_, PhyAddrPointer_28_, PhyAddrPointer_27_, 
        PhyAddrPointer_26_, PhyAddrPointer_25_, test_so16, PhyAddrPointer_23_, 
        PhyAddrPointer_22_, PhyAddrPointer_21_, PhyAddrPointer_20_, 
        PhyAddrPointer_19_, PhyAddrPointer_18_, PhyAddrPointer_17_, 
        PhyAddrPointer_16_, PhyAddrPointer_15_, PhyAddrPointer_14_, 
        PhyAddrPointer_13_, PhyAddrPointer_12_, PhyAddrPointer_11_, 
        PhyAddrPointer_10_, PhyAddrPointer_9_, PhyAddrPointer_8_, 
        PhyAddrPointer_7_, PhyAddrPointer_6_, PhyAddrPointer_5_, 
        PhyAddrPointer_4_, test_so15, PhyAddrPointer_2_, PhyAddrPointer_1_, 
        PhyAddrPointer_0_}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 
        1'b0}), .CI(1'b0), .SUM({N1029, N1027, N1026, N1025, N1024, N1023, 
        N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, 
        N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, 
        N1002, N1001, N1000, N999, N998, N997}), .CO() );
  b15_DW01_add_21 add_0_root_sub_1_root_sub_357_2 ( .A({N3467, 
        InstAddrPointer_30_, InstAddrPointer_29_, test_so8, 
        InstAddrPointer_27_, InstAddrPointer_26_, InstAddrPointer_25_, 
        InstAddrPointer_24_, InstAddrPointer_23_, InstAddrPointer_22_, 
        InstAddrPointer_21_, InstAddrPointer_20_, InstAddrPointer_19_, 
        InstAddrPointer_18_, InstAddrPointer_17_, InstAddrPointer_16_, 
        InstAddrPointer_15_, InstAddrPointer_14_, InstAddrPointer_13_, 
        InstAddrPointer_12_, InstAddrPointer_11_, InstAddrPointer_10_, 
        InstAddrPointer_9_, InstAddrPointer_8_, test_so7, InstAddrPointer_6_, 
        InstAddrPointer_5_, InstAddrPointer_4_, InstAddrPointer_3_, 
        InstAddrPointer_2_, InstAddrPointer_1_, N3469}), .B({n3679, n3681, 
        n3679, n3681, n3679, n3681, n3679, n3681, n3679, n3680, n3679, n3680, 
        n3679, n3680, n3679, n3680, n3679, n3680, n3679, n3680, n3680, n3680, 
        n3680, n3680, add_2_root_sub_1_root_sub_357_2_SUM_7_, 
        add_2_root_sub_1_root_sub_357_2_SUM_6_, 
        add_2_root_sub_1_root_sub_357_2_SUM_5_, 
        add_2_root_sub_1_root_sub_357_2_SUM_4_, 
        add_2_root_sub_1_root_sub_357_2_SUM_3_, 
        add_2_root_sub_1_root_sub_357_2_SUM_2_, n5316, N2385}), .CI(1'b0), 
        .SUM({N3026, N3025, N3024, N3023, N3022, N3021, N3020, N3019, N3018, 
        N3017, N3016, N3015, N3014, N3013, N3012, N3011, N3010, N3009, N3008, 
        N3007, N3006, N3005, N3004, N3003, N3002, N3001, N3000, N2999, N2998, 
        N2997, N2996, N2995}), .CO() );
  SDFFARX1 uWord_reg_0_ ( .D(n2541), .SI(rEIP_31_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3572), .Q(N3450), .QN() );
  SDFFARX1 uWord_reg_1_ ( .D(n2540), .SI(N3450), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3572), .Q(N3451), .QN() );
  SDFFARX1 uWord_reg_2_ ( .D(n2539), .SI(N3451), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3571), .Q(N3452), .QN() );
  SDFFARX1 uWord_reg_3_ ( .D(n2538), .SI(N3452), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3571), .Q(N3453), .QN() );
  SDFFARX1 uWord_reg_4_ ( .D(n2537), .SI(N3453), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3571), .Q(N3454), .QN() );
  SDFFARX1 uWord_reg_5_ ( .D(n2536), .SI(N3454), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3571), .Q(N3455), .QN() );
  SDFFARX1 uWord_reg_6_ ( .D(n2535), .SI(N3455), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3571), .Q(N3456), .QN() );
  SDFFARX1 uWord_reg_7_ ( .D(n2534), .SI(N3456), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3571), .Q(N3457), .QN() );
  SDFFARX1 uWord_reg_8_ ( .D(n2533), .SI(N3457), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3570), .Q(N3458), .QN() );
  SDFFARX1 uWord_reg_9_ ( .D(n2532), .SI(N3458), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3570), .Q(N3459), .QN() );
  SDFFARX1 uWord_reg_10_ ( .D(n2531), .SI(N3459), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3570), .Q(N3460), .QN() );
  SDFFARX1 uWord_reg_11_ ( .D(n2530), .SI(N3460), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3570), .Q(N3461), .QN() );
  SDFFARX1 uWord_reg_12_ ( .D(n2529), .SI(N3461), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3570), .Q(N3462), .QN() );
  SDFFARX1 uWord_reg_13_ ( .D(n2528), .SI(N3462), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3570), .Q(N3463), .QN() );
  SDFFARX1 uWord_reg_14_ ( .D(n2527), .SI(N3463), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3569), .Q(test_so20), .QN() );
  SDFFARX1 CodeFetch_reg ( .D(n2591), .SI(n5209), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3603), .Q(n4821), .QN() );
  SDFFARX1 MemoryFetch_reg ( .D(n2593), .SI(M_IO_n), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3602), .Q(n4820), .QN() );
  SDFFARX1 lWord_reg_15_ ( .D(n2589), .SI(N3448), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3580), .Q(N3449), .QN() );
  SDFFARX1 lWord_reg_0_ ( .D(n2572), .SI(W_R_n), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3579), .Q(N3434), .QN() );
  SDFFARX1 lWord_reg_1_ ( .D(n2571), .SI(N3434), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3579), .Q(N3435), .QN() );
  SDFFARX1 lWord_reg_2_ ( .D(n2570), .SI(N3435), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3579), .Q(test_so17), .QN() );
  SDFFARX1 lWord_reg_3_ ( .D(n2569), .SI(test_si18), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3578), .Q(N3437), .QN() );
  SDFFARX1 lWord_reg_4_ ( .D(n2568), .SI(N3437), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3578), .Q(N3438), .QN() );
  SDFFARX1 lWord_reg_5_ ( .D(n2567), .SI(N3438), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3578), .Q(N3439), .QN() );
  SDFFARX1 lWord_reg_6_ ( .D(n2566), .SI(N3439), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3577), .Q(N3440), .QN() );
  SDFFARX1 lWord_reg_7_ ( .D(n2565), .SI(N3440), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3577), .Q(N3441), .QN() );
  SDFFARX1 lWord_reg_8_ ( .D(n2564), .SI(N3441), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3577), .Q(N3442), .QN() );
  SDFFARX1 lWord_reg_9_ ( .D(n2563), .SI(N3442), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3576), .Q(N3443), .QN() );
  SDFFARX1 lWord_reg_10_ ( .D(n2562), .SI(N3443), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3576), .Q(N3444), .QN() );
  SDFFARX1 lWord_reg_11_ ( .D(n2561), .SI(N3444), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3576), .Q(N3445), .QN() );
  SDFFARX1 lWord_reg_12_ ( .D(n2560), .SI(N3445), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3575), .Q(N3446), .QN() );
  SDFFARX1 lWord_reg_13_ ( .D(n2559), .SI(N3446), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3575), .Q(N3447), .QN() );
  SDFFARX1 lWord_reg_14_ ( .D(n2558), .SI(N3447), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3575), .Q(N3448), .QN() );
  SDFFARX1 ByteEnable_reg_2_ ( .D(n2430), .SI(n5216), .SE(test_se), .CLK(CLOCK), .RSTB(n3542), .Q(n5213), .QN() );
  SDFFARX1 ByteEnable_reg_1_ ( .D(n2428), .SI(n5218), .SE(test_se), .CLK(CLOCK), .RSTB(n3542), .Q(n5216), .QN() );
  SDFFARX1 ByteEnable_reg_3_ ( .D(n2432), .SI(n5213), .SE(test_se), .CLK(CLOCK), .RSTB(n3543), .Q(n5209), .QN(n3693) );
  SDFFARX1 ReadRequest_reg ( .D(n2595), .SI(PhyAddrPointer_31_), .SE(test_se), 
        .CLK(CLOCK), .RSTB(n3602), .Q(n4816), .QN(n1595) );
  SDFFARX1 ByteEnable_reg_0_ ( .D(n2426), .SI(BE_n[3]), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3542), .Q(n5218), .QN(n3692) );
  SDFFARX1 DataWidth_reg_0_ ( .D(n2835), .SI(D_C_n), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3610), .Q(test_so2), .QN(n1416) );
  SDFFARX1 DataWidth_reg_1_ ( .D(n2834), .SI(test_si3), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3610), .Q(n2864), .QN(n1415) );
  SDFFARX1 RequestPending_reg ( .D(n2841), .SI(n4816), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3611), .Q(n2889), .QN(n1596) );
  SDFFARX1 D_C_n_reg ( .D(n2590), .SI(n4821), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3602), .Q(D_C_n), .QN(n3872) );
  SDFFARX1 ADS_n_reg ( .D(n2837), .SI(test_si1), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3610), .Q(ADS_n), .QN() );
  SDFFARX1 rEIP_reg_30_ ( .D(n2626), .SI(rEIP_29_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3600), .Q(rEIP_30_), .QN(n2901) );
  SDFFARX1 M_IO_n_reg ( .D(n2592), .SI(n2915), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3602), .Q(M_IO_n), .QN() );
  SDFFARX1 W_R_n_reg ( .D(n2594), .SI(n2867), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3602), .Q(W_R_n), .QN() );
  SDFFARX1 BE_n_reg_3_ ( .D(n2431), .SI(BE_n[2]), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3543), .Q(BE_n[3]), .QN() );
  SDFFARX1 BE_n_reg_2_ ( .D(n2429), .SI(BE_n[1]), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3542), .Q(BE_n[2]), .QN() );
  SDFFARX1 BE_n_reg_1_ ( .D(n2427), .SI(BE_n[0]), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3542), .Q(BE_n[1]), .QN() );
  SDFFARX1 BE_n_reg_0_ ( .D(n2425), .SI(Address[29]), .SE(test_se), .CLK(CLOCK), .RSTB(n3542), .Q(BE_n[0]), .QN() );
  SDFFARX1 Datao_reg_0_ ( .D(n2463), .SI(n2864), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3569), .Q(Datao[0]), .QN() );
  SDFFARX1 Datao_reg_1_ ( .D(n2462), .SI(Datao[0]), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3569), .Q(Datao[1]), .QN() );
  SDFFARX1 Datao_reg_2_ ( .D(n2461), .SI(Datao[1]), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3569), .Q(Datao[2]), .QN() );
  SDFFARX1 Datao_reg_3_ ( .D(n2460), .SI(Datao[2]), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3569), .Q(Datao[3]), .QN() );
  SDFFARX1 Datao_reg_4_ ( .D(n2459), .SI(Datao[3]), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3569), .Q(Datao[4]), .QN() );
  SDFFARX1 Datao_reg_5_ ( .D(n2458), .SI(Datao[4]), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3568), .Q(Datao[5]), .QN() );
  SDFFARX1 Datao_reg_6_ ( .D(n2457), .SI(Datao[5]), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3568), .Q(Datao[6]), .QN() );
  SDFFARX1 Datao_reg_7_ ( .D(n2456), .SI(Datao[6]), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3568), .Q(Datao[7]), .QN() );
  SDFFARX1 Datao_reg_8_ ( .D(n2455), .SI(Datao[7]), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3568), .Q(Datao[8]), .QN() );
  SDFFARX1 Datao_reg_9_ ( .D(n2454), .SI(Datao[8]), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3568), .Q(Datao[9]), .QN() );
  SDFFARX1 Datao_reg_10_ ( .D(n2453), .SI(Datao[9]), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3568), .Q(Datao[10]), .QN() );
  SDFFARX1 Datao_reg_11_ ( .D(n2452), .SI(Datao[10]), .SE(test_se), .CLK(CLOCK), .RSTB(n3567), .Q(Datao[11]), .QN() );
  SDFFARX1 Datao_reg_12_ ( .D(n2451), .SI(Datao[11]), .SE(test_se), .CLK(CLOCK), .RSTB(n3567), .Q(Datao[12]), .QN() );
  SDFFARX1 Datao_reg_13_ ( .D(n2450), .SI(Datao[12]), .SE(test_se), .CLK(CLOCK), .RSTB(n3567), .Q(Datao[13]), .QN() );
  SDFFARX1 Datao_reg_14_ ( .D(n2449), .SI(Datao[13]), .SE(test_se), .CLK(CLOCK), .RSTB(n3567), .Q(Datao[14]), .QN() );
  SDFFARX1 Datao_reg_15_ ( .D(n2448), .SI(Datao[14]), .SE(test_se), .CLK(CLOCK), .RSTB(n3567), .Q(Datao[15]), .QN() );
  SDFFARX1 Datao_reg_16_ ( .D(n2447), .SI(Datao[15]), .SE(test_se), .CLK(CLOCK), .RSTB(n3567), .Q(Datao[16]), .QN() );
  SDFFARX1 Datao_reg_17_ ( .D(n2446), .SI(Datao[16]), .SE(test_se), .CLK(CLOCK), .RSTB(n3566), .Q(Datao[17]), .QN() );
  SDFFARX1 Datao_reg_18_ ( .D(n2445), .SI(Datao[17]), .SE(test_se), .CLK(CLOCK), .RSTB(n3566), .Q(Datao[18]), .QN() );
  SDFFARX1 Datao_reg_19_ ( .D(n2444), .SI(Datao[18]), .SE(test_se), .CLK(CLOCK), .RSTB(n3566), .Q(Datao[19]), .QN() );
  SDFFARX1 Datao_reg_20_ ( .D(n2443), .SI(test_si4), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3566), .Q(Datao[20]), .QN() );
  SDFFARX1 Datao_reg_21_ ( .D(n2442), .SI(Datao[20]), .SE(test_se), .CLK(CLOCK), .RSTB(n3566), .Q(Datao[21]), .QN() );
  SDFFARX1 Datao_reg_22_ ( .D(n2441), .SI(Datao[21]), .SE(test_se), .CLK(CLOCK), .RSTB(n3566), .Q(Datao[22]), .QN() );
  SDFFARX1 Datao_reg_23_ ( .D(n2440), .SI(Datao[22]), .SE(test_se), .CLK(CLOCK), .RSTB(n3565), .Q(Datao[23]), .QN() );
  SDFFARX1 Datao_reg_24_ ( .D(n2439), .SI(Datao[23]), .SE(test_se), .CLK(CLOCK), .RSTB(n3565), .Q(Datao[24]), .QN() );
  SDFFARX1 Datao_reg_25_ ( .D(n2438), .SI(Datao[24]), .SE(test_se), .CLK(CLOCK), .RSTB(n3565), .Q(Datao[25]), .QN() );
  SDFFARX1 Datao_reg_26_ ( .D(n2437), .SI(Datao[25]), .SE(test_se), .CLK(CLOCK), .RSTB(n3565), .Q(Datao[26]), .QN() );
  SDFFARX1 Datao_reg_27_ ( .D(n2436), .SI(Datao[26]), .SE(test_se), .CLK(CLOCK), .RSTB(n3565), .Q(Datao[27]), .QN() );
  SDFFARX1 Datao_reg_28_ ( .D(n2435), .SI(Datao[27]), .SE(test_se), .CLK(CLOCK), .RSTB(n3565), .Q(Datao[28]), .QN() );
  SDFFARX1 Datao_reg_29_ ( .D(n2434), .SI(Datao[28]), .SE(test_se), .CLK(CLOCK), .RSTB(n3564), .Q(Datao[29]), .QN() );
  SDFFARX1 Datao_reg_30_ ( .D(n2433), .SI(Datao[29]), .SE(test_se), .CLK(CLOCK), .RSTB(n3564), .Q(Datao[30]), .QN() );
  SDFFARX1 Address_reg_0_ ( .D(n2625), .SI(ADS_n), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3585), .Q(Address[0]), .QN() );
  SDFFARX1 Address_reg_1_ ( .D(n2624), .SI(Address[0]), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3585), .Q(Address[1]), .QN() );
  SDFFARX1 Address_reg_2_ ( .D(n2623), .SI(Address[1]), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3585), .Q(Address[2]), .QN() );
  SDFFARX1 Address_reg_3_ ( .D(n2622), .SI(Address[2]), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3585), .Q(Address[3]), .QN() );
  SDFFARX1 Address_reg_4_ ( .D(n2621), .SI(Address[3]), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3585), .Q(Address[4]), .QN() );
  SDFFARX1 Address_reg_5_ ( .D(n2620), .SI(Address[4]), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3584), .Q(Address[5]), .QN() );
  SDFFARX1 Address_reg_6_ ( .D(n2619), .SI(Address[5]), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3584), .Q(Address[6]), .QN() );
  SDFFARX1 Address_reg_7_ ( .D(n2618), .SI(Address[6]), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3584), .Q(Address[7]), .QN() );
  SDFFARX1 Address_reg_8_ ( .D(n2617), .SI(Address[7]), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3584), .Q(Address[8]), .QN() );
  SDFFARX1 Address_reg_9_ ( .D(n2616), .SI(Address[8]), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3584), .Q(Address[9]), .QN() );
  SDFFARX1 Address_reg_10_ ( .D(n2615), .SI(Address[9]), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3584), .Q(Address[10]), .QN() );
  SDFFARX1 Address_reg_11_ ( .D(n2614), .SI(Address[10]), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3583), .Q(Address[11]), .QN() );
  SDFFARX1 Address_reg_12_ ( .D(n2613), .SI(Address[11]), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3583), .Q(Address[12]), .QN() );
  SDFFARX1 Address_reg_13_ ( .D(n2612), .SI(Address[12]), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3583), .Q(Address[13]), .QN() );
  SDFFARX1 Address_reg_14_ ( .D(n2611), .SI(Address[13]), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3583), .Q(Address[14]), .QN() );
  SDFFARX1 Address_reg_15_ ( .D(n2610), .SI(Address[14]), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3583), .Q(Address[15]), .QN() );
  SDFFARX1 Address_reg_16_ ( .D(n2609), .SI(Address[15]), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3583), .Q(Address[16]), .QN() );
  SDFFARX1 Address_reg_17_ ( .D(n2608), .SI(Address[16]), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3582), .Q(Address[17]), .QN() );
  SDFFARX1 Address_reg_18_ ( .D(n2607), .SI(Address[17]), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3582), .Q(Address[18]), .QN() );
  SDFFARX1 Address_reg_19_ ( .D(n2606), .SI(Address[18]), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3582), .Q(Address[19]), .QN() );
  SDFFARX1 Address_reg_20_ ( .D(n2605), .SI(test_si2), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3582), .Q(Address[20]), .QN() );
  SDFFARX1 Address_reg_21_ ( .D(n2604), .SI(Address[20]), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3582), .Q(Address[21]), .QN() );
  SDFFARX1 Address_reg_22_ ( .D(n2603), .SI(Address[21]), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3582), .Q(Address[22]), .QN() );
  SDFFARX1 Address_reg_23_ ( .D(n2602), .SI(Address[22]), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3581), .Q(Address[23]), .QN() );
  SDFFARX1 Address_reg_24_ ( .D(n2601), .SI(Address[23]), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3581), .Q(Address[24]), .QN() );
  SDFFARX1 Address_reg_25_ ( .D(n2600), .SI(Address[24]), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3581), .Q(Address[25]), .QN() );
  SDFFARX1 Address_reg_26_ ( .D(n2599), .SI(Address[25]), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3581), .Q(Address[26]), .QN() );
  SDFFARX1 Address_reg_27_ ( .D(n2598), .SI(Address[26]), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3581), .Q(Address[27]), .QN() );
  SDFFARX1 Address_reg_28_ ( .D(n2597), .SI(Address[27]), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3581), .Q(Address[28]), .QN() );
  SDFFARX1 Address_reg_29_ ( .D(n2596), .SI(Address[28]), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3580), .Q(Address[29]), .QN() );
  SDFFARX1 PhyAddrPointer_reg_31_ ( .D(n2464), .SI(PhyAddrPointer_30_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3601), .Q(PhyAddrPointer_31_), .QN(n1558) );
  SDFFARX1 EAX_reg_30_ ( .D(n2543), .SI(EAX_29_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3580), .Q(test_so5), .QN() );
  SDFFARX1 More_reg ( .D(n2657), .SI(n4820), .SE(test_se), .CLK(CLOCK), .RSTB(
        n3608), .Q(n5326), .QN(n3873) );
  SDFFARX1 EAX_reg_23_ ( .D(n2550), .SI(EAX_22_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3573), .Q(EAX_23_), .QN() );
  SDFFARX1 EAX_reg_24_ ( .D(n2549), .SI(EAX_23_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3573), .Q(EAX_24_), .QN() );
  SDFFARX1 EAX_reg_25_ ( .D(n2548), .SI(EAX_24_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3573), .Q(EAX_25_), .QN() );
  SDFFARX1 EAX_reg_26_ ( .D(n2547), .SI(EAX_25_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3573), .Q(EAX_26_), .QN() );
  SDFFARX1 EAX_reg_27_ ( .D(n2546), .SI(EAX_26_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3572), .Q(EAX_27_), .QN() );
  SDFFARX1 EAX_reg_28_ ( .D(n2545), .SI(EAX_27_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3572), .Q(EAX_28_), .QN() );
  SDFFARX1 EAX_reg_29_ ( .D(n2544), .SI(EAX_28_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3572), .Q(EAX_29_), .QN() );
  SDFFARX1 Flush_reg ( .D(n2794), .SI(N1954), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3608), .Q(n2870), .QN(n1590) );
  SDFFARX1 PhyAddrPointer_reg_30_ ( .D(n2465), .SI(PhyAddrPointer_29_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3600), .Q(PhyAddrPointer_30_), .QN(n1559) );
  SDFFARX1 PhyAddrPointer_reg_29_ ( .D(n2466), .SI(PhyAddrPointer_28_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3600), .Q(PhyAddrPointer_29_), .QN(n1560) );
  SDFFARX1 PhyAddrPointer_reg_24_ ( .D(n2471), .SI(PhyAddrPointer_23_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3592), .Q(test_so16), .QN(n1565) );
  SDFFARX1 PhyAddrPointer_reg_25_ ( .D(n2470), .SI(test_si17), .SE(test_se), 
        .CLK(CLOCK), .RSTB(n3592), .Q(PhyAddrPointer_25_), .QN(n1564) );
  SDFFARX1 PhyAddrPointer_reg_26_ ( .D(n2469), .SI(PhyAddrPointer_25_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3591), .Q(PhyAddrPointer_26_), .QN(n1563) );
  SDFFARX1 PhyAddrPointer_reg_27_ ( .D(n2468), .SI(PhyAddrPointer_26_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3591), .Q(PhyAddrPointer_27_), .QN(n1562) );
  SDFFARX1 PhyAddrPointer_reg_28_ ( .D(n2467), .SI(PhyAddrPointer_27_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3591), .Q(PhyAddrPointer_28_), .QN(n1561) );
  SDFFARX1 InstAddrPointer_reg_31_ ( .D(n2832), .SI(InstAddrPointer_30_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3601), .Q(N3467), .QN(n3869) );
  SDFFARX1 EBX_reg_23_ ( .D(n2802), .SI(EBX_22_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3604), .Q(EBX_23_), .QN() );
  SDFFARX1 EBX_reg_24_ ( .D(n2801), .SI(EBX_23_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3604), .Q(EBX_24_), .QN() );
  SDFFARX1 EBX_reg_25_ ( .D(n2800), .SI(EBX_24_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3604), .Q(EBX_25_), .QN() );
  SDFFARX1 EBX_reg_26_ ( .D(n2799), .SI(EBX_25_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3604), .Q(EBX_26_), .QN() );
  SDFFARX1 EBX_reg_27_ ( .D(n2798), .SI(EBX_26_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3603), .Q(EBX_27_), .QN() );
  SDFFARX1 EBX_reg_28_ ( .D(n2797), .SI(EBX_27_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3603), .Q(EBX_28_), .QN() );
  SDFFARX1 EBX_reg_29_ ( .D(n2796), .SI(EBX_28_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3603), .Q(EBX_29_), .QN() );
  SDFFARX1 EBX_reg_30_ ( .D(n2795), .SI(EBX_29_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3603), .Q(EBX_30_), .QN() );
  SDFFARX1 InstAddrPointer_reg_30_ ( .D(n2496), .SI(InstAddrPointer_29_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3590), .Q(InstAddrPointer_30_), .QN(
        n3868) );
  SDFFARX1 InstAddrPointer_reg_23_ ( .D(n2503), .SI(InstAddrPointer_22_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3586), .Q(InstAddrPointer_23_), .QN(
        n3846) );
  SDFFARX1 InstAddrPointer_reg_24_ ( .D(n2502), .SI(InstAddrPointer_23_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3586), .Q(InstAddrPointer_24_), .QN(
        n3845) );
  SDFFARX1 InstAddrPointer_reg_25_ ( .D(n2501), .SI(InstAddrPointer_24_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3586), .Q(InstAddrPointer_25_), .QN(
        n3844) );
  SDFFARX1 InstAddrPointer_reg_26_ ( .D(n2500), .SI(InstAddrPointer_25_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3586), .Q(InstAddrPointer_26_), .QN(
        n3843) );
  SDFFARX1 InstAddrPointer_reg_27_ ( .D(n2499), .SI(InstAddrPointer_26_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3586), .Q(InstAddrPointer_27_), .QN(
        n3842) );
  SDFFARX1 InstAddrPointer_reg_28_ ( .D(n2498), .SI(InstAddrPointer_27_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3586), .Q(test_so8), .QN(n3841) );
  SDFFARX1 InstAddrPointer_reg_29_ ( .D(n2497), .SI(test_si9), .SE(test_se), 
        .CLK(CLOCK), .RSTB(n3585), .Q(InstAddrPointer_29_), .QN(n3840) );
  SDFFARX1 EBX_reg_31_ ( .D(n2826), .SI(EBX_30_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3608), .Q(N1954), .QN() );
  SDFFARX1 rEIP_reg_14_ ( .D(n2642), .SI(rEIP_13_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3595), .Q(rEIP_14_), .QN(n4744) );
  SDFFARX1 rEIP_reg_15_ ( .D(n2641), .SI(rEIP_14_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3595), .Q(rEIP_15_), .QN(n4749) );
  SDFFARX1 rEIP_reg_16_ ( .D(n2640), .SI(rEIP_15_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3595), .Q(rEIP_16_), .QN(n4754) );
  SDFFARX1 rEIP_reg_17_ ( .D(n2639), .SI(rEIP_16_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3594), .Q(rEIP_17_), .QN(n4759) );
  SDFFARX1 rEIP_reg_18_ ( .D(n2638), .SI(rEIP_17_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3594), .Q(rEIP_18_), .QN(n4764) );
  SDFFARX1 rEIP_reg_19_ ( .D(n2637), .SI(rEIP_18_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3594), .Q(rEIP_19_), .QN(n4769) );
  SDFFARX1 rEIP_reg_20_ ( .D(n2636), .SI(rEIP_19_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3593), .Q(rEIP_20_), .QN(n2891) );
  SDFFARX1 rEIP_reg_21_ ( .D(n2635), .SI(rEIP_20_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3593), .Q(rEIP_21_), .QN(n2892) );
  SDFFARX1 rEIP_reg_22_ ( .D(n2634), .SI(rEIP_21_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3593), .Q(rEIP_22_), .QN(n2893) );
  SDFFARX1 rEIP_reg_23_ ( .D(n2633), .SI(rEIP_22_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3592), .Q(rEIP_23_), .QN(n2894) );
  SDFFARX1 rEIP_reg_24_ ( .D(n2632), .SI(rEIP_23_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3592), .Q(rEIP_24_), .QN(n2895) );
  SDFFARX1 rEIP_reg_25_ ( .D(n2631), .SI(rEIP_24_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3592), .Q(rEIP_25_), .QN(n2896) );
  SDFFARX1 rEIP_reg_26_ ( .D(n2630), .SI(rEIP_25_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3591), .Q(test_so19), .QN(n2897) );
  SDFFARX1 rEIP_reg_27_ ( .D(n2629), .SI(test_si20), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3591), .Q(rEIP_27_), .QN(n2898) );
  SDFFARX1 rEIP_reg_28_ ( .D(n2628), .SI(rEIP_27_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3591), .Q(rEIP_28_), .QN(n2899) );
  SDFFARX1 rEIP_reg_29_ ( .D(n2627), .SI(rEIP_28_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3590), .Q(rEIP_29_), .QN(n2900) );
  SDFFARX1 EAX_reg_15_ ( .D(n2573), .SI(N3360), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3574), .Q(N3361), .QN(n3823) );
  SDFFARX1 State2_reg_3_ ( .D(n2828), .SI(n2865), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3609), .Q(n4097), .QN() );
  SDFFARX1 EAX_reg_31_ ( .D(n2542), .SI(test_si6), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3572), .Q(EAX_31_), .QN(n3822) );
  SDFFARX1 EAX_reg_16_ ( .D(n2557), .SI(N3361), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3574), .Q(EAX_16_), .QN() );
  SDFFARX1 EAX_reg_17_ ( .D(n2556), .SI(EAX_16_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3574), .Q(EAX_17_), .QN() );
  SDFFARX1 EAX_reg_18_ ( .D(n2555), .SI(EAX_17_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3574), .Q(EAX_18_), .QN() );
  SDFFARX1 EAX_reg_19_ ( .D(n2554), .SI(EAX_18_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3574), .Q(EAX_19_), .QN() );
  SDFFARX1 EAX_reg_20_ ( .D(n2553), .SI(EAX_19_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3574), .Q(EAX_20_), .QN() );
  SDFFARX1 EAX_reg_21_ ( .D(n2552), .SI(EAX_20_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3573), .Q(EAX_21_), .QN() );
  SDFFARX1 EAX_reg_22_ ( .D(n2551), .SI(EAX_21_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3573), .Q(EAX_22_), .QN() );
  SDFFARX1 State2_reg_1_ ( .D(n2827), .SI(n2842), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3603), .Q(n2844), .QN(n1491) );
  SDFFARX1 State2_reg_0_ ( .D(n2830), .SI(n2889), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3610), .Q(n2842), .QN(n1492) );
  SDFFARX1 State2_reg_2_ ( .D(n2829), .SI(n2844), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3609), .Q(n2865), .QN(n1490) );
  SDFFARX1 State_reg_1_ ( .D(n2839), .SI(n4045), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3611), .Q(n2847), .QN(n1435) );
  SDFFARX1 StateBS16_reg ( .D(n2836), .SI(n4097), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3610), .Q(n2868), .QN(n1472) );
  SDFFARX1 State_reg_2_ ( .D(n2840), .SI(n2847), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3611), .Q(n2867), .QN(n1434) );
  SDFFARX1 State_reg_0_ ( .D(n2838), .SI(n2868), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3610), .Q(n4045), .QN(n1436) );
  SDFFARX1 PhyAddrPointer_reg_8_ ( .D(n2487), .SI(PhyAddrPointer_7_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3597), .Q(PhyAddrPointer_8_), .QN(n1581)
         );
  SDFFARX1 PhyAddrPointer_reg_9_ ( .D(n2486), .SI(PhyAddrPointer_8_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3597), .Q(PhyAddrPointer_9_), .QN(n1580)
         );
  SDFFARX1 PhyAddrPointer_reg_10_ ( .D(n2485), .SI(PhyAddrPointer_9_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3597), .Q(PhyAddrPointer_10_), .QN(n1579) );
  SDFFARX1 PhyAddrPointer_reg_11_ ( .D(n2484), .SI(PhyAddrPointer_10_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3596), .Q(PhyAddrPointer_11_), .QN(n1578) );
  SDFFARX1 PhyAddrPointer_reg_12_ ( .D(n2483), .SI(PhyAddrPointer_11_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3596), .Q(PhyAddrPointer_12_), .QN(n1577) );
  SDFFARX1 PhyAddrPointer_reg_13_ ( .D(n2482), .SI(PhyAddrPointer_12_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3596), .Q(PhyAddrPointer_13_), .QN(n1576) );
  SDFFARX1 PhyAddrPointer_reg_14_ ( .D(n2481), .SI(PhyAddrPointer_13_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3595), .Q(PhyAddrPointer_14_), .QN(n1575) );
  SDFFARX1 PhyAddrPointer_reg_15_ ( .D(n2480), .SI(PhyAddrPointer_14_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3595), .Q(PhyAddrPointer_15_), .QN(n1574) );
  SDFFARX1 PhyAddrPointer_reg_16_ ( .D(n2479), .SI(PhyAddrPointer_15_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3595), .Q(PhyAddrPointer_16_), .QN(n1573) );
  SDFFARX1 PhyAddrPointer_reg_17_ ( .D(n2478), .SI(PhyAddrPointer_16_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3594), .Q(PhyAddrPointer_17_), .QN(n1572) );
  SDFFARX1 PhyAddrPointer_reg_18_ ( .D(n2477), .SI(PhyAddrPointer_17_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3594), .Q(PhyAddrPointer_18_), .QN(n1571) );
  SDFFARX1 PhyAddrPointer_reg_19_ ( .D(n2476), .SI(PhyAddrPointer_18_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3594), .Q(PhyAddrPointer_19_), .QN(n1570) );
  SDFFARX1 PhyAddrPointer_reg_20_ ( .D(n2475), .SI(PhyAddrPointer_19_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3593), .Q(PhyAddrPointer_20_), .QN(n1569) );
  SDFFARX1 PhyAddrPointer_reg_21_ ( .D(n2474), .SI(PhyAddrPointer_20_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3593), .Q(PhyAddrPointer_21_), .QN(n1568) );
  SDFFARX1 PhyAddrPointer_reg_22_ ( .D(n2473), .SI(PhyAddrPointer_21_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3593), .Q(PhyAddrPointer_22_), .QN(n1567) );
  SDFFARX1 PhyAddrPointer_reg_23_ ( .D(n2472), .SI(PhyAddrPointer_22_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3592), .Q(PhyAddrPointer_23_), .QN(n1566) );
  SDFFARX1 EBX_reg_15_ ( .D(n2810), .SI(EBX_14_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3605), .Q(EBX_15_), .QN() );
  SDFFARX1 EBX_reg_16_ ( .D(n2809), .SI(EBX_15_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3605), .Q(EBX_16_), .QN() );
  SDFFARX1 EBX_reg_17_ ( .D(n2808), .SI(EBX_16_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3605), .Q(EBX_17_), .QN() );
  SDFFARX1 EBX_reg_18_ ( .D(n2807), .SI(EBX_17_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3605), .Q(EBX_18_), .QN() );
  SDFFARX1 EBX_reg_19_ ( .D(n2806), .SI(EBX_18_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3605), .Q(test_so6), .QN() );
  SDFFARX1 EBX_reg_20_ ( .D(n2805), .SI(test_si7), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3605), .Q(EBX_20_), .QN() );
  SDFFARX1 EBX_reg_21_ ( .D(n2804), .SI(EBX_20_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3604), .Q(EBX_21_), .QN() );
  SDFFARX1 EBX_reg_22_ ( .D(n2803), .SI(EBX_21_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3604), .Q(EBX_22_), .QN() );
  SDFFARX1 InstAddrPointer_reg_16_ ( .D(n2510), .SI(InstAddrPointer_15_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3588), .Q(InstAddrPointer_16_), .QN(
        n3853) );
  SDFFARX1 InstAddrPointer_reg_17_ ( .D(n2509), .SI(InstAddrPointer_16_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3587), .Q(InstAddrPointer_17_), .QN(
        n3852) );
  SDFFARX1 InstAddrPointer_reg_18_ ( .D(n2508), .SI(InstAddrPointer_17_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3587), .Q(InstAddrPointer_18_), .QN(
        n3851) );
  SDFFARX1 InstAddrPointer_reg_19_ ( .D(n2507), .SI(InstAddrPointer_18_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3587), .Q(InstAddrPointer_19_), .QN(
        n3850) );
  SDFFARX1 InstAddrPointer_reg_20_ ( .D(n2506), .SI(InstAddrPointer_19_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3587), .Q(InstAddrPointer_20_), .QN(
        n3849) );
  SDFFARX1 InstAddrPointer_reg_21_ ( .D(n2505), .SI(InstAddrPointer_20_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3587), .Q(InstAddrPointer_21_), .QN(
        n3848) );
  SDFFARX1 InstAddrPointer_reg_22_ ( .D(n2504), .SI(InstAddrPointer_21_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3587), .Q(InstAddrPointer_22_), .QN(
        n3847) );
  SDFFARX1 InstQueueWr_Addr_reg_2_ ( .D(n2787), .SI(N3991), .SE(test_se), 
        .CLK(CLOCK), .RSTB(n3609), .Q(N3990), .QN(n1554) );
  SDFFARX1 InstQueueWr_Addr_reg_3_ ( .D(n2786), .SI(N3990), .SE(test_se), 
        .CLK(CLOCK), .RSTB(n3609), .Q(N3989), .QN(n1553) );
  SDFFARX1 PhyAddrPointer_reg_0_ ( .D(n2495), .SI(n5326), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3600), .Q(PhyAddrPointer_0_), .QN(n1589) );
  SDFFARX1 rEIP_reg_5_ ( .D(n2651), .SI(rEIP_4_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3601), .Q(rEIP_5_), .QN(n4700) );
  SDFFARX1 rEIP_reg_2_ ( .D(n2654), .SI(rEIP_1_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3599), .Q(rEIP_2_), .QN(n4680) );
  SDFFARX1 rEIP_reg_3_ ( .D(n2653), .SI(rEIP_2_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3599), .Q(rEIP_3_), .QN(n4686) );
  SDFFARX1 rEIP_reg_4_ ( .D(n2652), .SI(rEIP_3_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3598), .Q(rEIP_4_), .QN(n4692) );
  SDFFARX1 rEIP_reg_6_ ( .D(n2650), .SI(rEIP_5_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3598), .Q(test_so18), .QN(n4704) );
  SDFFARX1 rEIP_reg_7_ ( .D(n2649), .SI(test_si19), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3598), .Q(rEIP_7_), .QN(n4709) );
  SDFFARX1 rEIP_reg_8_ ( .D(n2648), .SI(rEIP_7_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3597), .Q(rEIP_8_), .QN(n4714) );
  SDFFARX1 rEIP_reg_9_ ( .D(n2647), .SI(rEIP_8_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3597), .Q(rEIP_9_), .QN(n4719) );
  SDFFARX1 rEIP_reg_10_ ( .D(n2646), .SI(rEIP_9_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3597), .Q(rEIP_10_), .QN(n4724) );
  SDFFARX1 rEIP_reg_11_ ( .D(n2645), .SI(rEIP_10_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3596), .Q(rEIP_11_), .QN(n4729) );
  SDFFARX1 rEIP_reg_12_ ( .D(n2644), .SI(rEIP_11_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3596), .Q(rEIP_12_), .QN(n4734) );
  SDFFARX1 rEIP_reg_13_ ( .D(n2643), .SI(rEIP_12_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3596), .Q(rEIP_13_), .QN(n4739) );
  SDFFARX1 InstQueueRd_Addr_reg_4_ ( .D(n2790), .SI(InstQueueRd_Addr[3]), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3601), .Q(InstQueueRd_Addr[4]), .QN(
        n3871) );
  SDFFARX1 rEIP_reg_1_ ( .D(n2655), .SI(rEIP_0_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3599), .Q(rEIP_1_), .QN(n2888) );
  SDFFARX1 EAX_reg_7_ ( .D(n2581), .SI(N3352), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3577), .Q(N3353), .QN(n3831) );
  SDFFARX1 EAX_reg_8_ ( .D(n2580), .SI(N3353), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3577), .Q(N3354), .QN(n3830) );
  SDFFARX1 EAX_reg_9_ ( .D(n2579), .SI(N3354), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3576), .Q(test_so4), .QN(n3829) );
  SDFFARX1 EAX_reg_10_ ( .D(n2578), .SI(test_si5), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3576), .Q(N3356), .QN(n3828) );
  SDFFARX1 EAX_reg_11_ ( .D(n2577), .SI(N3356), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3576), .Q(N3357), .QN(n3827) );
  SDFFARX1 EAX_reg_12_ ( .D(n2576), .SI(N3357), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3575), .Q(N3358), .QN(n3826) );
  SDFFARX1 EAX_reg_13_ ( .D(n2575), .SI(N3358), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3575), .Q(N3359), .QN(n3825) );
  SDFFARX1 EAX_reg_14_ ( .D(n2574), .SI(N3359), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3575), .Q(N3360), .QN(n3824) );
  SDFFARX1 InstQueueWr_Addr_reg_0_ ( .D(n2789), .SI(InstQueueRd_Addr[4]), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3609), .Q(N1239), .QN(n1556) );
  SDFFARX1 InstQueueWr_Addr_reg_1_ ( .D(n2788), .SI(N1239), .SE(test_se), 
        .CLK(CLOCK), .RSTB(n3609), .Q(N3991), .QN(n1555) );
  SDFFARX1 rEIP_reg_0_ ( .D(n2656), .SI(N3449), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3600), .Q(rEIP_0_), .QN(n2845) );
  SDFFARX1 PhyAddrPointer_reg_5_ ( .D(n2490), .SI(PhyAddrPointer_4_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3600), .Q(PhyAddrPointer_5_), .QN(n1584)
         );
  SDFFARX1 PhyAddrPointer_reg_3_ ( .D(n2492), .SI(PhyAddrPointer_2_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3599), .Q(test_so15), .QN(n1586) );
  SDFFARX1 PhyAddrPointer_reg_4_ ( .D(n2491), .SI(test_si16), .SE(test_se), 
        .CLK(CLOCK), .RSTB(n3598), .Q(PhyAddrPointer_4_), .QN(n1585) );
  SDFFARX1 PhyAddrPointer_reg_6_ ( .D(n2489), .SI(PhyAddrPointer_5_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3598), .Q(PhyAddrPointer_6_), .QN(n1583)
         );
  SDFFARX1 PhyAddrPointer_reg_7_ ( .D(n2488), .SI(PhyAddrPointer_6_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3598), .Q(PhyAddrPointer_7_), .QN(n1582)
         );
  SDFFARX1 rEIP_reg_31_ ( .D(n2833), .SI(rEIP_30_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3601), .Q(rEIP_31_), .QN(n2866) );
  SDFFARX1 EBX_reg_8_ ( .D(n2817), .SI(EBX_7_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3607), .Q(EBX_8_), .QN() );
  SDFFARX1 EBX_reg_9_ ( .D(n2816), .SI(EBX_8_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3606), .Q(EBX_9_), .QN() );
  SDFFARX1 EBX_reg_10_ ( .D(n2815), .SI(EBX_9_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3606), .Q(EBX_10_), .QN() );
  SDFFARX1 EBX_reg_11_ ( .D(n2814), .SI(EBX_10_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3606), .Q(EBX_11_), .QN() );
  SDFFARX1 EBX_reg_12_ ( .D(n2813), .SI(EBX_11_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3606), .Q(EBX_12_), .QN() );
  SDFFARX1 EBX_reg_13_ ( .D(n2812), .SI(EBX_12_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3606), .Q(EBX_13_), .QN() );
  SDFFARX1 EBX_reg_14_ ( .D(n2811), .SI(EBX_13_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3606), .Q(EBX_14_), .QN() );
  SDFFARX1 InstAddrPointer_reg_8_ ( .D(n2518), .SI(test_si8), .SE(test_se), 
        .CLK(CLOCK), .RSTB(n3589), .Q(InstAddrPointer_8_), .QN(n3861) );
  SDFFARX1 InstAddrPointer_reg_9_ ( .D(n2517), .SI(InstAddrPointer_8_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3589), .Q(InstAddrPointer_9_), .QN(n3860) );
  SDFFARX1 InstAddrPointer_reg_10_ ( .D(n2516), .SI(InstAddrPointer_9_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3589), .Q(InstAddrPointer_10_), .QN(
        n3859) );
  SDFFARX1 InstAddrPointer_reg_11_ ( .D(n2515), .SI(InstAddrPointer_10_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3588), .Q(InstAddrPointer_11_), .QN(
        n3858) );
  SDFFARX1 InstAddrPointer_reg_12_ ( .D(n2514), .SI(InstAddrPointer_11_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3588), .Q(InstAddrPointer_12_), .QN(
        n3857) );
  SDFFARX1 InstAddrPointer_reg_13_ ( .D(n2513), .SI(InstAddrPointer_12_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3588), .Q(InstAddrPointer_13_), .QN(
        n3856) );
  SDFFARX1 InstAddrPointer_reg_14_ ( .D(n2512), .SI(InstAddrPointer_13_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3588), .Q(InstAddrPointer_14_), .QN(
        n3855) );
  SDFFARX1 InstAddrPointer_reg_15_ ( .D(n2511), .SI(InstAddrPointer_14_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3588), .Q(InstAddrPointer_15_), .QN(
        n3854) );
  SDFFARX1 PhyAddrPointer_reg_1_ ( .D(n2494), .SI(PhyAddrPointer_0_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3599), .Q(PhyAddrPointer_1_), .QN(n1588)
         );
  SDFFARX1 PhyAddrPointer_reg_2_ ( .D(n2493), .SI(PhyAddrPointer_1_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3599), .Q(PhyAddrPointer_2_), .QN(n1587)
         );
  SDFFARX1 EAX_reg_1_ ( .D(n2587), .SI(N3346), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3579), .Q(N3347), .QN(n3837) );
  SDFFARX1 EAX_reg_2_ ( .D(n2586), .SI(N3347), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3579), .Q(N3348), .QN(n3836) );
  SDFFARX1 EAX_reg_3_ ( .D(n2585), .SI(N3348), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3578), .Q(N3349), .QN(n3835) );
  SDFFARX1 EAX_reg_4_ ( .D(n2584), .SI(N3349), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3578), .Q(N3350), .QN(n3834) );
  SDFFARX1 EAX_reg_5_ ( .D(n2583), .SI(N3350), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3578), .Q(N3351), .QN(n3833) );
  SDFFARX1 EAX_reg_6_ ( .D(n2582), .SI(N3351), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3577), .Q(N3352), .QN(n3832) );
  SDFFARX1 InstQueue_reg_14__7_ ( .D(n2666), .SI(n2874), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3563), .Q(n2875), .QN(n3813) );
  SDFFARX1 InstQueue_reg_14__6_ ( .D(n2667), .SI(n2873), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3563), .Q(n2874), .QN(n3812) );
  SDFFARX1 InstQueue_reg_14__5_ ( .D(n2668), .SI(n2872), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3562), .Q(n2873), .QN(n3811) );
  SDFFARX1 InstQueue_reg_14__4_ ( .D(n2669), .SI(n2871), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3562), .Q(n2872), .QN(n3810) );
  SDFFARX1 InstQueue_reg_1__7_ ( .D(n2770), .SI(n4250), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3545), .Q(n4253), .QN(n3709) );
  SDFFARX1 InstQueue_reg_1__6_ ( .D(n2771), .SI(n4247), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3545), .Q(n4250), .QN(n3708) );
  SDFFARX1 InstQueue_reg_1__5_ ( .D(n2772), .SI(n4244), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3545), .Q(n4247), .QN(n3707) );
  SDFFARX1 InstQueue_reg_0__7_ ( .D(n2778), .SI(N2554), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3544), .Q(N2555), .QN(n3701) );
  SDFFARX1 InstQueue_reg_0__6_ ( .D(n2779), .SI(N2553), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3544), .Q(N2554), .QN(n3700) );
  SDFFARX1 InstQueue_reg_0__5_ ( .D(n2780), .SI(N2552), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3544), .Q(N2553), .QN(n3699) );
  SDFFARX1 InstQueue_reg_0__4_ ( .D(n2781), .SI(N2551), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3544), .Q(N2552), .QN(n3698) );
  SDFFARX1 InstQueue_reg_5__7_ ( .D(n2738), .SI(n4365), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3551), .Q(n4368), .QN(n3741) );
  SDFFARX1 InstQueue_reg_5__6_ ( .D(n2739), .SI(n4362), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3551), .Q(n4365), .QN(n3740) );
  SDFFARX1 InstQueue_reg_5__5_ ( .D(n2740), .SI(n4359), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3550), .Q(n4362), .QN(n3739) );
  SDFFARX1 InstQueue_reg_5__4_ ( .D(n2741), .SI(n4355), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3550), .Q(n4359), .QN(n3738) );
  SDFFARX1 InstQueue_reg_4__7_ ( .D(n2746), .SI(n4333), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3549), .Q(n4336), .QN(n3733) );
  SDFFARX1 InstQueue_reg_4__6_ ( .D(n2747), .SI(n4330), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3549), .Q(n4333), .QN(n3732) );
  SDFFARX1 InstQueue_reg_4__5_ ( .D(n2748), .SI(n4326), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3549), .Q(n4330), .QN(n3731) );
  SDFFARX1 InstQueue_reg_4__4_ ( .D(n2749), .SI(n4323), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3549), .Q(n4326), .QN(n3730) );
  SDFFARX1 InstQueue_reg_2__7_ ( .D(n2762), .SI(n2859), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3547), .Q(n2860), .QN(n3717) );
  SDFFARX1 InstQueue_reg_2__6_ ( .D(n2763), .SI(n2858), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3547), .Q(n2859), .QN(n3716) );
  SDFFARX1 InstQueue_reg_2__5_ ( .D(n2764), .SI(n2857), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3546), .Q(n2858), .QN(n3715) );
  SDFFARX1 InstQueue_reg_2__4_ ( .D(n2765), .SI(n2863), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3546), .Q(n2857), .QN(n3714) );
  SDFFARX1 InstQueue_reg_12__7_ ( .D(n2682), .SI(n4557), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3560), .Q(n4560), .QN(n3797) );
  SDFFARX1 InstQueue_reg_12__6_ ( .D(n2683), .SI(n4554), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3560), .Q(n4557), .QN(n3796) );
  SDFFARX1 InstQueue_reg_12__5_ ( .D(n2684), .SI(n4551), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3560), .Q(n4554), .QN(n3795) );
  SDFFARX1 InstQueue_reg_12__4_ ( .D(n2685), .SI(n4547), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3560), .Q(n4551), .QN(n3794) );
  SDFFARX1 InstQueue_reg_10__7_ ( .D(n2698), .SI(n2852), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3557), .Q(n2853), .QN(n3781) );
  SDFFARX1 InstQueue_reg_10__6_ ( .D(n2699), .SI(n2851), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3557), .Q(n2852), .QN(n3780) );
  SDFFARX1 InstQueue_reg_10__5_ ( .D(n2700), .SI(n2850), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3557), .Q(n2851), .QN(n3779) );
  SDFFARX1 InstQueue_reg_10__4_ ( .D(n2701), .SI(n2849), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3557), .Q(n2850), .QN(n3778) );
  SDFFARX1 InstQueue_reg_8__7_ ( .D(n2714), .SI(n4446), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3555), .Q(test_so12), .QN(n3765) );
  SDFFARX1 InstQueue_reg_8__6_ ( .D(n2715), .SI(n4443), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3555), .Q(n4446), .QN(n3764) );
  SDFFARX1 InstQueue_reg_8__5_ ( .D(n2716), .SI(n4439), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3554), .Q(n4443), .QN(n3763) );
  SDFFARX1 InstQueue_reg_8__4_ ( .D(n2717), .SI(n4436), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3554), .Q(n4439), .QN(n3762) );
  SDFFARX1 InstQueue_reg_6__7_ ( .D(n2730), .SI(n2881), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3552), .Q(n2882), .QN(n3749) );
  SDFFARX1 InstQueue_reg_6__6_ ( .D(n2731), .SI(n2880), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3552), .Q(n2881), .QN(n3748) );
  SDFFARX1 InstQueue_reg_6__5_ ( .D(n2732), .SI(n2879), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3552), .Q(n2880), .QN(n3747) );
  SDFFARX1 InstQueue_reg_6__4_ ( .D(n2733), .SI(n2886), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3552), .Q(n2879), .QN(n3746) );
  SDFFARX1 InstQueue_reg_13__7_ ( .D(n2674), .SI(n4590), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3561), .Q(n4593), .QN(n3805) );
  SDFFARX1 InstQueue_reg_13__6_ ( .D(n2675), .SI(n4587), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3561), .Q(n4590), .QN(n3804) );
  SDFFARX1 InstQueue_reg_13__5_ ( .D(n2676), .SI(n4584), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3561), .Q(n4587), .QN(n3803) );
  SDFFARX1 InstQueue_reg_9__7_ ( .D(n2706), .SI(n4477), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3556), .Q(n4480), .QN(n3773) );
  SDFFARX1 InstQueue_reg_9__6_ ( .D(n2707), .SI(n4474), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3556), .Q(n4477), .QN(n3772) );
  SDFFARX1 InstQueue_reg_9__5_ ( .D(n2708), .SI(n4471), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3556), .Q(n4474), .QN(n3771) );
  SDFFARX1 InstQueue_reg_9__4_ ( .D(n2709), .SI(n4467), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3556), .Q(n4471), .QN(n3770) );
  SDFFARX1 InstQueue_reg_3__7_ ( .D(n2754), .SI(n2919), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3548), .Q(n2920), .QN(n3725) );
  SDFFARX1 InstQueue_reg_3__6_ ( .D(n2755), .SI(test_si11), .SE(test_se), 
        .CLK(CLOCK), .RSTB(n3548), .Q(n2919), .QN(n3724) );
  SDFFARX1 InstQueue_reg_3__5_ ( .D(n2756), .SI(n2917), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3548), .Q(test_so10), .QN(n3723) );
  SDFFARX1 InstQueue_reg_15__7_ ( .D(n2658), .SI(n2914), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3564), .Q(n2915), .QN(n3821) );
  SDFFARX1 InstQueue_reg_15__6_ ( .D(n2659), .SI(n2913), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3564), .Q(n2914), .QN(n3820) );
  SDFFARX1 InstQueue_reg_15__5_ ( .D(n2660), .SI(n2912), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3564), .Q(n2913), .QN(n3819) );
  SDFFARX1 InstQueue_reg_11__7_ ( .D(n2690), .SI(n2909), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3559), .Q(n2910), .QN(n3789) );
  SDFFARX1 InstQueue_reg_11__6_ ( .D(n2691), .SI(n2908), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3559), .Q(n2909), .QN(n3788) );
  SDFFARX1 InstQueue_reg_11__5_ ( .D(n2692), .SI(test_si14), .SE(test_se), 
        .CLK(CLOCK), .RSTB(n3558), .Q(n2908), .QN(n3787) );
  SDFFARX1 InstQueue_reg_11__4_ ( .D(n2693), .SI(n2927), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3558), .Q(test_so13), .QN(n3786) );
  SDFFARX1 InstQueue_reg_7__7_ ( .D(n2722), .SI(n2905), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3553), .Q(n2906), .QN(n3757) );
  SDFFARX1 InstQueue_reg_7__6_ ( .D(n2723), .SI(n2904), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3553), .Q(n2905), .QN(n3756) );
  SDFFARX1 InstQueue_reg_7__5_ ( .D(n2724), .SI(n2903), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3553), .Q(n2904), .QN(n3755) );
  SDFFARX1 InstQueue_reg_7__4_ ( .D(n2725), .SI(n2902), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3553), .Q(n2903), .QN(n3754) );
  SDFFARX1 EBX_reg_1_ ( .D(n2824), .SI(EBX_0_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3608), .Q(EBX_1_), .QN() );
  SDFFARX1 EBX_reg_2_ ( .D(n2823), .SI(EBX_1_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3608), .Q(EBX_2_), .QN() );
  SDFFARX1 EBX_reg_3_ ( .D(n2822), .SI(EBX_2_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3607), .Q(EBX_3_), .QN() );
  SDFFARX1 EBX_reg_4_ ( .D(n2821), .SI(EBX_3_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3607), .Q(EBX_4_), .QN() );
  SDFFARX1 EBX_reg_5_ ( .D(n2820), .SI(EBX_4_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3607), .Q(EBX_5_), .QN() );
  SDFFARX1 EBX_reg_6_ ( .D(n2819), .SI(EBX_5_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3607), .Q(EBX_6_), .QN() );
  SDFFARX1 EBX_reg_7_ ( .D(n2818), .SI(EBX_6_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3607), .Q(EBX_7_), .QN() );
  SDFFARX1 EAX_reg_0_ ( .D(n2588), .SI(Datao[30]), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3579), .Q(N3346), .QN(n3838) );
  SDFFARX1 InstAddrPointer_reg_5_ ( .D(n2521), .SI(InstAddrPointer_4_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3601), .Q(InstAddrPointer_5_), .QN(n3870) );
  SDFFARX1 InstAddrPointer_reg_3_ ( .D(n2523), .SI(InstAddrPointer_2_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3590), .Q(InstAddrPointer_3_), .QN(n3865) );
  SDFFARX1 InstAddrPointer_reg_4_ ( .D(n2522), .SI(InstAddrPointer_3_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3589), .Q(InstAddrPointer_4_), .QN(n3864) );
  SDFFARX1 InstAddrPointer_reg_6_ ( .D(n2520), .SI(InstAddrPointer_5_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3589), .Q(InstAddrPointer_6_), .QN(n3863) );
  SDFFARX1 InstAddrPointer_reg_7_ ( .D(n2519), .SI(InstAddrPointer_6_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3589), .Q(test_so7), .QN(n3862) );
  SDFFARX1 InstAddrPointer_reg_2_ ( .D(n2524), .SI(InstAddrPointer_1_), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3590), .Q(InstAddrPointer_2_), .QN(n3866) );
  SDFFARX1 EBX_reg_0_ ( .D(n2825), .SI(EAX_31_), .SE(test_se), .CLK(CLOCK), 
        .RSTB(n3608), .Q(EBX_0_), .QN() );
  SDFFARX1 InstAddrPointer_reg_1_ ( .D(n2525), .SI(N3469), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3590), .Q(InstAddrPointer_1_), .QN(n3867) );
  SDFFARX1 InstQueue_reg_14__3_ ( .D(n2670), .SI(n2878), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3562), .Q(n2871), .QN(n3809) );
  SDFFARX1 InstQueue_reg_14__2_ ( .D(n2671), .SI(test_si15), .SE(test_se), 
        .CLK(CLOCK), .RSTB(n3562), .Q(n2878), .QN(n3808) );
  SDFFARX1 InstQueue_reg_14__1_ ( .D(n2672), .SI(n2876), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3562), .Q(test_so14), .QN(n3807) );
  SDFFARX1 InstQueue_reg_14__0_ ( .D(n2673), .SI(n4593), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3562), .Q(n2876), .QN(n3806) );
  SDFFARX1 InstQueue_reg_1__4_ ( .D(n2773), .SI(n4241), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3545), .Q(n4244), .QN(n3706) );
  SDFFARX1 InstQueue_reg_1__3_ ( .D(n2774), .SI(n4238), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3545), .Q(n4241), .QN(n3705) );
  SDFFARX1 InstQueue_reg_1__2_ ( .D(n2775), .SI(n4234), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3545), .Q(n4238), .QN(n3704) );
  SDFFARX1 InstQueue_reg_1__1_ ( .D(n2776), .SI(test_si10), .SE(test_se), 
        .CLK(CLOCK), .RSTB(n3544), .Q(n4234), .QN(n3703) );
  SDFFARX1 InstQueue_reg_1__0_ ( .D(n2777), .SI(N2555), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3544), .Q(test_so9), .QN(n3702) );
  SDFFARX1 InstQueue_reg_0__3_ ( .D(n2782), .SI(N2550), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3543), .Q(N2551), .QN(n3697) );
  SDFFARX1 InstQueue_reg_0__2_ ( .D(n2783), .SI(N2549), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3543), .Q(N2550), .QN(n3696) );
  SDFFARX1 InstQueue_reg_0__1_ ( .D(n2784), .SI(N2548), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3543), .Q(N2549), .QN(n3695) );
  SDFFARX1 InstQueue_reg_0__0_ ( .D(n2785), .SI(N3989), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3543), .Q(N2548), .QN(n3694) );
  SDFFARX1 InstQueue_reg_5__3_ ( .D(n2742), .SI(n4352), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3550), .Q(n4355), .QN(n3737) );
  SDFFARX1 InstQueue_reg_5__2_ ( .D(n2743), .SI(n4349), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3550), .Q(n4352), .QN(n3736) );
  SDFFARX1 InstQueue_reg_5__1_ ( .D(n2744), .SI(n4345), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3550), .Q(n4349), .QN(n3735) );
  SDFFARX1 InstQueue_reg_5__0_ ( .D(n2745), .SI(n4336), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3550), .Q(n4345), .QN(n3734) );
  SDFFARX1 InstQueue_reg_4__3_ ( .D(n2750), .SI(n4320), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3549), .Q(n4323), .QN(n3729) );
  SDFFARX1 InstQueue_reg_4__2_ ( .D(n2751), .SI(n4317), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3549), .Q(n4320), .QN(n3728) );
  SDFFARX1 InstQueue_reg_4__1_ ( .D(n2752), .SI(n4313), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3548), .Q(n4317), .QN(n3727) );
  SDFFARX1 InstQueue_reg_4__0_ ( .D(n2753), .SI(n2920), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3548), .Q(n4313), .QN(n3726) );
  SDFFARX1 InstQueue_reg_2__3_ ( .D(n2766), .SI(n2862), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3546), .Q(n2863), .QN(n3713) );
  SDFFARX1 InstQueue_reg_2__2_ ( .D(n2767), .SI(n2861), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3546), .Q(n2862), .QN(n3712) );
  SDFFARX1 InstQueue_reg_2__1_ ( .D(n2768), .SI(n2848), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3546), .Q(n2861), .QN(n3711) );
  SDFFARX1 InstQueue_reg_2__0_ ( .D(n2769), .SI(n4253), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3546), .Q(n2848), .QN(n3710) );
  SDFFARX1 InstQueue_reg_12__3_ ( .D(n2686), .SI(n4544), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3559), .Q(n4547), .QN(n3793) );
  SDFFARX1 InstQueue_reg_12__2_ ( .D(n2687), .SI(n4541), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3559), .Q(n4544), .QN(n3792) );
  SDFFARX1 InstQueue_reg_12__1_ ( .D(n2688), .SI(n4537), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3559), .Q(n4541), .QN(n3791) );
  SDFFARX1 InstQueue_reg_12__0_ ( .D(n2689), .SI(n2910), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3559), .Q(n4537), .QN(n3790) );
  SDFFARX1 InstQueue_reg_10__3_ ( .D(n2702), .SI(n2856), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3557), .Q(n2849), .QN(n3777) );
  SDFFARX1 InstQueue_reg_10__2_ ( .D(n2703), .SI(n2855), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3557), .Q(n2856), .QN(n3776) );
  SDFFARX1 InstQueue_reg_10__1_ ( .D(n2704), .SI(n2854), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3556), .Q(n2855), .QN(n3775) );
  SDFFARX1 InstQueue_reg_10__0_ ( .D(n2705), .SI(n4480), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3556), .Q(n2854), .QN(n3774) );
  SDFFARX1 InstQueue_reg_8__3_ ( .D(n2718), .SI(n4433), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3554), .Q(n4436), .QN(n3761) );
  SDFFARX1 InstQueue_reg_8__2_ ( .D(n2719), .SI(n4430), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3554), .Q(n4433), .QN(n3760) );
  SDFFARX1 InstQueue_reg_8__1_ ( .D(n2720), .SI(n4426), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3554), .Q(n4430), .QN(n3759) );
  SDFFARX1 InstQueue_reg_8__0_ ( .D(n2721), .SI(n2906), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3554), .Q(n4426), .QN(n3758) );
  SDFFARX1 InstQueue_reg_6__3_ ( .D(n2734), .SI(test_si12), .SE(test_se), 
        .CLK(CLOCK), .RSTB(n3551), .Q(n2886), .QN(n3745) );
  SDFFARX1 InstQueue_reg_6__2_ ( .D(n2735), .SI(n2884), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3551), .Q(test_so11), .QN(n3744) );
  SDFFARX1 InstQueue_reg_6__1_ ( .D(n2736), .SI(n2869), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3551), .Q(n2884), .QN(n3743) );
  SDFFARX1 InstQueue_reg_6__0_ ( .D(n2737), .SI(n4368), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3551), .Q(n2869), .QN(n3742) );
  SDFFARX1 InstQueue_reg_13__4_ ( .D(n2677), .SI(n4580), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3561), .Q(n4584), .QN(n3802) );
  SDFFARX1 InstQueue_reg_13__3_ ( .D(n2678), .SI(n4577), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3561), .Q(n4580), .QN(n3801) );
  SDFFARX1 InstQueue_reg_13__2_ ( .D(n2679), .SI(n4574), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3561), .Q(n4577), .QN(n3800) );
  SDFFARX1 InstQueue_reg_13__1_ ( .D(n2680), .SI(n4570), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3560), .Q(n4574), .QN(n3799) );
  SDFFARX1 InstQueue_reg_13__0_ ( .D(n2681), .SI(n4560), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3560), .Q(n4570), .QN(n3798) );
  SDFFARX1 InstQueue_reg_9__3_ ( .D(n2710), .SI(n4464), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3555), .Q(n4467), .QN(n3769) );
  SDFFARX1 InstQueue_reg_9__2_ ( .D(n2711), .SI(n4461), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3555), .Q(n4464), .QN(n3768) );
  SDFFARX1 InstQueue_reg_9__1_ ( .D(n2712), .SI(n4457), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3555), .Q(n4461), .QN(n3767) );
  SDFFARX1 InstQueue_reg_9__0_ ( .D(n2713), .SI(test_si13), .SE(test_se), 
        .CLK(CLOCK), .RSTB(n3555), .Q(n4457), .QN(n3766) );
  SDFFARX1 InstQueue_reg_3__4_ ( .D(n2757), .SI(n2933), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3548), .Q(n2917), .QN(n3722) );
  SDFFARX1 InstQueue_reg_3__3_ ( .D(n2758), .SI(n2932), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3547), .Q(n2933), .QN(n3721) );
  SDFFARX1 InstQueue_reg_3__2_ ( .D(n2759), .SI(n2931), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3547), .Q(n2932), .QN(n3720) );
  SDFFARX1 InstQueue_reg_3__1_ ( .D(n2760), .SI(n2916), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3547), .Q(n2931), .QN(n3719) );
  SDFFARX1 InstQueue_reg_3__0_ ( .D(n2761), .SI(n2860), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3547), .Q(n2916), .QN(n3718) );
  SDFFARX1 InstQueue_reg_15__4_ ( .D(n2661), .SI(n2911), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3564), .Q(n2912), .QN(n3818) );
  SDFFARX1 InstQueue_reg_15__3_ ( .D(n2662), .SI(n2930), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3563), .Q(n2911), .QN(n3817) );
  SDFFARX1 InstQueue_reg_15__2_ ( .D(n2663), .SI(n2929), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3563), .Q(n2930), .QN(n3816) );
  SDFFARX1 InstQueue_reg_15__1_ ( .D(n2664), .SI(n2928), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3563), .Q(n2929), .QN(n3815) );
  SDFFARX1 InstQueue_reg_15__0_ ( .D(n2665), .SI(n2875), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3563), .Q(n2928), .QN(n3814) );
  SDFFARX1 InstQueue_reg_11__3_ ( .D(n2694), .SI(n2926), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3558), .Q(n2927), .QN(n3785) );
  SDFFARX1 InstQueue_reg_11__2_ ( .D(n2695), .SI(n2925), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3558), .Q(n2926), .QN(n3784) );
  SDFFARX1 InstQueue_reg_11__1_ ( .D(n2696), .SI(n2924), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3558), .Q(n2925), .QN(n3783) );
  SDFFARX1 InstQueue_reg_11__0_ ( .D(n2697), .SI(n2853), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3558), .Q(n2924), .QN(n3782) );
  SDFFARX1 InstQueue_reg_7__3_ ( .D(n2726), .SI(n2923), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3553), .Q(n2902), .QN(n3753) );
  SDFFARX1 InstQueue_reg_7__2_ ( .D(n2727), .SI(n2922), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3553), .Q(n2923), .QN(n3752) );
  SDFFARX1 InstQueue_reg_7__1_ ( .D(n2728), .SI(n2921), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3552), .Q(n2922), .QN(n3751) );
  SDFFARX1 InstQueue_reg_7__0_ ( .D(n2729), .SI(n2882), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3552), .Q(n2921), .QN(n3750) );
  SDFFARX1 InstQueueRd_Addr_reg_1_ ( .D(n2792), .SI(N2737), .SE(test_se), 
        .CLK(CLOCK), .RSTB(n3580), .Q(InstQueueRd_Addr[1]), .QN(n1550) );
  SDFFARX1 InstAddrPointer_reg_0_ ( .D(n2526), .SI(n2870), .SE(test_se), .CLK(
        CLOCK), .RSTB(n3590), .Q(N3469), .QN(n1557) );
  SDFFARX1 InstQueueRd_Addr_reg_0_ ( .D(n2793), .SI(N3467), .SE(test_se), 
        .CLK(CLOCK), .RSTB(n3580), .Q(N2737), .QN(n1552) );
  SDFFARX1 InstQueueRd_Addr_reg_2_ ( .D(n2791), .SI(InstQueueRd_Addr[1]), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3580), .Q(InstQueueRd_Addr[2]), .QN(
        n3839) );
  SDFFARX1 InstQueueRd_Addr_reg_3_ ( .D(n2831), .SI(InstQueueRd_Addr[2]), .SE(
        test_se), .CLK(CLOCK), .RSTB(n3602), .Q(InstQueueRd_Addr[3]), .QN(
        n1548) );
  XNOR2X1 U2310 ( .IN1(Datai[23]), .IN2(n2975), .Q(n2843) );
  AND2X1 U2311 ( .IN1(N1764), .IN2(mult_add_463_aco_A_0_), .Q(n2846) );
  XNOR2X1 U2312 ( .IN1(add_495_carry[4]), .IN2(InstQueueRd_Addr[4]), .Q(n2883)
         );
  OR2X1 U2313 ( .IN1(n1548), .IN2(n2870), .Q(n2887) );
  INVX0 U2314 ( .IN(Datai[13]), .QN(n2934) );
  INVX0 U2315 ( .IN(n2934), .QN(n2935) );
  INVX0 U2316 ( .IN(Datai[10]), .QN(n2936) );
  INVX0 U2317 ( .IN(n2936), .QN(n2937) );
  INVX0 U2318 ( .IN(Datai[14]), .QN(n2938) );
  INVX0 U2319 ( .IN(n2938), .QN(n2939) );
  INVX0 U2320 ( .IN(Datai[8]), .QN(n2940) );
  INVX0 U2321 ( .IN(n2940), .QN(n2941) );
  INVX0 U2322 ( .IN(Datai[11]), .QN(n2942) );
  INVX0 U2323 ( .IN(n2942), .QN(n2943) );
  INVX0 U2324 ( .IN(Datai[9]), .QN(n2944) );
  INVX0 U2325 ( .IN(n2944), .QN(n2945) );
  INVX0 U2326 ( .IN(Datai[12]), .QN(n2946) );
  INVX0 U2327 ( .IN(n2946), .QN(n2947) );
  INVX0 U2328 ( .IN(READY_n), .QN(n2948) );
  INVX0 U2329 ( .IN(n2948), .QN(n2949) );
  NBUFFX2 U2330 ( .IN(n3459), .Q(n3458) );
  NBUFFX2 U2331 ( .IN(n3460), .Q(n3457) );
  NBUFFX2 U2332 ( .IN(n3460), .Q(n3456) );
  NBUFFX2 U2333 ( .IN(n3461), .Q(n3455) );
  NBUFFX2 U2334 ( .IN(n3461), .Q(n3454) );
  NBUFFX2 U2335 ( .IN(n3474), .Q(n3466) );
  NBUFFX2 U2336 ( .IN(n3473), .Q(n3468) );
  NBUFFX2 U2337 ( .IN(n3473), .Q(n3469) );
  NBUFFX2 U2338 ( .IN(n3472), .Q(n3470) );
  NBUFFX2 U2339 ( .IN(n3474), .Q(n3467) );
  NBUFFX2 U2340 ( .IN(n3472), .Q(n3471) );
  INVX0 U2341 ( .IN(n3195), .QN(n3185) );
  INVX0 U2342 ( .IN(n3184), .QN(n3194) );
  INVX0 U2343 ( .IN(n3203), .QN(n3187) );
  INVX0 U2344 ( .IN(n3203), .QN(n3186) );
  INVX0 U2345 ( .IN(n3203), .QN(n3188) );
  INVX0 U2346 ( .IN(n3204), .QN(n3193) );
  INVX0 U2347 ( .IN(n3204), .QN(n3192) );
  INVX0 U2348 ( .IN(n3204), .QN(n3191) );
  INVX0 U2349 ( .IN(n3203), .QN(n3190) );
  INVX0 U2350 ( .IN(n3203), .QN(n3189) );
  INVX0 U2351 ( .IN(n3137), .QN(n3140) );
  INVX0 U2352 ( .IN(n3146), .QN(n3141) );
  INVX0 U2353 ( .IN(n3146), .QN(n3142) );
  INVX0 U2354 ( .IN(n3145), .QN(n3143) );
  INVX0 U2355 ( .IN(n3145), .QN(n3144) );
  NBUFFX2 U2356 ( .IN(n3462), .Q(n3453) );
  NBUFFX2 U2357 ( .IN(n3463), .Q(n3462) );
  NBUFFX2 U2358 ( .IN(n3475), .Q(n3465) );
  NBUFFX2 U2359 ( .IN(n3476), .Q(n3475) );
  NBUFFX2 U2360 ( .IN(n3447), .Q(n3446) );
  NBUFFX2 U2361 ( .IN(n3448), .Q(n3445) );
  NBUFFX2 U2362 ( .IN(n3448), .Q(n3444) );
  NBUFFX2 U2363 ( .IN(n3449), .Q(n3443) );
  NBUFFX2 U2364 ( .IN(n3449), .Q(n3442) );
  NBUFFX2 U2365 ( .IN(n3477), .Q(n3473) );
  NBUFFX2 U2366 ( .IN(n3464), .Q(n3460) );
  NBUFFX2 U2367 ( .IN(n3477), .Q(n3472) );
  NBUFFX2 U2368 ( .IN(n3463), .Q(n3461) );
  NBUFFX2 U2369 ( .IN(n3464), .Q(n3459) );
  NBUFFX2 U2370 ( .IN(n3476), .Q(n3474) );
  INVX0 U2371 ( .IN(n3182), .QN(n3195) );
  INVX0 U2372 ( .IN(n3183), .QN(n3197) );
  INVX0 U2373 ( .IN(n3183), .QN(n3198) );
  INVX0 U2374 ( .IN(n3183), .QN(n3199) );
  INVX0 U2375 ( .IN(n3183), .QN(n3202) );
  INVX0 U2376 ( .IN(n3183), .QN(n3201) );
  INVX0 U2377 ( .IN(n3183), .QN(n3196) );
  INVX0 U2378 ( .IN(n3183), .QN(n3200) );
  INVX0 U2379 ( .IN(n3183), .QN(n3203) );
  INVX0 U2380 ( .IN(n3183), .QN(n3204) );
  NBUFFX2 U2381 ( .IN(n3646), .Q(n3542) );
  NBUFFX2 U2382 ( .IN(n3646), .Q(n3543) );
  NBUFFX2 U2383 ( .IN(n3645), .Q(n3544) );
  NBUFFX2 U2384 ( .IN(n3645), .Q(n3545) );
  NBUFFX2 U2385 ( .IN(n3644), .Q(n3546) );
  NBUFFX2 U2386 ( .IN(n3644), .Q(n3547) );
  NBUFFX2 U2387 ( .IN(n3643), .Q(n3548) );
  NBUFFX2 U2388 ( .IN(n3643), .Q(n3549) );
  NBUFFX2 U2389 ( .IN(n3642), .Q(n3550) );
  NBUFFX2 U2390 ( .IN(n3642), .Q(n3551) );
  NBUFFX2 U2391 ( .IN(n3641), .Q(n3552) );
  NBUFFX2 U2392 ( .IN(n3641), .Q(n3553) );
  NBUFFX2 U2393 ( .IN(n3640), .Q(n3554) );
  NBUFFX2 U2394 ( .IN(n3640), .Q(n3555) );
  NBUFFX2 U2395 ( .IN(n3639), .Q(n3556) );
  NBUFFX2 U2396 ( .IN(n3639), .Q(n3557) );
  NBUFFX2 U2397 ( .IN(n3638), .Q(n3558) );
  NBUFFX2 U2398 ( .IN(n3638), .Q(n3559) );
  NBUFFX2 U2399 ( .IN(n3637), .Q(n3560) );
  NBUFFX2 U2400 ( .IN(n3637), .Q(n3561) );
  NBUFFX2 U2401 ( .IN(n3636), .Q(n3562) );
  NBUFFX2 U2402 ( .IN(n3636), .Q(n3563) );
  NBUFFX2 U2403 ( .IN(n3635), .Q(n3564) );
  NBUFFX2 U2404 ( .IN(n3635), .Q(n3565) );
  NBUFFX2 U2405 ( .IN(n3634), .Q(n3566) );
  NBUFFX2 U2406 ( .IN(n3634), .Q(n3567) );
  NBUFFX2 U2407 ( .IN(n3633), .Q(n3568) );
  NBUFFX2 U2408 ( .IN(n3633), .Q(n3569) );
  NBUFFX2 U2409 ( .IN(n3632), .Q(n3570) );
  NBUFFX2 U2410 ( .IN(n3632), .Q(n3571) );
  NBUFFX2 U2411 ( .IN(n3631), .Q(n3572) );
  NBUFFX2 U2412 ( .IN(n3631), .Q(n3573) );
  NBUFFX2 U2413 ( .IN(n3630), .Q(n3574) );
  NBUFFX2 U2414 ( .IN(n3630), .Q(n3575) );
  NBUFFX2 U2415 ( .IN(n3629), .Q(n3576) );
  NBUFFX2 U2416 ( .IN(n3629), .Q(n3577) );
  NBUFFX2 U2417 ( .IN(n3628), .Q(n3578) );
  NBUFFX2 U2418 ( .IN(n3628), .Q(n3579) );
  NBUFFX2 U2419 ( .IN(n3627), .Q(n3580) );
  NBUFFX2 U2420 ( .IN(n3627), .Q(n3581) );
  NBUFFX2 U2421 ( .IN(n3626), .Q(n3582) );
  NBUFFX2 U2422 ( .IN(n3626), .Q(n3583) );
  NBUFFX2 U2423 ( .IN(n3625), .Q(n3584) );
  NBUFFX2 U2424 ( .IN(n3625), .Q(n3585) );
  NBUFFX2 U2425 ( .IN(n3624), .Q(n3586) );
  NBUFFX2 U2426 ( .IN(n3624), .Q(n3587) );
  NBUFFX2 U2427 ( .IN(n3623), .Q(n3588) );
  NBUFFX2 U2428 ( .IN(n3623), .Q(n3589) );
  NBUFFX2 U2429 ( .IN(n3622), .Q(n3590) );
  NBUFFX2 U2430 ( .IN(n3622), .Q(n3591) );
  NBUFFX2 U2431 ( .IN(n3621), .Q(n3592) );
  NBUFFX2 U2432 ( .IN(n3621), .Q(n3593) );
  NBUFFX2 U2433 ( .IN(n3620), .Q(n3594) );
  NBUFFX2 U2434 ( .IN(n3620), .Q(n3595) );
  NBUFFX2 U2435 ( .IN(n3619), .Q(n3596) );
  NBUFFX2 U2436 ( .IN(n3619), .Q(n3597) );
  NBUFFX2 U2437 ( .IN(n3618), .Q(n3598) );
  NBUFFX2 U2438 ( .IN(n3618), .Q(n3599) );
  NBUFFX2 U2439 ( .IN(n3617), .Q(n3600) );
  NBUFFX2 U2440 ( .IN(n3617), .Q(n3601) );
  NBUFFX2 U2441 ( .IN(n3616), .Q(n3602) );
  NBUFFX2 U2442 ( .IN(n3616), .Q(n3603) );
  NBUFFX2 U2443 ( .IN(n3615), .Q(n3604) );
  NBUFFX2 U2444 ( .IN(n3615), .Q(n3605) );
  INVX0 U2445 ( .IN(n3113), .QN(n3108) );
  INVX0 U2446 ( .IN(n3125), .QN(n3121) );
  INVX0 U2447 ( .IN(n3163), .QN(n3164) );
  INVX0 U2448 ( .IN(n3170), .QN(n3166) );
  INVX0 U2449 ( .IN(n3170), .QN(n3165) );
  INVX0 U2450 ( .IN(n3896), .QN(n3146) );
  INVX0 U2451 ( .IN(n3135), .QN(n3145) );
  INVX0 U2452 ( .IN(n3133), .QN(n3150) );
  INVX0 U2453 ( .IN(n3135), .QN(n3156) );
  INVX0 U2454 ( .IN(n3135), .QN(n3155) );
  INVX0 U2455 ( .IN(n3132), .QN(n3149) );
  INVX0 U2456 ( .IN(n3135), .QN(n3154) );
  INVX0 U2457 ( .IN(n3114), .QN(n3109) );
  INVX0 U2458 ( .IN(n3169), .QN(n3168) );
  INVX0 U2459 ( .IN(n3169), .QN(n3167) );
  INVX0 U2460 ( .IN(n3134), .QN(n3153) );
  INVX0 U2461 ( .IN(n3132), .QN(n3147) );
  INVX0 U2462 ( .IN(n3132), .QN(n3148) );
  INVX0 U2463 ( .IN(n3134), .QN(n3152) );
  INVX0 U2464 ( .IN(n3134), .QN(n3151) );
  NBUFFX2 U2465 ( .IN(n3272), .Q(n3270) );
  NBUFFX2 U2466 ( .IN(n3273), .Q(n3269) );
  NBUFFX2 U2467 ( .IN(n3273), .Q(n3268) );
  NBUFFX2 U2468 ( .IN(n3274), .Q(n3267) );
  NBUFFX2 U2469 ( .IN(n3274), .Q(n3266) );
  NBUFFX2 U2470 ( .IN(n3272), .Q(n3271) );
  NBUFFX2 U2471 ( .IN(n3275), .Q(n3264) );
  NBUFFX2 U2472 ( .IN(n3275), .Q(n3265) );
  NBUFFX2 U2473 ( .IN(n3335), .Q(n3325) );
  NBUFFX2 U2474 ( .IN(n3335), .Q(n3326) );
  NBUFFX2 U2475 ( .IN(n3334), .Q(n3327) );
  NBUFFX2 U2476 ( .IN(n3333), .Q(n3329) );
  NBUFFX2 U2477 ( .IN(n3332), .Q(n3331) );
  NBUFFX2 U2478 ( .IN(n3334), .Q(n3328) );
  NBUFFX2 U2479 ( .IN(n3333), .Q(n3330) );
  NBUFFX2 U2480 ( .IN(n3284), .Q(n3282) );
  NBUFFX2 U2481 ( .IN(n3308), .Q(n3306) );
  NBUFFX2 U2482 ( .IN(n3285), .Q(n3281) );
  NBUFFX2 U2483 ( .IN(n3309), .Q(n3305) );
  NBUFFX2 U2484 ( .IN(n3285), .Q(n3280) );
  NBUFFX2 U2485 ( .IN(n3309), .Q(n3304) );
  NBUFFX2 U2486 ( .IN(n3286), .Q(n3279) );
  NBUFFX2 U2487 ( .IN(n3310), .Q(n3303) );
  NBUFFX2 U2488 ( .IN(n3286), .Q(n3278) );
  NBUFFX2 U2489 ( .IN(n3310), .Q(n3302) );
  NBUFFX2 U2490 ( .IN(n3284), .Q(n3283) );
  NBUFFX2 U2491 ( .IN(n3308), .Q(n3307) );
  NBUFFX2 U2492 ( .IN(n3287), .Q(n3276) );
  NBUFFX2 U2493 ( .IN(n3311), .Q(n3300) );
  NBUFFX2 U2494 ( .IN(n3287), .Q(n3277) );
  NBUFFX2 U2495 ( .IN(n3311), .Q(n3301) );
  NBUFFX2 U2496 ( .IN(n3296), .Q(n3294) );
  NBUFFX2 U2497 ( .IN(n3320), .Q(n3318) );
  NBUFFX2 U2498 ( .IN(n3297), .Q(n3293) );
  NBUFFX2 U2499 ( .IN(n3321), .Q(n3317) );
  NBUFFX2 U2500 ( .IN(n3297), .Q(n3292) );
  NBUFFX2 U2501 ( .IN(n3321), .Q(n3316) );
  NBUFFX2 U2502 ( .IN(n3298), .Q(n3291) );
  NBUFFX2 U2503 ( .IN(n3322), .Q(n3315) );
  NBUFFX2 U2504 ( .IN(n3298), .Q(n3290) );
  NBUFFX2 U2505 ( .IN(n3322), .Q(n3314) );
  NBUFFX2 U2506 ( .IN(n3296), .Q(n3295) );
  NBUFFX2 U2507 ( .IN(n3320), .Q(n3319) );
  NBUFFX2 U2508 ( .IN(n3299), .Q(n3288) );
  NBUFFX2 U2509 ( .IN(n3323), .Q(n3312) );
  NBUFFX2 U2510 ( .IN(n3299), .Q(n3289) );
  NBUFFX2 U2511 ( .IN(n3323), .Q(n3313) );
  NBUFFX2 U2512 ( .IN(n4832), .Q(n3477) );
  NBUFFX2 U2513 ( .IN(n4832), .Q(n3476) );
  NBUFFX2 U2514 ( .IN(n4831), .Q(n3463) );
  NBUFFX2 U2515 ( .IN(n4831), .Q(n3464) );
  NBUFFX2 U2516 ( .IN(n3452), .Q(n3448) );
  NBUFFX2 U2517 ( .IN(n3451), .Q(n3449) );
  NBUFFX2 U2518 ( .IN(n3452), .Q(n3447) );
  NBUFFX2 U2519 ( .IN(n3450), .Q(n3441) );
  NBUFFX2 U2520 ( .IN(n3451), .Q(n3450) );
  INVX0 U2521 ( .IN(n2952), .QN(n3102) );
  INVX0 U2522 ( .IN(n2951), .QN(n3103) );
  NBUFFX2 U2523 ( .IN(n4824), .Q(n3407) );
  NBUFFX2 U2524 ( .IN(n4824), .Q(n3406) );
  NBUFFX2 U2525 ( .IN(n4824), .Q(n3405) );
  NBUFFX2 U2526 ( .IN(n4824), .Q(n3408) );
  NBUFFX2 U2527 ( .IN(n4824), .Q(n3409) );
  NBUFFX2 U2528 ( .IN(n4824), .Q(n3410) );
  NBUFFX2 U2529 ( .IN(n3373), .Q(n3372) );
  NBUFFX2 U2530 ( .IN(n3374), .Q(n3371) );
  NBUFFX2 U2531 ( .IN(n3374), .Q(n3370) );
  NBUFFX2 U2532 ( .IN(n3375), .Q(n3369) );
  NBUFFX2 U2533 ( .IN(n3375), .Q(n3368) );
  NBUFFX2 U2534 ( .IN(n3365), .Q(n3357) );
  NBUFFX2 U2535 ( .IN(n3365), .Q(n3358) );
  NBUFFX2 U2536 ( .IN(n3364), .Q(n3359) );
  NBUFFX2 U2537 ( .IN(n3364), .Q(n3360) );
  NBUFFX2 U2538 ( .IN(n3363), .Q(n3361) );
  NBUFFX2 U2539 ( .IN(n3523), .Q(n3516) );
  NBUFFX2 U2540 ( .IN(n3522), .Q(n3517) );
  NBUFFX2 U2541 ( .IN(n3522), .Q(n3518) );
  NBUFFX2 U2542 ( .IN(n3521), .Q(n3519) );
  NBUFFX2 U2543 ( .IN(n3521), .Q(n3520) );
  NBUFFX2 U2544 ( .IN(n3523), .Q(n3515) );
  NBUFFX2 U2545 ( .IN(n3486), .Q(n3484) );
  NBUFFX2 U2546 ( .IN(n3510), .Q(n3508) );
  NBUFFX2 U2547 ( .IN(n3487), .Q(n3483) );
  NBUFFX2 U2548 ( .IN(n3511), .Q(n3507) );
  NBUFFX2 U2549 ( .IN(n3487), .Q(n3482) );
  NBUFFX2 U2550 ( .IN(n3511), .Q(n3506) );
  NBUFFX2 U2551 ( .IN(n3488), .Q(n3481) );
  NBUFFX2 U2552 ( .IN(n3512), .Q(n3505) );
  NBUFFX2 U2553 ( .IN(n3488), .Q(n3480) );
  NBUFFX2 U2554 ( .IN(n3512), .Q(n3504) );
  NBUFFX2 U2555 ( .IN(n3489), .Q(n3478) );
  NBUFFX2 U2556 ( .IN(n3513), .Q(n3502) );
  NBUFFX2 U2557 ( .IN(n3489), .Q(n3479) );
  NBUFFX2 U2558 ( .IN(n3513), .Q(n3503) );
  NBUFFX2 U2559 ( .IN(n3486), .Q(n3485) );
  NBUFFX2 U2560 ( .IN(n3510), .Q(n3509) );
  NBUFFX2 U2561 ( .IN(n3363), .Q(n3362) );
  INVX0 U2562 ( .IN(n3393), .QN(n3392) );
  INVX0 U2563 ( .IN(n3184), .QN(n3182) );
  INVX0 U2564 ( .IN(n3394), .QN(n3391) );
  INVX0 U2565 ( .IN(n3397), .QN(n3390) );
  INVX0 U2566 ( .IN(n3184), .QN(n3183) );
  NBUFFX2 U2567 ( .IN(n3348), .Q(n3337) );
  NBUFFX2 U2568 ( .IN(n3348), .Q(n3338) );
  NBUFFX2 U2569 ( .IN(n3347), .Q(n3339) );
  NBUFFX2 U2570 ( .IN(n3347), .Q(n3340) );
  NBUFFX2 U2571 ( .IN(n3346), .Q(n3341) );
  NBUFFX2 U2572 ( .IN(n3346), .Q(n3342) );
  NBUFFX2 U2573 ( .IN(n3345), .Q(n3343) );
  NBUFFX2 U2574 ( .IN(n3345), .Q(n3344) );
  NBUFFX2 U2575 ( .IN(n3614), .Q(n3606) );
  NBUFFX2 U2576 ( .IN(n3614), .Q(n3607) );
  NBUFFX2 U2577 ( .IN(n3613), .Q(n3608) );
  NBUFFX2 U2578 ( .IN(n3613), .Q(n3609) );
  NBUFFX2 U2579 ( .IN(n3647), .Q(n3646) );
  NBUFFX2 U2580 ( .IN(n3647), .Q(n3645) );
  NBUFFX2 U2581 ( .IN(n3648), .Q(n3644) );
  NBUFFX2 U2582 ( .IN(n3648), .Q(n3643) );
  NBUFFX2 U2583 ( .IN(n3649), .Q(n3642) );
  NBUFFX2 U2584 ( .IN(n3649), .Q(n3641) );
  NBUFFX2 U2585 ( .IN(n3650), .Q(n3640) );
  NBUFFX2 U2586 ( .IN(n3650), .Q(n3639) );
  NBUFFX2 U2587 ( .IN(n3651), .Q(n3638) );
  NBUFFX2 U2588 ( .IN(n3651), .Q(n3637) );
  NBUFFX2 U2589 ( .IN(n3652), .Q(n3636) );
  NBUFFX2 U2590 ( .IN(n3652), .Q(n3635) );
  NBUFFX2 U2591 ( .IN(n3653), .Q(n3634) );
  NBUFFX2 U2592 ( .IN(n3653), .Q(n3633) );
  NBUFFX2 U2593 ( .IN(n3654), .Q(n3632) );
  NBUFFX2 U2594 ( .IN(n3654), .Q(n3631) );
  NBUFFX2 U2595 ( .IN(n3655), .Q(n3630) );
  NBUFFX2 U2596 ( .IN(n3655), .Q(n3629) );
  NBUFFX2 U2597 ( .IN(n3656), .Q(n3628) );
  NBUFFX2 U2598 ( .IN(n3656), .Q(n3627) );
  NBUFFX2 U2599 ( .IN(n3657), .Q(n3626) );
  NBUFFX2 U2600 ( .IN(n3657), .Q(n3625) );
  NBUFFX2 U2601 ( .IN(n3658), .Q(n3624) );
  NBUFFX2 U2602 ( .IN(n3658), .Q(n3623) );
  NBUFFX2 U2603 ( .IN(n3659), .Q(n3622) );
  NBUFFX2 U2604 ( .IN(n3659), .Q(n3621) );
  NBUFFX2 U2605 ( .IN(n3660), .Q(n3620) );
  NBUFFX2 U2606 ( .IN(n3660), .Q(n3619) );
  NBUFFX2 U2607 ( .IN(n3661), .Q(n3618) );
  NBUFFX2 U2608 ( .IN(n3661), .Q(n3617) );
  NBUFFX2 U2609 ( .IN(n3662), .Q(n3616) );
  NBUFFX2 U2610 ( .IN(n3662), .Q(n3615) );
  INVX0 U2611 ( .IN(n3112), .QN(n3107) );
  INVX0 U2612 ( .IN(n3129), .QN(n3122) );
  INVX0 U2613 ( .IN(n3125), .QN(n3124) );
  INVX0 U2614 ( .IN(n3115), .QN(n3111) );
  INVX0 U2615 ( .IN(n3893), .QN(n3113) );
  INVX0 U2616 ( .IN(n3893), .QN(n3115) );
  INVX0 U2617 ( .IN(n3893), .QN(n3116) );
  INVX0 U2618 ( .IN(n3894), .QN(n3125) );
  INVX0 U2619 ( .IN(n3119), .QN(n3128) );
  INVX0 U2620 ( .IN(n3119), .QN(n3126) );
  INVX0 U2621 ( .IN(n3119), .QN(n3129) );
  INVX0 U2622 ( .IN(n3124), .QN(n3127) );
  INVX0 U2623 ( .IN(n3138), .QN(n3133) );
  INVX0 U2624 ( .IN(n3897), .QN(n3170) );
  INVX0 U2625 ( .IN(n3136), .QN(n3135) );
  INVX0 U2626 ( .IN(n3166), .QN(n3180) );
  INVX0 U2627 ( .IN(n3161), .QN(n3181) );
  INVX0 U2628 ( .IN(n3114), .QN(n3110) );
  INVX0 U2629 ( .IN(n3127), .QN(n3123) );
  INVX0 U2630 ( .IN(n3106), .QN(n3114) );
  INVX0 U2631 ( .IN(n3106), .QN(n3118) );
  INVX0 U2632 ( .IN(n3106), .QN(n3117) );
  INVX0 U2633 ( .IN(n3120), .QN(n3131) );
  INVX0 U2634 ( .IN(n3120), .QN(n3130) );
  INVX0 U2635 ( .IN(n3139), .QN(n3132) );
  INVX0 U2636 ( .IN(n3137), .QN(n3134) );
  INVX0 U2637 ( .IN(n3158), .QN(n3169) );
  INVX0 U2638 ( .IN(n3160), .QN(n3175) );
  INVX0 U2639 ( .IN(n3158), .QN(n3174) );
  INVX0 U2640 ( .IN(n3160), .QN(n3179) );
  INVX0 U2641 ( .IN(n3157), .QN(n3171) );
  INVX0 U2642 ( .IN(n3160), .QN(n3178) );
  INVX0 U2643 ( .IN(n3157), .QN(n3172) );
  INVX0 U2644 ( .IN(n3159), .QN(n3177) );
  INVX0 U2645 ( .IN(n3158), .QN(n3173) );
  INVX0 U2646 ( .IN(n3159), .QN(n3176) );
  AND4X1 U2647 ( .IN1(n4113), .IN2(n3104), .IN3(n4811), .IN4(n3185), .Q(n2950)
         );
  NBUFFX2 U2648 ( .IN(n4060), .Q(n3232) );
  NBUFFX2 U2649 ( .IN(n4060), .Q(n3231) );
  NBUFFX2 U2650 ( .IN(n4060), .Q(n3233) );
  NBUFFX2 U2651 ( .IN(n4060), .Q(n3234) );
  NBUFFX2 U2652 ( .IN(n4060), .Q(n3235) );
  NBUFFX2 U2653 ( .IN(n4060), .Q(n3236) );
  NBUFFX2 U2654 ( .IN(n3336), .Q(n3324) );
  NBUFFX2 U2655 ( .IN(n4076), .Q(n3336) );
  NBUFFX2 U2656 ( .IN(n3249), .Q(n3239) );
  NBUFFX2 U2657 ( .IN(n3248), .Q(n3240) );
  NBUFFX2 U2658 ( .IN(n3249), .Q(n3238) );
  NBUFFX2 U2659 ( .IN(n3247), .Q(n3242) );
  NBUFFX2 U2660 ( .IN(n3247), .Q(n3243) );
  NBUFFX2 U2661 ( .IN(n3246), .Q(n3244) );
  NBUFFX2 U2662 ( .IN(n3246), .Q(n3245) );
  NBUFFX2 U2663 ( .IN(n4076), .Q(n3332) );
  NBUFFX2 U2664 ( .IN(n4076), .Q(n3335) );
  NBUFFX2 U2665 ( .IN(n4076), .Q(n3334) );
  NBUFFX2 U2666 ( .IN(n4076), .Q(n3333) );
  NBUFFX2 U2667 ( .IN(n4070), .Q(n3273) );
  NBUFFX2 U2668 ( .IN(n4070), .Q(n3274) );
  NBUFFX2 U2669 ( .IN(n4070), .Q(n3272) );
  NBUFFX2 U2670 ( .IN(n4070), .Q(n3275) );
  NBUFFX2 U2671 ( .IN(n4830), .Q(n3451) );
  NBUFFX2 U2672 ( .IN(n4830), .Q(n3452) );
  NBUFFX2 U2673 ( .IN(n4060), .Q(n3237) );
  NBUFFX2 U2674 ( .IN(n4072), .Q(n3285) );
  NBUFFX2 U2675 ( .IN(n4073), .Q(n3297) );
  NBUFFX2 U2676 ( .IN(n4074), .Q(n3309) );
  NBUFFX2 U2677 ( .IN(n4075), .Q(n3321) );
  NBUFFX2 U2678 ( .IN(n4072), .Q(n3286) );
  NBUFFX2 U2679 ( .IN(n4073), .Q(n3298) );
  NBUFFX2 U2680 ( .IN(n4074), .Q(n3310) );
  NBUFFX2 U2681 ( .IN(n4075), .Q(n3322) );
  NBUFFX2 U2682 ( .IN(n4072), .Q(n3284) );
  NBUFFX2 U2683 ( .IN(n4073), .Q(n3296) );
  NBUFFX2 U2684 ( .IN(n4074), .Q(n3308) );
  NBUFFX2 U2685 ( .IN(n4075), .Q(n3320) );
  NBUFFX2 U2686 ( .IN(n4072), .Q(n3287) );
  NBUFFX2 U2687 ( .IN(n4073), .Q(n3299) );
  NBUFFX2 U2688 ( .IN(n4074), .Q(n3311) );
  NBUFFX2 U2689 ( .IN(n4075), .Q(n3323) );
  AND4X1 U2690 ( .IN1(n4113), .IN2(n3104), .IN3(n4811), .IN4(n3185), .Q(n2951)
         );
  AND4X1 U2691 ( .IN1(n4113), .IN2(n3104), .IN3(n4811), .IN4(n3185), .Q(n2952)
         );
  NBUFFX2 U2692 ( .IN(n4825), .Q(n3413) );
  NBUFFX2 U2693 ( .IN(n4825), .Q(n3412) );
  NBUFFX2 U2694 ( .IN(n4825), .Q(n3411) );
  NBUFFX2 U2695 ( .IN(n4825), .Q(n3414) );
  NBUFFX2 U2696 ( .IN(n4825), .Q(n3416) );
  NBUFFX2 U2697 ( .IN(n4825), .Q(n3415) );
  NBUFFX2 U2698 ( .IN(n4827), .Q(n3429) );
  NBUFFX2 U2699 ( .IN(n4827), .Q(n3428) );
  NBUFFX2 U2700 ( .IN(n4827), .Q(n3427) );
  NBUFFX2 U2701 ( .IN(n4827), .Q(n3426) );
  NBUFFX2 U2702 ( .IN(n4827), .Q(n3425) );
  NBUFFX2 U2703 ( .IN(n4827), .Q(n3424) );
  NBUFFX2 U2704 ( .IN(n5203), .Q(n3525) );
  NBUFFX2 U2705 ( .IN(n5203), .Q(n3526) );
  NBUFFX2 U2706 ( .IN(n5203), .Q(n3527) );
  NBUFFX2 U2707 ( .IN(n5203), .Q(n3528) );
  NBUFFX2 U2708 ( .IN(n5203), .Q(n3529) );
  NBUFFX2 U2709 ( .IN(n5203), .Q(n3530) );
  NBUFFX2 U2710 ( .IN(n3538), .Q(n3537) );
  NBUFFX2 U2711 ( .IN(n3539), .Q(n3536) );
  NBUFFX2 U2712 ( .IN(n3539), .Q(n3535) );
  NBUFFX2 U2713 ( .IN(n3540), .Q(n3534) );
  NBUFFX2 U2714 ( .IN(n3540), .Q(n3533) );
  NBUFFX2 U2715 ( .IN(n3376), .Q(n3367) );
  NBUFFX2 U2716 ( .IN(n4119), .Q(n3376) );
  NBUFFX2 U2717 ( .IN(n3366), .Q(n3356) );
  NBUFFX2 U2718 ( .IN(n4118), .Q(n3366) );
  NBUFFX2 U2719 ( .IN(n3498), .Q(n3496) );
  NBUFFX2 U2720 ( .IN(n3499), .Q(n3495) );
  NBUFFX2 U2721 ( .IN(n3499), .Q(n3494) );
  NBUFFX2 U2722 ( .IN(n3500), .Q(n3493) );
  NBUFFX2 U2723 ( .IN(n3500), .Q(n3492) );
  NBUFFX2 U2724 ( .IN(n3501), .Q(n3490) );
  NBUFFX2 U2725 ( .IN(n3501), .Q(n3491) );
  NBUFFX2 U2726 ( .IN(n3498), .Q(n3497) );
  NBUFFX2 U2727 ( .IN(n3248), .Q(n3241) );
  NBUFFX2 U2728 ( .IN(n5074), .Q(n3522) );
  NBUFFX2 U2729 ( .IN(n5074), .Q(n3521) );
  NBUFFX2 U2730 ( .IN(n5074), .Q(n3523) );
  NBUFFX2 U2731 ( .IN(n4118), .Q(n3365) );
  NBUFFX2 U2732 ( .IN(n4118), .Q(n3364) );
  NBUFFX2 U2733 ( .IN(n4118), .Q(n3363) );
  NBUFFX2 U2734 ( .IN(n4119), .Q(n3373) );
  NBUFFX2 U2735 ( .IN(n4119), .Q(n3374) );
  NBUFFX2 U2736 ( .IN(n4119), .Q(n3375) );
  NBUFFX2 U2737 ( .IN(n5203), .Q(n3531) );
  NBUFFX2 U2738 ( .IN(n4827), .Q(n3430) );
  NBUFFX2 U2739 ( .IN(n5073), .Q(n3511) );
  NBUFFX2 U2740 ( .IN(n5073), .Q(n3512) );
  NBUFFX2 U2741 ( .IN(n5073), .Q(n3513) );
  NBUFFX2 U2742 ( .IN(n5073), .Q(n3510) );
  NBUFFX2 U2743 ( .IN(n5071), .Q(n3487) );
  NBUFFX2 U2744 ( .IN(n5071), .Q(n3488) );
  NBUFFX2 U2745 ( .IN(n5071), .Q(n3489) );
  NBUFFX2 U2746 ( .IN(n5071), .Q(n3486) );
  NBUFFX2 U2747 ( .IN(n3524), .Q(n3514) );
  NBUFFX2 U2748 ( .IN(n5074), .Q(n3524) );
  INVX0 U2749 ( .IN(n4103), .QN(n4012) );
  INVX0 U2750 ( .IN(n4181), .QN(n4221) );
  INVX0 U2751 ( .IN(n4164), .QN(n3393) );
  INVX0 U2752 ( .IN(n3389), .QN(n3395) );
  INVX0 U2753 ( .IN(n3389), .QN(n3394) );
  INVX0 U2754 ( .IN(n4164), .QN(n3396) );
  INVX0 U2755 ( .IN(n4015), .QN(n3184) );
  NBUFFX2 U2756 ( .IN(n3385), .Q(n3383) );
  NBUFFX2 U2757 ( .IN(n3388), .Q(n3384) );
  INVX0 U2758 ( .IN(n3392), .QN(n3397) );
  INVX0 U2759 ( .IN(n3392), .QN(n3398) );
  NBUFFX2 U2760 ( .IN(n3387), .Q(n3378) );
  NBUFFX2 U2761 ( .IN(n3387), .Q(n3379) );
  NBUFFX2 U2762 ( .IN(n3386), .Q(n3380) );
  NBUFFX2 U2763 ( .IN(n3386), .Q(n3381) );
  NBUFFX2 U2764 ( .IN(n3385), .Q(n3382) );
  NBUFFX2 U2765 ( .IN(n4111), .Q(n3345) );
  NBUFFX2 U2766 ( .IN(n4111), .Q(n3348) );
  NBUFFX2 U2767 ( .IN(n4111), .Q(n3347) );
  NBUFFX2 U2768 ( .IN(n4111), .Q(n3346) );
  NBUFFX2 U2769 ( .IN(n3612), .Q(n3610) );
  NBUFFX2 U2770 ( .IN(n3612), .Q(n3611) );
  NBUFFX2 U2771 ( .IN(n3673), .Q(n3647) );
  NBUFFX2 U2772 ( .IN(n3673), .Q(n3648) );
  NBUFFX2 U2773 ( .IN(n3672), .Q(n3649) );
  NBUFFX2 U2774 ( .IN(n3672), .Q(n3650) );
  NBUFFX2 U2775 ( .IN(n3671), .Q(n3651) );
  NBUFFX2 U2776 ( .IN(n3671), .Q(n3652) );
  NBUFFX2 U2777 ( .IN(n3670), .Q(n3653) );
  NBUFFX2 U2778 ( .IN(n3670), .Q(n3654) );
  NBUFFX2 U2779 ( .IN(n3669), .Q(n3655) );
  NBUFFX2 U2780 ( .IN(n3669), .Q(n3656) );
  NBUFFX2 U2781 ( .IN(n3668), .Q(n3657) );
  NBUFFX2 U2782 ( .IN(n3668), .Q(n3658) );
  NBUFFX2 U2783 ( .IN(n3667), .Q(n3659) );
  NBUFFX2 U2784 ( .IN(n3667), .Q(n3660) );
  NBUFFX2 U2785 ( .IN(n3666), .Q(n3661) );
  NBUFFX2 U2786 ( .IN(n3666), .Q(n3662) );
  NBUFFX2 U2787 ( .IN(n3663), .Q(n3614) );
  NBUFFX2 U2788 ( .IN(n3663), .Q(n3613) );
  INVX0 U2789 ( .IN(n3893), .QN(n3112) );
  INVX0 U2790 ( .IN(n3170), .QN(n3161) );
  INVX0 U2791 ( .IN(n3125), .QN(n3119) );
  INVX0 U2792 ( .IN(n3896), .QN(n3138) );
  INVX0 U2793 ( .IN(n3896), .QN(n3136) );
  INVX0 U2794 ( .IN(n3896), .QN(n3139) );
  NBUFFX2 U2795 ( .IN(n2953), .Q(n3680) );
  INVX0 U2796 ( .IN(n3889), .QN(n3881) );
  INVX0 U2797 ( .IN(n3163), .QN(n3158) );
  INVX0 U2798 ( .IN(n3162), .QN(n3160) );
  INVX0 U2799 ( .IN(n3163), .QN(n3157) );
  INVX0 U2800 ( .IN(n3125), .QN(n3120) );
  INVX0 U2801 ( .IN(n3113), .QN(n3106) );
  INVX0 U2802 ( .IN(n3162), .QN(n3159) );
  INVX0 U2803 ( .IN(n3896), .QN(n3137) );
  NBUFFX2 U2804 ( .IN(n2953), .Q(n3679) );
  INVX0 U2805 ( .IN(n4021), .QN(mult_add_463_aco_A_0_) );
  NOR3X0 U2806 ( .IN1(N3423), .IN2(N3427), .IN3(N3424), .QN(n3689) );
  INVX0 U2807 ( .IN(N3417), .QN(N3424) );
  INVX0 U2808 ( .IN(N3418), .QN(N3423) );
  NBUFFX2 U2809 ( .IN(n2953), .Q(n3681) );
  NBUFFX2 U2810 ( .IN(n4068), .Q(n3262) );
  NBUFFX2 U2811 ( .IN(n4068), .Q(n3261) );
  NBUFFX2 U2812 ( .IN(n4068), .Q(n3260) );
  NBUFFX2 U2813 ( .IN(n4068), .Q(n3259) );
  NBUFFX2 U2814 ( .IN(n4068), .Q(n3257) );
  NBUFFX2 U2815 ( .IN(n4068), .Q(n3258) );
  NBUFFX2 U2816 ( .IN(n4828), .Q(n3437) );
  NBUFFX2 U2817 ( .IN(n4068), .Q(n3263) );
  NBUFFX2 U2818 ( .IN(n4062), .Q(n3248) );
  NBUFFX2 U2819 ( .IN(n4062), .Q(n3247) );
  NBUFFX2 U2820 ( .IN(n4062), .Q(n3246) );
  NBUFFX2 U2821 ( .IN(n4062), .Q(n3249) );
  NBUFFX2 U2822 ( .IN(n4826), .Q(n3419) );
  NBUFFX2 U2823 ( .IN(n4826), .Q(n3418) );
  NBUFFX2 U2824 ( .IN(n4826), .Q(n3417) );
  NBUFFX2 U2825 ( .IN(n4058), .Q(n3219) );
  NBUFFX2 U2826 ( .IN(n4058), .Q(n3218) );
  NBUFFX2 U2827 ( .IN(n4826), .Q(n3420) );
  NBUFFX2 U2828 ( .IN(n4826), .Q(n3422) );
  NBUFFX2 U2829 ( .IN(n4826), .Q(n3421) );
  NBUFFX2 U2830 ( .IN(n4117), .Q(n3349) );
  NBUFFX2 U2831 ( .IN(n3440), .Q(n3432) );
  NBUFFX2 U2832 ( .IN(n3439), .Q(n3433) );
  NBUFFX2 U2833 ( .IN(n3438), .Q(n3435) );
  NBUFFX2 U2834 ( .IN(n3438), .Q(n3436) );
  NBUFFX2 U2835 ( .IN(n3439), .Q(n3434) );
  NBUFFX2 U2836 ( .IN(n3440), .Q(n3431) );
  NBUFFX2 U2837 ( .IN(n4058), .Q(n3220) );
  NBUFFX2 U2838 ( .IN(n4058), .Q(n3221) );
  NBUFFX2 U2839 ( .IN(n4058), .Q(n3222) );
  NBUFFX2 U2840 ( .IN(n4058), .Q(n3223) );
  NBUFFX2 U2841 ( .IN(n4117), .Q(n3355) );
  NBUFFX2 U2842 ( .IN(n4826), .Q(n3423) );
  NBUFFX2 U2843 ( .IN(n5204), .Q(n3538) );
  NBUFFX2 U2844 ( .IN(n5204), .Q(n3539) );
  NBUFFX2 U2845 ( .IN(n5204), .Q(n3540) );
  NBUFFX2 U2846 ( .IN(n5072), .Q(n3499) );
  NBUFFX2 U2847 ( .IN(n5072), .Q(n3500) );
  NBUFFX2 U2848 ( .IN(n5072), .Q(n3501) );
  NBUFFX2 U2849 ( .IN(n5072), .Q(n3498) );
  NBUFFX2 U2850 ( .IN(n4058), .Q(n3224) );
  NBUFFX2 U2851 ( .IN(n3541), .Q(n3532) );
  NBUFFX2 U2852 ( .IN(n5204), .Q(n3541) );
  NOR2X0 U2853 ( .IN1(n4594), .IN2(n3396), .QN(n4568) );
  NOR2X0 U2854 ( .IN1(n4617), .IN2(n3394), .QN(n4599) );
  NOR2X0 U2855 ( .IN1(n4255), .IN2(n3393), .QN(n4227) );
  NOR2X0 U2856 ( .IN1(n4620), .IN2(n3394), .QN(n4623) );
  INVX0 U2857 ( .IN(n4594), .QN(n4530) );
  INVX0 U2858 ( .IN(n4255), .QN(n4222) );
  INVX0 U2859 ( .IN(n3396), .QN(n3389) );
  NBUFFX2 U2860 ( .IN(n4117), .Q(n3350) );
  NBUFFX2 U2861 ( .IN(n4117), .Q(n3351) );
  NBUFFX2 U2862 ( .IN(n4117), .Q(n3352) );
  NBUFFX2 U2863 ( .IN(n4117), .Q(n3353) );
  NBUFFX2 U2864 ( .IN(n4117), .Q(n3354) );
  NBUFFX2 U2865 ( .IN(n4156), .Q(n3385) );
  INVX0 U2866 ( .IN(n4620), .QN(n4186) );
  INVX0 U2867 ( .IN(n4617), .QN(n4563) );
  INVX0 U2868 ( .IN(n2956), .QN(n3104) );
  INVX0 U2869 ( .IN(n2956), .QN(n3105) );
  NBUFFX2 U2870 ( .IN(n4024), .Q(n3205) );
  NBUFFX2 U2871 ( .IN(n4024), .Q(n3206) );
  NBUFFX2 U2872 ( .IN(n4024), .Q(n3207) );
  NBUFFX2 U2873 ( .IN(n4024), .Q(n3209) );
  NBUFFX2 U2874 ( .IN(n4024), .Q(n3208) );
  NBUFFX2 U2875 ( .IN(n4024), .Q(n3210) );
  NBUFFX2 U2876 ( .IN(n4813), .Q(n3404) );
  NBUFFX2 U2877 ( .IN(n4813), .Q(n3403) );
  NBUFFX2 U2878 ( .IN(n4813), .Q(n3402) );
  NBUFFX2 U2879 ( .IN(n4813), .Q(n3401) );
  NBUFFX2 U2880 ( .IN(n4813), .Q(n3400) );
  NBUFFX2 U2881 ( .IN(n4813), .Q(n3399) );
  NBUFFX2 U2882 ( .IN(n4049), .Q(n3212) );
  NBUFFX2 U2883 ( .IN(n4049), .Q(n3217) );
  NBUFFX2 U2884 ( .IN(n4049), .Q(n3216) );
  NBUFFX2 U2885 ( .IN(n4049), .Q(n3215) );
  NBUFFX2 U2886 ( .IN(n4049), .Q(n3214) );
  NBUFFX2 U2887 ( .IN(n4049), .Q(n3213) );
  NBUFFX2 U2888 ( .IN(n4024), .Q(n3211) );
  NBUFFX2 U2889 ( .IN(n4156), .Q(n3387) );
  NBUFFX2 U2890 ( .IN(n4156), .Q(n3386) );
  NBUFFX2 U2891 ( .IN(n3388), .Q(n3377) );
  NBUFFX2 U2892 ( .IN(n4156), .Q(n3388) );
  NBUFFX2 U2893 ( .IN(n3674), .Q(n3673) );
  NBUFFX2 U2894 ( .IN(n3674), .Q(n3672) );
  NBUFFX2 U2895 ( .IN(n3675), .Q(n3671) );
  NBUFFX2 U2896 ( .IN(n3675), .Q(n3670) );
  NBUFFX2 U2897 ( .IN(n3676), .Q(n3669) );
  NBUFFX2 U2898 ( .IN(n3676), .Q(n3668) );
  NBUFFX2 U2899 ( .IN(n3677), .Q(n3667) );
  NBUFFX2 U2900 ( .IN(n3677), .Q(n3666) );
  NBUFFX2 U2901 ( .IN(n3665), .Q(n3663) );
  NBUFFX2 U2902 ( .IN(n3664), .Q(n3612) );
  NBUFFX2 U2903 ( .IN(n3665), .Q(n3664) );
  NAND2X0 U2904 ( .IN1(add_2_root_sub_1_root_sub_357_2_carry[7]), .IN2(N2392), 
        .QN(n2953) );
  NAND2X0 U2905 ( .IN1(N2737), .IN2(InstQueueRd_Addr[1]), .QN(n3889) );
  INVX0 U2906 ( .IN(n3887), .QN(n3884) );
  INVX0 U2907 ( .IN(n3897), .QN(n3163) );
  INVX0 U2908 ( .IN(n3897), .QN(n3162) );
  NBUFFX2 U2909 ( .IN(n4059), .Q(n3227) );
  NBUFFX2 U2910 ( .IN(n4059), .Q(n3226) );
  NBUFFX2 U2911 ( .IN(n4059), .Q(n3225) );
  NBUFFX2 U2912 ( .IN(n4063), .Q(n3251) );
  NBUFFX2 U2913 ( .IN(n4063), .Q(n3252) );
  NBUFFX2 U2914 ( .IN(n4063), .Q(n3253) );
  NBUFFX2 U2915 ( .IN(n4059), .Q(n3230) );
  NOR2X0 U2916 ( .IN1(n2954), .IN2(n4091), .QN(n5060) );
  INVX0 U2917 ( .IN(n3332), .QN(n2954) );
  NAND2X0 U2918 ( .IN1(r679_carry[4]), .IN2(n3871), .QN(n2955) );
  NBUFFX2 U2919 ( .IN(n4059), .Q(n3228) );
  NBUFFX2 U2920 ( .IN(n4059), .Q(n3229) );
  NBUFFX2 U2921 ( .IN(n4063), .Q(n3250) );
  NBUFFX2 U2922 ( .IN(n4063), .Q(n3254) );
  NBUFFX2 U2923 ( .IN(n4063), .Q(n3255) );
  NBUFFX2 U2924 ( .IN(n4828), .Q(n3438) );
  NBUFFX2 U2925 ( .IN(n4828), .Q(n3439) );
  NBUFFX2 U2926 ( .IN(n4828), .Q(n3440) );
  NBUFFX2 U2927 ( .IN(n4063), .Q(n3256) );
  AO22X1 U2928 ( .IN1(Datai[1]), .IN2(n3384), .IN3(n4089), .IN4(n4628), .Q(
        n4193) );
  AO22X1 U2929 ( .IN1(Datai[2]), .IN2(n3384), .IN3(n4089), .IN4(n4631), .Q(
        n4197) );
  AO22X1 U2930 ( .IN1(Datai[0]), .IN2(n3384), .IN3(n4089), .IN4(n4126), .Q(
        n4188) );
  AO22X1 U2931 ( .IN1(n3086), .IN2(n3384), .IN3(n4089), .IN4(n4635), .Q(n4201)
         );
  AO22X1 U2932 ( .IN1(n3088), .IN2(n3384), .IN3(n4089), .IN4(n4638), .Q(n4205)
         );
  AO22X1 U2933 ( .IN1(Datai[5]), .IN2(n3383), .IN3(n4089), .IN4(n4641), .Q(
        n4210) );
  AO22X1 U2934 ( .IN1(Datai[6]), .IN2(n3383), .IN3(n4089), .IN4(n4644), .Q(
        n4214) );
  AO22X1 U2935 ( .IN1(Datai[7]), .IN2(n3383), .IN3(n4089), .IN4(n4647), .Q(
        n4218) );
  NOR2X0 U2936 ( .IN1(n4370), .IN2(n3393), .QN(n4343) );
  NOR2X0 U2937 ( .IN1(n4562), .IN2(n3395), .QN(n4535) );
  NOR2X0 U2938 ( .IN1(n4303), .IN2(n3393), .QN(n4261) );
  NOR2X0 U2939 ( .IN1(n4256), .IN2(n3393), .QN(n4183) );
  NOR2X0 U2940 ( .IN1(n4417), .IN2(n3393), .QN(n4376) );
  NOR2X0 U2941 ( .IN1(n4418), .IN2(n3393), .QN(n4399) );
  NOR2X0 U2942 ( .IN1(n4369), .IN2(n3393), .QN(n4311) );
  NOR2X0 U2943 ( .IN1(n4304), .IN2(n3395), .QN(n4285) );
  NOR2X0 U2944 ( .IN1(n4482), .IN2(n3395), .QN(n4424) );
  NOR2X0 U2945 ( .IN1(n4561), .IN2(n3395), .QN(n4512) );
  NOR2X0 U2946 ( .IN1(n4506), .IN2(n3394), .QN(n4488) );
  INVX0 U2947 ( .IN(n4370), .QN(n4305) );
  INVX0 U2948 ( .IN(n4369), .QN(n4280) );
  INVX0 U2949 ( .IN(n4482), .QN(n4394) );
  INVX0 U2950 ( .IN(n4173), .QN(n4419) );
  INVX0 U2951 ( .IN(n3996), .QN(n3877) );
  INVX0 U2952 ( .IN(n4562), .QN(n4507) );
  INVX0 U2953 ( .IN(n3998), .QN(n3875) );
  INVX0 U2954 ( .IN(n4091), .QN(n4017) );
  INVX0 U2955 ( .IN(n4174), .QN(n4254) );
  INVX0 U2956 ( .IN(n3089), .QN(n3090) );
  INVX0 U2957 ( .IN(n3081), .QN(n3082) );
  INVX0 U2958 ( .IN(n3093), .QN(n3094) );
  INVX0 U2959 ( .IN(n3083), .QN(n3084) );
  INVX0 U2960 ( .IN(n3091), .QN(n3092) );
  INVX0 U2961 ( .IN(n3079), .QN(n3080) );
  INVX0 U2962 ( .IN(n3087), .QN(n3088) );
  INVX0 U2963 ( .IN(n3085), .QN(n3086) );
  NOR2X0 U2964 ( .IN1(n2948), .IN2(n2868), .QN(n5309) );
  INVX0 U2965 ( .IN(n4095), .QN(n4089) );
  INVX0 U2966 ( .IN(n4417), .QN(n4337) );
  INVX0 U2967 ( .IN(n4418), .QN(n4371) );
  INVX0 U2968 ( .IN(n4303), .QN(n4220) );
  INVX0 U2969 ( .IN(n4304), .QN(n4257) );
  INVX0 U2970 ( .IN(n4561), .QN(n4483) );
  INVX0 U2971 ( .IN(n4506), .QN(n4450) );
  INVX0 U2972 ( .IN(n4256), .QN(n4219) );
  AND3X1 U2973 ( .IN1(n2842), .IN2(n4097), .IN3(n4649), .Q(n2956) );
  OAI21X1 U2974 ( .IN1(N3485), .IN2(N3486), .IN3(N3484), .QN(n3690) );
  NBUFFX2 U2975 ( .IN(n5315), .Q(n3674) );
  NBUFFX2 U2976 ( .IN(n5315), .Q(n3675) );
  NBUFFX2 U2977 ( .IN(n5315), .Q(n3676) );
  NBUFFX2 U2978 ( .IN(n5315), .Q(n3677) );
  NBUFFX2 U2979 ( .IN(n3678), .Q(n3665) );
  NBUFFX2 U2980 ( .IN(n5315), .Q(n3678) );
  INVX0 U2981 ( .IN(N2386), .QN(n5316) );
  NAND2X0 U2982 ( .IN1(n1550), .IN2(N2737), .QN(n3887) );
  INVX0 U2983 ( .IN(N3419), .QN(n3688) );
  NAND2X0 U2984 ( .IN1(n1552), .IN2(InstQueueRd_Addr[1]), .QN(n3996) );
  NAND2X0 U2985 ( .IN1(n1550), .IN2(n1552), .QN(n3998) );
  AND2X1 U2986 ( .IN1(N1763), .IN2(mult_add_463_aco_A_0_), .Q(n2957) );
  AND2X1 U2987 ( .IN1(N1762), .IN2(mult_add_463_aco_A_0_), .Q(n2958) );
  AND2X1 U2988 ( .IN1(N1761), .IN2(mult_add_463_aco_A_0_), .Q(n2959) );
  AND2X1 U2989 ( .IN1(N1760), .IN2(mult_add_463_aco_A_0_), .Q(n2960) );
  AND2X1 U2990 ( .IN1(N1759), .IN2(mult_add_463_aco_A_0_), .Q(n2961) );
  AND2X1 U2991 ( .IN1(N1758), .IN2(mult_add_463_aco_A_0_), .Q(n2962) );
  AND2X1 U2992 ( .IN1(N1757), .IN2(mult_add_463_aco_A_0_), .Q(n2963) );
  AND2X1 U2993 ( .IN1(N1756), .IN2(mult_add_463_aco_A_0_), .Q(n2964) );
  AND2X1 U2994 ( .IN1(N1755), .IN2(mult_add_463_aco_A_0_), .Q(n2965) );
  AND2X1 U2995 ( .IN1(N1754), .IN2(mult_add_463_aco_A_0_), .Q(n2966) );
  AND2X1 U2996 ( .IN1(N1753), .IN2(mult_add_463_aco_A_0_), .Q(n2967) );
  AND2X1 U2997 ( .IN1(N1752), .IN2(mult_add_463_aco_A_0_), .Q(n2968) );
  AND2X1 U2998 ( .IN1(N1751), .IN2(mult_add_463_aco_A_0_), .Q(n2969) );
  AND2X1 U2999 ( .IN1(N1750), .IN2(mult_add_463_aco_A_0_), .Q(n2970) );
  FADDX1 U3000 ( .A(N3989), .B(n1548), .CI(r679_carry[3]), .CO(r679_carry[4]), 
        .S(r680_B_3_) );
  FADDX1 U3001 ( .A(N3991), .B(n1550), .CI(r679_carry[1]), .CO(r679_carry[2]), 
        .S(r680_B_1_) );
  FADDX1 U3002 ( .A(N3990), .B(n3839), .CI(r679_carry[2]), .CO(r679_carry[3]), 
        .S(r680_B_2_) );
  NAND3X0 U3003 ( .IN1(n5200), .IN2(n2844), .IN3(n1490), .QN(n4174) );
  NAND3X0 U3004 ( .IN1(n1491), .IN2(n2865), .IN3(n4116), .QN(n4091) );
  NOR2X0 U3005 ( .IN1(n2971), .IN2(n3398), .QN(n4216) );
  XNOR2X1 U3006 ( .IN1(Datai[31]), .IN2(add_div_313_carry[7]), .Q(n2971) );
  NBUFFX2 U3007 ( .IN(N655), .Q(n3097) );
  NBUFFX2 U3008 ( .IN(N656), .Q(n3096) );
  NBUFFX2 U3009 ( .IN(N657), .Q(n3095) );
  NOR2X0 U3010 ( .IN1(n2972), .IN2(n3398), .QN(n4203) );
  XNOR2X1 U3011 ( .IN1(Datai[28]), .IN2(add_div_313_carry[4]), .Q(n2972) );
  NOR2X0 U3012 ( .IN1(n2973), .IN2(n3397), .QN(n4208) );
  XNOR2X1 U3013 ( .IN1(Datai[29]), .IN2(add_div_313_carry[5]), .Q(n2973) );
  NOR2X0 U3014 ( .IN1(n2974), .IN2(n3397), .QN(n4212) );
  XNOR2X1 U3015 ( .IN1(Datai[30]), .IN2(add_div_313_carry[6]), .Q(n2974) );
  NAND2X0 U3016 ( .IN1(add_div_311_carry[6]), .IN2(Datai[22]), .QN(n2975) );
  INVX0 U3017 ( .IN(Datai[7]), .QN(n3093) );
  INVX0 U3018 ( .IN(Datai[6]), .QN(n3091) );
  INVX0 U3019 ( .IN(Datai[5]), .QN(n3089) );
  INVX0 U3020 ( .IN(Datai[4]), .QN(n3087) );
  INVX0 U3021 ( .IN(Datai[3]), .QN(n3085) );
  INVX0 U3022 ( .IN(Datai[2]), .QN(n3083) );
  INVX0 U3023 ( .IN(Datai[1]), .QN(n3081) );
  INVX0 U3024 ( .IN(Datai[0]), .QN(n3079) );
  NOR2X0 U3025 ( .IN1(n2976), .IN2(n3398), .QN(n4185) );
  XNOR2X1 U3026 ( .IN1(Datai[24]), .IN2(N811), .Q(n2976) );
  NOR2X0 U3027 ( .IN1(n2977), .IN2(n3397), .QN(n4191) );
  XNOR2X1 U3028 ( .IN1(Datai[25]), .IN2(add_div_313_carry[1]), .Q(n2977) );
  NOR2X0 U3029 ( .IN1(n2978), .IN2(n3398), .QN(n4195) );
  XNOR2X1 U3030 ( .IN1(Datai[26]), .IN2(add_div_313_carry[2]), .Q(n2978) );
  NOR2X0 U3031 ( .IN1(n2979), .IN2(n3397), .QN(n4199) );
  XNOR2X1 U3032 ( .IN1(Datai[27]), .IN2(add_div_313_carry[3]), .Q(n2979) );
  NOR3X0 U3033 ( .IN1(N3493), .IN2(n3690), .IN3(n2887), .QN(n3691) );
  HADDX1 U3034 ( .A0(InstQueueRd_Addr[1]), .B0(N2737), .C1(r698_carry[2]), 
        .SO(N2700) );
  HADDX1 U3035 ( .A0(InstQueueRd_Addr[3]), .B0(r698_carry[3]), .C1(
        r698_carry[4]), .SO(N2702) );
  HADDX1 U3036 ( .A0(InstQueueRd_Addr[2]), .B0(r698_carry[2]), .C1(
        r698_carry[3]), .SO(N2701) );
  NBUFFX2 U3037 ( .IN(N651), .Q(n3101) );
  NBUFFX2 U3038 ( .IN(N652), .Q(n3100) );
  NBUFFX2 U3039 ( .IN(N653), .Q(n3099) );
  NBUFFX2 U3040 ( .IN(N654), .Q(n3098) );
  HADDX1 U3041 ( .A0(InstQueueRd_Addr[4]), .B0(r698_carry[4]), .C1(N2704), 
        .SO(N2703) );
  XOR2X1 U3042 ( .IN1(Datai[22]), .IN2(add_div_311_carry[6]), .Q(N657) );
  AND2X1 U3043 ( .IN1(add_div_311_carry[5]), .IN2(Datai[21]), .Q(
        add_div_311_carry[6]) );
  XOR2X1 U3044 ( .IN1(Datai[21]), .IN2(add_div_311_carry[5]), .Q(N656) );
  AND2X1 U3045 ( .IN1(add_div_311_carry[4]), .IN2(Datai[20]), .Q(
        add_div_311_carry[5]) );
  XOR2X1 U3046 ( .IN1(Datai[20]), .IN2(add_div_311_carry[4]), .Q(N655) );
  AND2X1 U3047 ( .IN1(add_div_311_carry[3]), .IN2(Datai[19]), .Q(
        add_div_311_carry[4]) );
  XOR2X1 U3048 ( .IN1(Datai[19]), .IN2(add_div_311_carry[3]), .Q(N654) );
  AND2X1 U3049 ( .IN1(add_div_311_carry[2]), .IN2(Datai[18]), .Q(
        add_div_311_carry[3]) );
  XOR2X1 U3050 ( .IN1(Datai[18]), .IN2(add_div_311_carry[2]), .Q(N653) );
  AND2X1 U3051 ( .IN1(add_div_311_carry[1]), .IN2(Datai[17]), .Q(
        add_div_311_carry[2]) );
  XOR2X1 U3052 ( .IN1(Datai[17]), .IN2(add_div_311_carry[1]), .Q(N652) );
  AND2X1 U3053 ( .IN1(add_div_311_A_0_), .IN2(Datai[16]), .Q(
        add_div_311_carry[1]) );
  XOR2X1 U3054 ( .IN1(Datai[16]), .IN2(add_div_311_A_0_), .Q(N651) );
  AND2X1 U3055 ( .IN1(add_div_313_carry[6]), .IN2(Datai[30]), .Q(
        add_div_313_carry[7]) );
  AND2X1 U3056 ( .IN1(add_div_313_carry[5]), .IN2(Datai[29]), .Q(
        add_div_313_carry[6]) );
  AND2X1 U3057 ( .IN1(add_div_313_carry[4]), .IN2(Datai[28]), .Q(
        add_div_313_carry[5]) );
  AND2X1 U3058 ( .IN1(add_div_313_carry[3]), .IN2(Datai[27]), .Q(
        add_div_313_carry[4]) );
  AND2X1 U3059 ( .IN1(add_div_313_carry[2]), .IN2(Datai[26]), .Q(
        add_div_313_carry[3]) );
  AND2X1 U3060 ( .IN1(add_div_313_carry[1]), .IN2(Datai[25]), .Q(
        add_div_313_carry[2]) );
  AND2X1 U3061 ( .IN1(N811), .IN2(Datai[24]), .Q(add_div_313_carry[1]) );
  XOR2X1 U3062 ( .IN1(test_so5), .IN2(add_div_457_carry[14]), .Q(N1764) );
  AND2X1 U3063 ( .IN1(add_div_457_carry[13]), .IN2(EAX_29_), .Q(
        add_div_457_carry[14]) );
  XOR2X1 U3064 ( .IN1(EAX_29_), .IN2(add_div_457_carry[13]), .Q(N1763) );
  AND2X1 U3065 ( .IN1(add_div_457_carry[12]), .IN2(EAX_28_), .Q(
        add_div_457_carry[13]) );
  XOR2X1 U3066 ( .IN1(EAX_28_), .IN2(add_div_457_carry[12]), .Q(N1762) );
  AND2X1 U3067 ( .IN1(add_div_457_carry[11]), .IN2(EAX_27_), .Q(
        add_div_457_carry[12]) );
  XOR2X1 U3068 ( .IN1(EAX_27_), .IN2(add_div_457_carry[11]), .Q(N1761) );
  AND2X1 U3069 ( .IN1(add_div_457_carry[10]), .IN2(EAX_26_), .Q(
        add_div_457_carry[11]) );
  XOR2X1 U3070 ( .IN1(EAX_26_), .IN2(add_div_457_carry[10]), .Q(N1760) );
  AND2X1 U3071 ( .IN1(add_div_457_carry[9]), .IN2(EAX_25_), .Q(
        add_div_457_carry[10]) );
  XOR2X1 U3072 ( .IN1(EAX_25_), .IN2(add_div_457_carry[9]), .Q(N1759) );
  AND2X1 U3073 ( .IN1(add_div_457_carry[8]), .IN2(EAX_24_), .Q(
        add_div_457_carry[9]) );
  XOR2X1 U3074 ( .IN1(EAX_24_), .IN2(add_div_457_carry[8]), .Q(N1758) );
  AND2X1 U3075 ( .IN1(add_div_457_carry[7]), .IN2(EAX_23_), .Q(
        add_div_457_carry[8]) );
  XOR2X1 U3076 ( .IN1(EAX_23_), .IN2(add_div_457_carry[7]), .Q(N1757) );
  AND2X1 U3077 ( .IN1(add_div_457_carry[6]), .IN2(EAX_22_), .Q(
        add_div_457_carry[7]) );
  XOR2X1 U3078 ( .IN1(EAX_22_), .IN2(add_div_457_carry[6]), .Q(N1756) );
  AND2X1 U3079 ( .IN1(add_div_457_carry[5]), .IN2(EAX_21_), .Q(
        add_div_457_carry[6]) );
  XOR2X1 U3080 ( .IN1(EAX_21_), .IN2(add_div_457_carry[5]), .Q(N1755) );
  AND2X1 U3081 ( .IN1(add_div_457_carry[4]), .IN2(EAX_20_), .Q(
        add_div_457_carry[5]) );
  XOR2X1 U3082 ( .IN1(EAX_20_), .IN2(add_div_457_carry[4]), .Q(N1754) );
  AND2X1 U3083 ( .IN1(add_div_457_carry[3]), .IN2(EAX_19_), .Q(
        add_div_457_carry[4]) );
  XOR2X1 U3084 ( .IN1(EAX_19_), .IN2(add_div_457_carry[3]), .Q(N1753) );
  AND2X1 U3085 ( .IN1(add_div_457_carry[2]), .IN2(EAX_18_), .Q(
        add_div_457_carry[3]) );
  XOR2X1 U3086 ( .IN1(EAX_18_), .IN2(add_div_457_carry[2]), .Q(N1752) );
  AND2X1 U3087 ( .IN1(add_div_457_carry[1]), .IN2(EAX_17_), .Q(
        add_div_457_carry[2]) );
  XOR2X1 U3088 ( .IN1(EAX_17_), .IN2(add_div_457_carry[1]), .Q(N1751) );
  AND2X1 U3089 ( .IN1(N1749), .IN2(EAX_16_), .Q(add_div_457_carry[1]) );
  XOR2X1 U3090 ( .IN1(EAX_16_), .IN2(N1749), .Q(N1750) );
  XOR2X1 U3091 ( .IN1(add_1_root_add_0_root_add_402_7_B_30_), .IN2(
        add_1_root_add_0_root_add_391_7_carry[30]), .Q(N2415) );
  AND2X1 U3092 ( .IN1(add_1_root_add_0_root_add_391_7_carry[29]), .IN2(
        add_1_root_add_0_root_add_402_7_B_29_), .Q(
        add_1_root_add_0_root_add_391_7_carry[30]) );
  XOR2X1 U3093 ( .IN1(add_1_root_add_0_root_add_402_7_B_29_), .IN2(
        add_1_root_add_0_root_add_391_7_carry[29]), .Q(N2414) );
  AND2X1 U3094 ( .IN1(add_1_root_add_0_root_add_391_7_carry[28]), .IN2(
        add_1_root_add_0_root_add_402_7_B_28_), .Q(
        add_1_root_add_0_root_add_391_7_carry[29]) );
  XOR2X1 U3095 ( .IN1(add_1_root_add_0_root_add_402_7_B_28_), .IN2(
        add_1_root_add_0_root_add_391_7_carry[28]), .Q(N2413) );
  AND2X1 U3096 ( .IN1(add_1_root_add_0_root_add_391_7_carry[27]), .IN2(
        add_1_root_add_0_root_add_402_7_B_27_), .Q(
        add_1_root_add_0_root_add_391_7_carry[28]) );
  XOR2X1 U3097 ( .IN1(add_1_root_add_0_root_add_402_7_B_27_), .IN2(
        add_1_root_add_0_root_add_391_7_carry[27]), .Q(N2412) );
  AND2X1 U3098 ( .IN1(add_1_root_add_0_root_add_391_7_carry[26]), .IN2(
        add_1_root_add_0_root_add_402_7_B_26_), .Q(
        add_1_root_add_0_root_add_391_7_carry[27]) );
  XOR2X1 U3099 ( .IN1(add_1_root_add_0_root_add_402_7_B_26_), .IN2(
        add_1_root_add_0_root_add_391_7_carry[26]), .Q(N2411) );
  AND2X1 U3100 ( .IN1(add_1_root_add_0_root_add_391_7_carry[25]), .IN2(
        add_1_root_add_0_root_add_402_7_B_25_), .Q(
        add_1_root_add_0_root_add_391_7_carry[26]) );
  XOR2X1 U3101 ( .IN1(add_1_root_add_0_root_add_402_7_B_25_), .IN2(
        add_1_root_add_0_root_add_391_7_carry[25]), .Q(N2410) );
  AND2X1 U3102 ( .IN1(add_1_root_add_0_root_add_391_7_carry[24]), .IN2(
        add_1_root_add_0_root_add_402_7_B_24_), .Q(
        add_1_root_add_0_root_add_391_7_carry[25]) );
  XOR2X1 U3103 ( .IN1(add_1_root_add_0_root_add_402_7_B_24_), .IN2(
        add_1_root_add_0_root_add_391_7_carry[24]), .Q(N2409) );
  AND2X1 U3104 ( .IN1(add_1_root_add_0_root_add_402_7_A_23_), .IN2(
        add_1_root_add_0_root_add_402_7_B_23_), .Q(
        add_1_root_add_0_root_add_391_7_carry[24]) );
  XOR2X1 U3105 ( .IN1(add_1_root_add_0_root_add_402_7_B_23_), .IN2(
        add_1_root_add_0_root_add_402_7_A_23_), .Q(N2408) );
  XOR2X1 U3106 ( .IN1(N2392), .IN2(add_2_root_sub_1_root_sub_357_2_carry[7]), 
        .Q(add_2_root_sub_1_root_sub_357_2_SUM_7_) );
  AND2X1 U3107 ( .IN1(add_2_root_sub_1_root_sub_357_2_carry[6]), .IN2(N2391), 
        .Q(add_2_root_sub_1_root_sub_357_2_carry[7]) );
  XOR2X1 U3108 ( .IN1(N2391), .IN2(add_2_root_sub_1_root_sub_357_2_carry[6]), 
        .Q(add_2_root_sub_1_root_sub_357_2_SUM_6_) );
  AND2X1 U3109 ( .IN1(add_2_root_sub_1_root_sub_357_2_carry[5]), .IN2(N2390), 
        .Q(add_2_root_sub_1_root_sub_357_2_carry[6]) );
  XOR2X1 U3110 ( .IN1(N2390), .IN2(add_2_root_sub_1_root_sub_357_2_carry[5]), 
        .Q(add_2_root_sub_1_root_sub_357_2_SUM_5_) );
  AND2X1 U3111 ( .IN1(add_2_root_sub_1_root_sub_357_2_carry[4]), .IN2(N2389), 
        .Q(add_2_root_sub_1_root_sub_357_2_carry[5]) );
  XOR2X1 U3112 ( .IN1(N2389), .IN2(add_2_root_sub_1_root_sub_357_2_carry[4]), 
        .Q(add_2_root_sub_1_root_sub_357_2_SUM_4_) );
  AND2X1 U3113 ( .IN1(add_2_root_sub_1_root_sub_357_2_carry[3]), .IN2(N2388), 
        .Q(add_2_root_sub_1_root_sub_357_2_carry[4]) );
  XOR2X1 U3114 ( .IN1(N2388), .IN2(add_2_root_sub_1_root_sub_357_2_carry[3]), 
        .Q(add_2_root_sub_1_root_sub_357_2_SUM_3_) );
  AND2X1 U3115 ( .IN1(N2386), .IN2(N2387), .Q(
        add_2_root_sub_1_root_sub_357_2_carry[3]) );
  XOR2X1 U3116 ( .IN1(N2387), .IN2(N2386), .Q(
        add_2_root_sub_1_root_sub_357_2_SUM_2_) );
  XOR2X1 U3117 ( .IN1(add_1_root_add_0_root_add_402_7_B_30_), .IN2(
        add_1_root_add_0_root_add_402_7_carry[30]), .Q(N2578) );
  AND2X1 U3118 ( .IN1(add_1_root_add_0_root_add_402_7_carry[29]), .IN2(
        add_1_root_add_0_root_add_402_7_B_29_), .Q(
        add_1_root_add_0_root_add_402_7_carry[30]) );
  XOR2X1 U3119 ( .IN1(add_1_root_add_0_root_add_402_7_B_29_), .IN2(
        add_1_root_add_0_root_add_402_7_carry[29]), .Q(N2577) );
  AND2X1 U3120 ( .IN1(add_1_root_add_0_root_add_402_7_carry[28]), .IN2(
        add_1_root_add_0_root_add_402_7_B_28_), .Q(
        add_1_root_add_0_root_add_402_7_carry[29]) );
  XOR2X1 U3121 ( .IN1(add_1_root_add_0_root_add_402_7_B_28_), .IN2(
        add_1_root_add_0_root_add_402_7_carry[28]), .Q(N2576) );
  AND2X1 U3122 ( .IN1(add_1_root_add_0_root_add_402_7_carry[27]), .IN2(
        add_1_root_add_0_root_add_402_7_B_27_), .Q(
        add_1_root_add_0_root_add_402_7_carry[28]) );
  XOR2X1 U3123 ( .IN1(add_1_root_add_0_root_add_402_7_B_27_), .IN2(
        add_1_root_add_0_root_add_402_7_carry[27]), .Q(N2575) );
  AND2X1 U3124 ( .IN1(add_1_root_add_0_root_add_402_7_carry[26]), .IN2(
        add_1_root_add_0_root_add_402_7_B_26_), .Q(
        add_1_root_add_0_root_add_402_7_carry[27]) );
  XOR2X1 U3125 ( .IN1(add_1_root_add_0_root_add_402_7_B_26_), .IN2(
        add_1_root_add_0_root_add_402_7_carry[26]), .Q(N2574) );
  AND2X1 U3126 ( .IN1(add_1_root_add_0_root_add_402_7_carry[25]), .IN2(
        add_1_root_add_0_root_add_402_7_B_25_), .Q(
        add_1_root_add_0_root_add_402_7_carry[26]) );
  XOR2X1 U3127 ( .IN1(add_1_root_add_0_root_add_402_7_B_25_), .IN2(
        add_1_root_add_0_root_add_402_7_carry[25]), .Q(N2573) );
  AND2X1 U3128 ( .IN1(add_1_root_add_0_root_add_402_7_carry[24]), .IN2(
        add_1_root_add_0_root_add_402_7_B_24_), .Q(
        add_1_root_add_0_root_add_402_7_carry[25]) );
  XOR2X1 U3129 ( .IN1(add_1_root_add_0_root_add_402_7_B_24_), .IN2(
        add_1_root_add_0_root_add_402_7_carry[24]), .Q(N2572) );
  AND2X1 U3130 ( .IN1(add_1_root_add_0_root_add_402_7_A_23_), .IN2(
        add_1_root_add_0_root_add_402_7_B_23_), .Q(
        add_1_root_add_0_root_add_402_7_carry[24]) );
  XOR2X1 U3131 ( .IN1(add_1_root_add_0_root_add_402_7_B_23_), .IN2(
        add_1_root_add_0_root_add_402_7_A_23_), .Q(N2571) );
  AND2X1 U3132 ( .IN1(InstQueueRd_Addr[3]), .IN2(add_495_carry[3]), .Q(
        add_495_carry[4]) );
  XOR2X1 U3133 ( .IN1(add_495_carry[3]), .IN2(InstQueueRd_Addr[3]), .Q(N2740)
         );
  AND2X1 U3134 ( .IN1(InstQueueRd_Addr[2]), .IN2(InstQueueRd_Addr[1]), .Q(
        add_495_carry[3]) );
  XOR2X1 U3135 ( .IN1(InstQueueRd_Addr[1]), .IN2(InstQueueRd_Addr[2]), .Q(
        N2739) );
  XOR2X1 U3136 ( .IN1(n3871), .IN2(r679_carry[4]), .Q(r680_B_4_) );
  OR2X1 U3137 ( .IN1(n1552), .IN2(N1239), .Q(r679_carry[1]) );
  XNOR2X1 U3138 ( .IN1(N1239), .IN2(n1552), .Q(gte_355_B_0_) );
  ISOLANDX1 U3139 ( .D(N3417), .ISO(N3989), .Q(n3686) );
  ISOLANDX1 U3140 ( .D(N1239), .ISO(N3420), .Q(n3683) );
  ISOLANDX1 U3141 ( .D(n3683), .ISO(N3419), .Q(n3682) );
  OAI222X1 U3142 ( .IN1(n3683), .IN2(n3688), .IN3(N3991), .IN4(n3682), .IN5(
        N3990), .IN6(N3423), .QN(n3684) );
  OA21X1 U3143 ( .IN1(N3418), .IN2(n1554), .IN3(n3684), .Q(n3685) );
  OA22X1 U3144 ( .IN1(n3686), .IN2(n3685), .IN3(N3417), .IN4(n1553), .Q(n3687)
         );
  NOR2X0 U3145 ( .IN1(N3427), .IN2(n3687), .QN(N3415) );
  OR2X1 U3146 ( .IN1(n3689), .IN2(N3427), .Q(N3428) );
  OR2X1 U3147 ( .IN1(n3691), .IN2(N3493), .Q(N3494) );
  INVX0 U3148 ( .IN(n3874), .QN(add_div_311_A_0_) );
  INVX0 U3149 ( .IN(RESET), .QN(n5315) );
  AO222X1 U3150 ( .IN1(n3875), .IN2(n3876), .IN3(n3877), .IN4(n3878), .IN5(
        n3879), .IN6(N2737), .Q(N2401) );
  AO221X1 U3151 ( .IN1(n3880), .IN2(n3875), .IN3(n3881), .IN4(n3878), .IN5(
        n3882), .Q(N2393) );
  AO22X1 U3152 ( .IN1(n3883), .IN2(n3877), .IN3(n3884), .IN4(n3876), .Q(n3882)
         );
  INVX0 U3153 ( .IN(n3885), .QN(n3878) );
  AO222X1 U3154 ( .IN1(n3881), .IN2(n3883), .IN3(n3880), .IN4(n3884), .IN5(
        n3886), .IN6(n1552), .Q(N2385) );
  OAI222X1 U3155 ( .IN1(n3885), .IN2(n3887), .IN3(n3888), .IN4(n3889), .IN5(
        N2737), .IN6(n3890), .QN(add_1_root_add_0_root_add_402_7_B_23_) );
  INVX0 U3156 ( .IN(n3879), .QN(n3890) );
  MUX21X1 U3157 ( .IN1(n3891), .IN2(n3883), .S(n1550), .Q(n3879) );
  AOI221X1 U3158 ( .IN1(n3758), .IN2(n3126), .IN3(n3790), .IN4(n3116), .IN5(
        n3892), .QN(n3883) );
  AO22X1 U3159 ( .IN1(n3726), .IN2(n3181), .IN3(n3694), .IN4(n3137), .Q(n3892)
         );
  OA221X1 U3160 ( .IN1(n3108), .IN2(n2876), .IN3(n3121), .IN4(n2854), .IN5(
        n3895), .Q(n3891) );
  OA22X1 U3161 ( .IN1(n3142), .IN2(n2848), .IN3(n3166), .IN4(n2869), .Q(n3895)
         );
  OA221X1 U3162 ( .IN1(n3814), .IN2(n3111), .IN3(n3782), .IN4(n3120), .IN5(
        n3898), .Q(n3888) );
  OA22X1 U3163 ( .IN1(n3718), .IN2(n3134), .IN3(n3750), .IN4(n3159), .Q(n3898)
         );
  AO221X1 U3164 ( .IN1(n3766), .IN2(n3130), .IN3(n3798), .IN4(n3117), .IN5(
        n3899), .Q(n3885) );
  AO22X1 U3165 ( .IN1(n3734), .IN2(n3181), .IN3(n3702), .IN4(n3156), .Q(n3899)
         );
  AO222X1 U3166 ( .IN1(n3900), .IN2(n3875), .IN3(n3901), .IN4(n3877), .IN5(
        n3902), .IN6(N2737), .Q(N2402) );
  AO221X1 U3167 ( .IN1(n3903), .IN2(n3875), .IN3(n3901), .IN4(n3881), .IN5(
        n3904), .Q(N2394) );
  AO22X1 U3168 ( .IN1(n3905), .IN2(n3877), .IN3(n3900), .IN4(n3884), .Q(n3904)
         );
  INVX0 U3169 ( .IN(n3906), .QN(n3901) );
  AO222X1 U3170 ( .IN1(n3905), .IN2(n3881), .IN3(n3903), .IN4(n3884), .IN5(
        n3907), .IN6(n1552), .Q(N2386) );
  OAI222X1 U3171 ( .IN1(n3887), .IN2(n3906), .IN3(n3908), .IN4(n3889), .IN5(
        N2737), .IN6(n3909), .QN(add_1_root_add_0_root_add_402_7_B_24_) );
  INVX0 U3172 ( .IN(n3902), .QN(n3909) );
  MUX21X1 U3173 ( .IN1(n3905), .IN2(n3910), .S(InstQueueRd_Addr[1]), .Q(n3902)
         );
  OA221X1 U3174 ( .IN1(n3106), .IN2(test_so14), .IN3(n3120), .IN4(n2855), 
        .IN5(n3911), .Q(n3910) );
  OA22X1 U3175 ( .IN1(n3140), .IN2(n2861), .IN3(n3164), .IN4(n2884), .Q(n3911)
         );
  AOI221X1 U3176 ( .IN1(n3759), .IN2(n3126), .IN3(n3791), .IN4(n3116), .IN5(
        n3912), .QN(n3905) );
  AO22X1 U3177 ( .IN1(n3727), .IN2(n3163), .IN3(n3695), .IN4(n3156), .Q(n3912)
         );
  OA221X1 U3178 ( .IN1(n3815), .IN2(n3111), .IN3(n3783), .IN4(n3120), .IN5(
        n3913), .Q(n3908) );
  OA22X1 U3179 ( .IN1(n3719), .IN2(n3134), .IN3(n3751), .IN4(n3159), .Q(n3913)
         );
  AO221X1 U3180 ( .IN1(n3767), .IN2(n3130), .IN3(n3799), .IN4(n3117), .IN5(
        n3914), .Q(n3906) );
  AO22X1 U3181 ( .IN1(n3735), .IN2(n3173), .IN3(n3703), .IN4(n3155), .Q(n3914)
         );
  AO222X1 U3182 ( .IN1(n3915), .IN2(n3875), .IN3(n3916), .IN4(n3877), .IN5(
        n3917), .IN6(N2737), .Q(N2403) );
  AO221X1 U3183 ( .IN1(n3918), .IN2(n3875), .IN3(n3916), .IN4(n3881), .IN5(
        n3919), .Q(N2395) );
  AO22X1 U3184 ( .IN1(n3920), .IN2(n3877), .IN3(n3915), .IN4(n3884), .Q(n3919)
         );
  INVX0 U3185 ( .IN(n3921), .QN(n3916) );
  AO222X1 U3186 ( .IN1(n3920), .IN2(n3881), .IN3(n3918), .IN4(n3884), .IN5(
        n3922), .IN6(n1552), .Q(N2387) );
  OAI222X1 U3187 ( .IN1(n3887), .IN2(n3921), .IN3(n3923), .IN4(n3889), .IN5(
        N2737), .IN6(n3924), .QN(add_1_root_add_0_root_add_402_7_B_25_) );
  INVX0 U3188 ( .IN(n3917), .QN(n3924) );
  MUX21X1 U3189 ( .IN1(n3920), .IN2(n3925), .S(InstQueueRd_Addr[1]), .Q(n3917)
         );
  OA221X1 U3190 ( .IN1(n3110), .IN2(n2878), .IN3(n3123), .IN4(n2856), .IN5(
        n3926), .Q(n3925) );
  OA22X1 U3191 ( .IN1(n3140), .IN2(n2862), .IN3(n3164), .IN4(test_so11), .Q(
        n3926) );
  AOI221X1 U3192 ( .IN1(n3760), .IN2(n3127), .IN3(n3792), .IN4(n3115), .IN5(
        n3927), .QN(n3920) );
  AO22X1 U3193 ( .IN1(n3728), .IN2(n3180), .IN3(n3696), .IN4(n3155), .Q(n3927)
         );
  OA221X1 U3194 ( .IN1(n3816), .IN2(n3110), .IN3(n3784), .IN4(n3120), .IN5(
        n3928), .Q(n3923) );
  OA22X1 U3195 ( .IN1(n3720), .IN2(n3134), .IN3(n3752), .IN4(n3159), .Q(n3928)
         );
  AO221X1 U3196 ( .IN1(n3768), .IN2(n3130), .IN3(n3800), .IN4(n3112), .IN5(
        n3929), .Q(n3921) );
  AO22X1 U3197 ( .IN1(n3736), .IN2(n3180), .IN3(n3704), .IN4(n3154), .Q(n3929)
         );
  AO222X1 U3198 ( .IN1(n3930), .IN2(n3875), .IN3(n3931), .IN4(n3877), .IN5(
        n3932), .IN6(N2737), .Q(N2404) );
  AO221X1 U3199 ( .IN1(n3933), .IN2(n3875), .IN3(n3931), .IN4(n3881), .IN5(
        n3934), .Q(N2396) );
  AO22X1 U3200 ( .IN1(n3935), .IN2(n3877), .IN3(n3930), .IN4(n3884), .Q(n3934)
         );
  INVX0 U3201 ( .IN(n3936), .QN(n3931) );
  AO222X1 U3202 ( .IN1(n3935), .IN2(n3881), .IN3(n3933), .IN4(n3884), .IN5(
        n3937), .IN6(n1552), .Q(N2388) );
  OAI222X1 U3203 ( .IN1(n3887), .IN2(n3936), .IN3(n3938), .IN4(n3889), .IN5(
        N2737), .IN6(n3939), .QN(add_1_root_add_0_root_add_402_7_B_26_) );
  INVX0 U3204 ( .IN(n3932), .QN(n3939) );
  MUX21X1 U3205 ( .IN1(n3935), .IN2(n3940), .S(InstQueueRd_Addr[1]), .Q(n3932)
         );
  OA221X1 U3206 ( .IN1(n3106), .IN2(n2871), .IN3(n3123), .IN4(n2849), .IN5(
        n3941), .Q(n3940) );
  OA22X1 U3207 ( .IN1(n3140), .IN2(n2863), .IN3(n3159), .IN4(n2886), .Q(n3941)
         );
  AOI221X1 U3208 ( .IN1(n3761), .IN2(n3126), .IN3(n3793), .IN4(n3115), .IN5(
        n3942), .QN(n3935) );
  AO22X1 U3209 ( .IN1(n3729), .IN2(n3179), .IN3(n3697), .IN4(n3154), .Q(n3942)
         );
  OA221X1 U3210 ( .IN1(n3817), .IN2(n3110), .IN3(n3785), .IN4(n3120), .IN5(
        n3943), .Q(n3938) );
  OA22X1 U3211 ( .IN1(n3721), .IN2(n3134), .IN3(n3753), .IN4(n3159), .Q(n3943)
         );
  AO221X1 U3212 ( .IN1(n3769), .IN2(n3130), .IN3(n3801), .IN4(n3112), .IN5(
        n3944), .Q(n3936) );
  AO22X1 U3213 ( .IN1(n3737), .IN2(n3173), .IN3(n3705), .IN4(n3153), .Q(n3944)
         );
  AO222X1 U3214 ( .IN1(n3945), .IN2(n3875), .IN3(n3946), .IN4(n3877), .IN5(
        n3947), .IN6(N2737), .Q(N2405) );
  AO221X1 U3215 ( .IN1(n3948), .IN2(n3875), .IN3(n3946), .IN4(n3881), .IN5(
        n3949), .Q(N2397) );
  AO22X1 U3216 ( .IN1(n3950), .IN2(n3877), .IN3(n3945), .IN4(n3884), .Q(n3949)
         );
  INVX0 U3217 ( .IN(n3951), .QN(n3946) );
  AO222X1 U3218 ( .IN1(n3950), .IN2(n3881), .IN3(n3948), .IN4(n3884), .IN5(
        n3952), .IN6(n1552), .Q(N2389) );
  OAI222X1 U3219 ( .IN1(n3887), .IN2(n3951), .IN3(n3953), .IN4(n3889), .IN5(
        N2737), .IN6(n3954), .QN(add_1_root_add_0_root_add_402_7_B_27_) );
  INVX0 U3220 ( .IN(n3947), .QN(n3954) );
  MUX21X1 U3221 ( .IN1(n3950), .IN2(n3955), .S(InstQueueRd_Addr[1]), .Q(n3947)
         );
  OA221X1 U3222 ( .IN1(n3106), .IN2(n2872), .IN3(n3123), .IN4(n2850), .IN5(
        n3956), .Q(n3955) );
  OA22X1 U3223 ( .IN1(n3141), .IN2(n2857), .IN3(n3159), .IN4(n2879), .Q(n3956)
         );
  AOI221X1 U3224 ( .IN1(n3762), .IN2(n3126), .IN3(n3794), .IN4(n3117), .IN5(
        n3957), .QN(n3950) );
  AO22X1 U3225 ( .IN1(n3730), .IN2(n3179), .IN3(n3698), .IN4(n3153), .Q(n3957)
         );
  OA221X1 U3226 ( .IN1(n3818), .IN2(n3106), .IN3(n3786), .IN4(n3120), .IN5(
        n3958), .Q(n3953) );
  OA22X1 U3227 ( .IN1(n3722), .IN2(n3134), .IN3(n3754), .IN4(n3157), .Q(n3958)
         );
  AO221X1 U3228 ( .IN1(n3770), .IN2(n3130), .IN3(n3802), .IN4(n3113), .IN5(
        n3959), .Q(n3951) );
  AO22X1 U3229 ( .IN1(n3738), .IN2(n3179), .IN3(n3706), .IN4(n3151), .Q(n3959)
         );
  AO222X1 U3230 ( .IN1(n3960), .IN2(n3875), .IN3(n3961), .IN4(n3877), .IN5(
        n3962), .IN6(N2737), .Q(N2406) );
  AO221X1 U3231 ( .IN1(n3963), .IN2(n3875), .IN3(n3961), .IN4(n3881), .IN5(
        n3964), .Q(N2398) );
  AO22X1 U3232 ( .IN1(n3965), .IN2(n3877), .IN3(n3960), .IN4(n3884), .Q(n3964)
         );
  INVX0 U3233 ( .IN(n3966), .QN(n3961) );
  AO222X1 U3234 ( .IN1(n3965), .IN2(n3881), .IN3(n3963), .IN4(n3884), .IN5(
        n3967), .IN6(n1552), .Q(N2390) );
  OAI222X1 U3235 ( .IN1(n3887), .IN2(n3966), .IN3(n3968), .IN4(n3889), .IN5(
        N2737), .IN6(n3969), .QN(add_1_root_add_0_root_add_402_7_B_28_) );
  INVX0 U3236 ( .IN(n3962), .QN(n3969) );
  MUX21X1 U3237 ( .IN1(n3970), .IN2(n3965), .S(n1550), .Q(n3962) );
  AOI221X1 U3238 ( .IN1(n3763), .IN2(n3127), .IN3(n3795), .IN4(n3115), .IN5(
        n3971), .QN(n3965) );
  AO22X1 U3239 ( .IN1(n3731), .IN2(n3178), .IN3(n3699), .IN4(n3148), .Q(n3971)
         );
  OA221X1 U3240 ( .IN1(n3107), .IN2(n2873), .IN3(n3123), .IN4(n2851), .IN5(
        n3972), .Q(n3970) );
  OA22X1 U3241 ( .IN1(n3141), .IN2(n2858), .IN3(n3159), .IN4(n2880), .Q(n3972)
         );
  OA221X1 U3242 ( .IN1(n3819), .IN2(n3110), .IN3(n3787), .IN4(n3123), .IN5(
        n3973), .Q(n3968) );
  OA22X1 U3243 ( .IN1(n3723), .IN2(n3134), .IN3(n3755), .IN4(n3159), .Q(n3973)
         );
  AO221X1 U3244 ( .IN1(n3771), .IN2(n3125), .IN3(n3803), .IN4(n3114), .IN5(
        n3974), .Q(n3966) );
  AO22X1 U3245 ( .IN1(n3739), .IN2(n3178), .IN3(n3707), .IN4(n3152), .Q(n3974)
         );
  AO222X1 U3246 ( .IN1(n3975), .IN2(n3875), .IN3(n3976), .IN4(n3877), .IN5(
        n3977), .IN6(N2737), .Q(N2407) );
  AO221X1 U3247 ( .IN1(n3978), .IN2(n3875), .IN3(n3976), .IN4(n3881), .IN5(
        n3979), .Q(N2399) );
  AO22X1 U3248 ( .IN1(n3980), .IN2(n3877), .IN3(n3975), .IN4(n3884), .Q(n3979)
         );
  INVX0 U3249 ( .IN(n3981), .QN(n3976) );
  AO222X1 U3250 ( .IN1(n3980), .IN2(n3881), .IN3(n3978), .IN4(n3884), .IN5(
        n3982), .IN6(n1552), .Q(N2391) );
  OAI222X1 U3251 ( .IN1(n3887), .IN2(n3981), .IN3(n3983), .IN4(n3889), .IN5(
        N2737), .IN6(n3984), .QN(add_1_root_add_0_root_add_402_7_B_29_) );
  INVX0 U3252 ( .IN(n3977), .QN(n3984) );
  MUX21X1 U3253 ( .IN1(n3985), .IN2(n3980), .S(n1550), .Q(n3977) );
  AOI221X1 U3254 ( .IN1(n3764), .IN2(n3127), .IN3(n3796), .IN4(n3115), .IN5(
        n3986), .QN(n3980) );
  AO22X1 U3255 ( .IN1(n3732), .IN2(n3177), .IN3(n3700), .IN4(n3152), .Q(n3986)
         );
  OA221X1 U3256 ( .IN1(n3107), .IN2(n2874), .IN3(n3120), .IN4(n2852), .IN5(
        n3987), .Q(n3985) );
  OA22X1 U3257 ( .IN1(n3141), .IN2(n2859), .IN3(n3157), .IN4(n2881), .Q(n3987)
         );
  OA221X1 U3258 ( .IN1(n3820), .IN2(n3106), .IN3(n3788), .IN4(n3120), .IN5(
        n3988), .Q(n3983) );
  OA22X1 U3259 ( .IN1(n3724), .IN2(n3144), .IN3(n3756), .IN4(n3157), .Q(n3988)
         );
  AO221X1 U3260 ( .IN1(n3772), .IN2(n3131), .IN3(n3804), .IN4(n3113), .IN5(
        n3989), .Q(n3981) );
  AO22X1 U3261 ( .IN1(n3740), .IN2(n3177), .IN3(n3708), .IN4(n3151), .Q(n3989)
         );
  AO222X1 U3262 ( .IN1(n3990), .IN2(n3875), .IN3(n3991), .IN4(n3877), .IN5(
        n3992), .IN6(N2737), .Q(add_1_root_add_0_root_add_402_7_A_23_) );
  AO221X1 U3263 ( .IN1(n3993), .IN2(n3875), .IN3(n3991), .IN4(n3881), .IN5(
        n3994), .Q(N2400) );
  AO22X1 U3264 ( .IN1(n3995), .IN2(n3877), .IN3(n3990), .IN4(n3884), .Q(n3994)
         );
  INVX0 U3265 ( .IN(n3997), .QN(n3991) );
  AO222X1 U3266 ( .IN1(n3995), .IN2(n3881), .IN3(n3993), .IN4(n3884), .IN5(
        n3999), .IN6(n1552), .Q(N2392) );
  OAI222X1 U3267 ( .IN1(n3887), .IN2(n3997), .IN3(n4000), .IN4(n3889), .IN5(
        N2737), .IN6(n4001), .QN(add_1_root_add_0_root_add_402_7_B_30_) );
  INVX0 U3268 ( .IN(n3992), .QN(n4001) );
  MUX21X1 U3269 ( .IN1(n4002), .IN2(n3995), .S(n1550), .Q(n3992) );
  AOI221X1 U3270 ( .IN1(n3765), .IN2(n3128), .IN3(n3797), .IN4(n3117), .IN5(
        n4003), .QN(n3995) );
  AO22X1 U3271 ( .IN1(n3733), .IN2(n3176), .IN3(n3701), .IN4(n3151), .Q(n4003)
         );
  OA221X1 U3272 ( .IN1(n3107), .IN2(n2875), .IN3(n3121), .IN4(n2853), .IN5(
        n4004), .Q(n4002) );
  OA22X1 U3273 ( .IN1(n3141), .IN2(n2860), .IN3(n3165), .IN4(n2882), .Q(n4004)
         );
  OA221X1 U3274 ( .IN1(n3821), .IN2(n3110), .IN3(n3789), .IN4(n3123), .IN5(
        n4005), .Q(n4000) );
  OA22X1 U3275 ( .IN1(n3725), .IN2(n3132), .IN3(n3757), .IN4(n3157), .Q(n4005)
         );
  AO221X1 U3276 ( .IN1(n3773), .IN2(n3125), .IN3(n3805), .IN4(n3114), .IN5(
        n4006), .Q(n3997) );
  AO22X1 U3277 ( .IN1(n3741), .IN2(n3176), .IN3(n3709), .IN4(n3150), .Q(n4006)
         );
  MUX21X1 U3278 ( .IN1(n4007), .IN2(n2889), .S(n4008), .Q(n2841) );
  NOR4X0 U3279 ( .IN1(n4009), .IN2(n4010), .IN3(n4011), .IN4(n4012), .QN(n4008) );
  NOR2X0 U3280 ( .IN1(n2949), .IN2(n4013), .QN(n4010) );
  NAND3X0 U3281 ( .IN1(n4014), .IN2(n3185), .IN3(n4016), .QN(n4007) );
  NAND2X0 U3282 ( .IN1(n4017), .IN2(n4018), .QN(n4014) );
  OAI221X1 U3283 ( .IN1(n4019), .IN2(n4020), .IN3(n2868), .IN4(n4021), .IN5(
        n2948), .QN(n4018) );
  AND2X1 U3284 ( .IN1(n4022), .IN2(n4023), .Q(n2840) );
  NAND4X0 U3285 ( .IN1(NA_n), .IN2(n3211), .IN3(n4025), .IN4(n4026), .QN(n4023) );
  NAND4X0 U3286 ( .IN1(n4027), .IN2(n4028), .IN3(n4029), .IN4(n4030), .QN(
        n4022) );
  NAND3X0 U3287 ( .IN1(n2949), .IN2(n4031), .IN3(n4032), .QN(n4029) );
  NAND2X0 U3288 ( .IN1(n1596), .IN2(n4033), .QN(n4031) );
  AO21X1 U3289 ( .IN1(n4026), .IN2(n4034), .IN3(n4033), .Q(n4028) );
  OR2X1 U3290 ( .IN1(n4025), .IN2(n2889), .Q(n4034) );
  NAND3X0 U3291 ( .IN1(n4027), .IN2(n4035), .IN3(n4036), .QN(n2839) );
  AO21X1 U3292 ( .IN1(n4037), .IN2(n4038), .IN3(n1596), .Q(n4035) );
  NAND2X0 U3293 ( .IN1(n4039), .IN2(n4033), .QN(n4038) );
  AND2X1 U3294 ( .IN1(n4040), .IN2(n4041), .Q(n4027) );
  NAND3X0 U3295 ( .IN1(n2867), .IN2(n2847), .IN3(n2949), .QN(n4041) );
  NAND4X0 U3296 ( .IN1(n4036), .IN2(n4042), .IN3(n4043), .IN4(n4044), .QN(
        n2838) );
  AO21X1 U3297 ( .IN1(n4037), .IN2(n4026), .IN3(n2889), .Q(n4043) );
  ISOLANDX1 U3298 ( .D(n4025), .ISO(n4032), .Q(n4037) );
  NAND3X0 U3299 ( .IN1(n1434), .IN2(n4045), .IN3(n1435), .QN(n4025) );
  NAND2X0 U3300 ( .IN1(n4039), .IN2(HOLD), .QN(n4042) );
  INVX0 U3301 ( .IN(n4026), .QN(n4039) );
  NAND2X0 U3302 ( .IN1(n4045), .IN2(n2867), .QN(n4026) );
  AOI22X1 U3303 ( .IN1(n4019), .IN2(n4046), .IN3(n4032), .IN4(n4047), .QN(
        n4036) );
  NAND2X0 U3304 ( .IN1(n2948), .IN2(n4033), .QN(n4047) );
  INVX0 U3305 ( .IN(HOLD), .QN(n4033) );
  INVX0 U3306 ( .IN(n4048), .QN(n4032) );
  OR4X1 U3307 ( .IN1(n3212), .IN2(HOLD), .IN3(NA_n), .IN4(n1596), .Q(n4046) );
  AO21X1 U3308 ( .IN1(n3211), .IN2(ADS_n), .IN3(n4050), .Q(n2837) );
  INVX0 U3309 ( .IN(n4051), .QN(n4050) );
  AO21X1 U3310 ( .IN1(n4051), .IN2(n2868), .IN3(n4052), .Q(n2836) );
  AO22X1 U3311 ( .IN1(n4051), .IN2(test_so2), .IN3(n4053), .IN4(n4054), .Q(
        n2835) );
  INVX0 U3312 ( .IN(BS16_n), .QN(n4054) );
  AO21X1 U3313 ( .IN1(n4051), .IN2(n2864), .IN3(n4052), .Q(n2834) );
  AO21X1 U3314 ( .IN1(BS16_n), .IN2(n4053), .IN3(n4055), .Q(n4052) );
  NOR2X0 U3315 ( .IN1(n4053), .IN2(n4055), .QN(n4051) );
  INVX0 U3316 ( .IN(n4044), .QN(n4055) );
  NAND2X0 U3317 ( .IN1(n4040), .IN2(n4048), .QN(n4053) );
  NAND3X0 U3318 ( .IN1(n2847), .IN2(n4045), .IN3(n1434), .QN(n4048) );
  OR2X1 U3319 ( .IN1(n4056), .IN2(n4057), .Q(n2833) );
  AO222X1 U3320 ( .IN1(rEIP_31_), .IN2(n2950), .IN3(N1062), .IN4(n3218), .IN5(
        n2956), .IN6(PhyAddrPointer_31_), .Q(n4057) );
  AO221X1 U3321 ( .IN1(n3225), .IN2(N1954), .IN3(N1800), .IN4(n3231), .IN5(
        n4061), .Q(n4056) );
  AO22X1 U3322 ( .IN1(N1029), .IN2(n3238), .IN3(N1987), .IN4(n3251), .Q(n4061)
         );
  NAND4X0 U3323 ( .IN1(n4064), .IN2(n4065), .IN3(n4066), .IN4(n4067), .QN(
        n2832) );
  OA22X1 U3324 ( .IN1(n3257), .IN2(n4069), .IN3(n3264), .IN4(n4071), .Q(n4067)
         );
  AOI22X1 U3325 ( .IN1(N1510), .IN2(n3276), .IN3(n34), .IN4(n3288), .QN(n4066)
         );
  AOI22X1 U3326 ( .IN1(N2887), .IN2(n3300), .IN3(N2447), .IN4(n3312), .QN(
        n4065) );
  OA22X1 U3327 ( .IN1(n3869), .IN2(n3324), .IN3(n2866), .IN4(n3194), .Q(n4064)
         );
  MUX21X1 U3328 ( .IN1(n4077), .IN2(n4078), .S(n4079), .Q(n2831) );
  AO22X1 U3329 ( .IN1(n4017), .IN2(n4080), .IN3(n4081), .IN4(n4082), .Q(n4077)
         );
  MUX21X1 U3330 ( .IN1(n4083), .IN2(n2842), .S(n4084), .Q(n2830) );
  NAND3X0 U3331 ( .IN1(n4085), .IN2(n4086), .IN3(n4087), .QN(n4083) );
  OA221X1 U3332 ( .IN1(N3494), .IN2(n4088), .IN3(n4016), .IN4(n2948), .IN5(
        n4013), .Q(n4087) );
  NAND2X0 U3333 ( .IN1(n4089), .IN2(InstQueueRd_Addr[4]), .QN(n4086) );
  NAND4X0 U3334 ( .IN1(n4090), .IN2(n4013), .IN3(n4091), .IN4(n4092), .QN(
        n2829) );
  OA221X1 U3335 ( .IN1(n2949), .IN2(n4093), .IN3(n1490), .IN4(n4094), .IN5(
        n3396), .Q(n4092) );
  NAND3X0 U3336 ( .IN1(n4088), .IN2(n4095), .IN3(n4096), .QN(n2828) );
  NAND2X0 U3337 ( .IN1(n4084), .IN2(n4097), .QN(n4096) );
  MUX21X1 U3338 ( .IN1(n4098), .IN2(n2844), .S(n4084), .Q(n2827) );
  INVX0 U3339 ( .IN(n4094), .QN(n4084) );
  NAND4X0 U3340 ( .IN1(n4016), .IN2(n4099), .IN3(n4085), .IN4(n4100), .QN(
        n4094) );
  AND3X1 U3341 ( .IN1(n4088), .IN2(n4095), .IN3(n4101), .Q(n4100) );
  OR2X1 U3342 ( .IN1(n4102), .IN2(n4091), .Q(n4101) );
  AND4X1 U3343 ( .IN1(n4103), .IN2(n4104), .IN3(n3105), .IN4(n3194), .Q(n4085)
         );
  NAND2X0 U3344 ( .IN1(n4017), .IN2(n4105), .QN(n4104) );
  NAND4X0 U3345 ( .IN1(N3415), .IN2(n4106), .IN3(n4107), .IN4(n4108), .QN(
        n4105) );
  NOR2X0 U3346 ( .IN1(N3428), .IN2(n4109), .QN(n4107) );
  AOI21X1 U3347 ( .IN1(n1590), .IN2(n3873), .IN3(n4110), .QN(n4109) );
  NAND2X0 U3348 ( .IN1(n3344), .IN2(n2948), .QN(n4099) );
  NOR2X0 U3349 ( .IN1(n4112), .IN2(n4009), .QN(n4016) );
  INVX0 U3350 ( .IN(n4093), .QN(n4009) );
  NAND3X0 U3351 ( .IN1(n4113), .IN2(n4091), .IN3(n4114), .QN(n4098) );
  MUX21X1 U3352 ( .IN1(n4115), .IN2(n4093), .S(n2949), .Q(n4114) );
  NAND3X0 U3353 ( .IN1(n1490), .IN2(n2844), .IN3(n4116), .QN(n4093) );
  AO22X1 U3354 ( .IN1(n3355), .IN2(N1954), .IN3(N1650), .IN4(n3362), .Q(n2826)
         );
  AO222X1 U3355 ( .IN1(N1619), .IN2(n3362), .IN3(N2548), .IN4(n3367), .IN5(
        n3355), .IN6(EBX_0_), .Q(n2825) );
  AO222X1 U3356 ( .IN1(N1620), .IN2(n3361), .IN3(N2549), .IN4(n3367), .IN5(
        n3355), .IN6(EBX_1_), .Q(n2824) );
  AO222X1 U3357 ( .IN1(N1621), .IN2(n3361), .IN3(N2550), .IN4(n3367), .IN5(
        n3354), .IN6(EBX_2_), .Q(n2823) );
  AO222X1 U3358 ( .IN1(N1622), .IN2(n3361), .IN3(N2551), .IN4(n3367), .IN5(
        n3354), .IN6(EBX_3_), .Q(n2822) );
  AO222X1 U3359 ( .IN1(N1623), .IN2(n3361), .IN3(N2552), .IN4(n3367), .IN5(
        n3354), .IN6(EBX_4_), .Q(n2821) );
  AO222X1 U3360 ( .IN1(N1624), .IN2(n3361), .IN3(N2553), .IN4(n3368), .IN5(
        n3354), .IN6(EBX_5_), .Q(n2820) );
  AO222X1 U3361 ( .IN1(N1625), .IN2(n3360), .IN3(N2554), .IN4(n3368), .IN5(
        n3354), .IN6(EBX_6_), .Q(n2819) );
  AO222X1 U3362 ( .IN1(N1626), .IN2(n3360), .IN3(N2555), .IN4(n3368), .IN5(
        n3353), .IN6(EBX_7_), .Q(n2818) );
  AO222X1 U3363 ( .IN1(N1627), .IN2(n3360), .IN3(N2393), .IN4(n3368), .IN5(
        n3353), .IN6(EBX_8_), .Q(n2817) );
  AO222X1 U3364 ( .IN1(N1628), .IN2(n3360), .IN3(N2394), .IN4(n3368), .IN5(
        n3353), .IN6(EBX_9_), .Q(n2816) );
  AO222X1 U3365 ( .IN1(N1629), .IN2(n3360), .IN3(N2395), .IN4(n3369), .IN5(
        n3353), .IN6(EBX_10_), .Q(n2815) );
  AO222X1 U3366 ( .IN1(N1630), .IN2(n3359), .IN3(N2396), .IN4(n3369), .IN5(
        n3353), .IN6(EBX_11_), .Q(n2814) );
  AO222X1 U3367 ( .IN1(N1631), .IN2(n3359), .IN3(N2397), .IN4(n3369), .IN5(
        n3352), .IN6(EBX_12_), .Q(n2813) );
  AO222X1 U3368 ( .IN1(N1632), .IN2(n3359), .IN3(N2398), .IN4(n3369), .IN5(
        n3352), .IN6(EBX_13_), .Q(n2812) );
  AO222X1 U3369 ( .IN1(N1633), .IN2(n3359), .IN3(N2399), .IN4(n3369), .IN5(
        n3352), .IN6(EBX_14_), .Q(n2811) );
  AO222X1 U3370 ( .IN1(N1634), .IN2(n3359), .IN3(N2400), .IN4(n3370), .IN5(
        n3352), .IN6(EBX_15_), .Q(n2810) );
  AO222X1 U3371 ( .IN1(N1635), .IN2(n3358), .IN3(N2401), .IN4(n3370), .IN5(
        n3351), .IN6(EBX_16_), .Q(n2809) );
  AO222X1 U3372 ( .IN1(N1636), .IN2(n3358), .IN3(N2402), .IN4(n3370), .IN5(
        n3351), .IN6(EBX_17_), .Q(n2808) );
  AO222X1 U3373 ( .IN1(N1637), .IN2(n3358), .IN3(N2403), .IN4(n3370), .IN5(
        n3351), .IN6(EBX_18_), .Q(n2807) );
  AO222X1 U3374 ( .IN1(N1638), .IN2(n3358), .IN3(N2404), .IN4(n3370), .IN5(
        n3351), .IN6(test_so6), .Q(n2806) );
  AO222X1 U3375 ( .IN1(N1639), .IN2(n3358), .IN3(N2405), .IN4(n3371), .IN5(
        n3351), .IN6(EBX_20_), .Q(n2805) );
  AO222X1 U3376 ( .IN1(N1640), .IN2(n3357), .IN3(N2406), .IN4(n3371), .IN5(
        n3350), .IN6(EBX_21_), .Q(n2804) );
  AO222X1 U3377 ( .IN1(N1641), .IN2(n3357), .IN3(N2407), .IN4(n3371), .IN5(
        n3350), .IN6(EBX_22_), .Q(n2803) );
  AO222X1 U3378 ( .IN1(N1642), .IN2(n3357), .IN3(N2571), .IN4(n3371), .IN5(
        n3350), .IN6(EBX_23_), .Q(n2802) );
  AO222X1 U3379 ( .IN1(N1643), .IN2(n3357), .IN3(N2572), .IN4(n3371), .IN5(
        n3352), .IN6(EBX_24_), .Q(n2801) );
  AO222X1 U3380 ( .IN1(N1644), .IN2(n3357), .IN3(N2573), .IN4(n3372), .IN5(
        n3350), .IN6(EBX_25_), .Q(n2800) );
  AO222X1 U3381 ( .IN1(N1645), .IN2(n3356), .IN3(N2574), .IN4(n3372), .IN5(
        n3350), .IN6(EBX_26_), .Q(n2799) );
  AO222X1 U3382 ( .IN1(N1646), .IN2(n3356), .IN3(N2575), .IN4(n3372), .IN5(
        n3349), .IN6(EBX_27_), .Q(n2798) );
  AO222X1 U3383 ( .IN1(N1647), .IN2(n3356), .IN3(N2576), .IN4(n3372), .IN5(
        n3349), .IN6(EBX_28_), .Q(n2797) );
  AO222X1 U3384 ( .IN1(N1648), .IN2(n3356), .IN3(N2577), .IN4(n3372), .IN5(
        n3349), .IN6(EBX_29_), .Q(n2796) );
  AO222X1 U3385 ( .IN1(N1649), .IN2(n3356), .IN3(N2578), .IN4(n3373), .IN5(
        n3349), .IN6(EBX_30_), .Q(n2795) );
  NOR2X0 U3386 ( .IN1(n3355), .IN2(n4120), .QN(n4119) );
  NOR2X0 U3387 ( .IN1(n4121), .IN2(n3349), .QN(n4118) );
  AO21X1 U3388 ( .IN1(n4122), .IN2(n4121), .IN3(n4091), .Q(n4117) );
  OR2X1 U3389 ( .IN1(n4120), .IN2(n4123), .Q(n4122) );
  NAND4X0 U3390 ( .IN1(n4124), .IN2(n4125), .IN3(n4126), .IN4(n4127), .QN(
        n4121) );
  NOR2X0 U3391 ( .IN1(n4128), .IN2(n4129), .QN(n4127) );
  MUX21X1 U3392 ( .IN1(n2870), .IN2(n4130), .S(n4131), .Q(n2794) );
  INVX0 U3393 ( .IN(n4106), .QN(n4130) );
  MUX21X1 U3394 ( .IN1(n4132), .IN2(N2737), .S(n4079), .Q(n2793) );
  AO222X1 U3395 ( .IN1(n4081), .IN2(n1552), .IN3(n1557), .IN4(n4133), .IN5(
        n4017), .IN6(n4134), .Q(n4132) );
  MUX21X1 U3396 ( .IN1(n4135), .IN2(InstQueueRd_Addr[1]), .S(n4079), .Q(n2792)
         );
  AO222X1 U3397 ( .IN1(n4081), .IN2(n4136), .IN3(n4137), .IN4(n4133), .IN5(
        n4017), .IN6(n4138), .Q(n4135) );
  MUX21X1 U3398 ( .IN1(n4139), .IN2(n4140), .S(n4079), .Q(n2791) );
  AO222X1 U3399 ( .IN1(n4141), .IN2(n4081), .IN3(n4142), .IN4(n4143), .IN5(
        n4017), .IN6(n4144), .Q(n4139) );
  NOR2X0 U3400 ( .IN1(n1557), .IN2(n4088), .QN(n4142) );
  MUX21X1 U3401 ( .IN1(n4145), .IN2(InstQueueRd_Addr[4]), .S(n4079), .Q(n2790)
         );
  AND3X1 U3402 ( .IN1(n4095), .IN2(n4146), .IN3(n4147), .Q(n4079) );
  NOR3X0 U3403 ( .IN1(n2883), .IN2(n4091), .IN3(n4148), .QN(n4145) );
  AO22X1 U3404 ( .IN1(n4149), .IN2(N1239), .IN3(n4150), .IN4(n4151), .Q(n2789)
         );
  OAI21X1 U3405 ( .IN1(n4088), .IN2(N3494), .IN3(n4152), .QN(n4150) );
  NAND2X0 U3406 ( .IN1(n4103), .IN2(n4151), .QN(n4149) );
  MUX21X1 U3407 ( .IN1(n4153), .IN2(n4154), .S(n1555), .Q(n2788) );
  OA21X1 U3408 ( .IN1(n4155), .IN2(n3388), .IN3(n4151), .Q(n4154) );
  NOR2X0 U3409 ( .IN1(n1556), .IN2(n4095), .QN(n4155) );
  NAND3X0 U3410 ( .IN1(n4151), .IN2(n3396), .IN3(n4152), .QN(n4153) );
  AO22X1 U3411 ( .IN1(n4157), .IN2(N3990), .IN3(n4158), .IN4(n4151), .Q(n2787)
         );
  AO222X1 U3412 ( .IN1(n4159), .IN2(n4089), .IN3(n4160), .IN4(n1554), .IN5(
        n4161), .IN6(n4162), .Q(n4158) );
  MUX21X1 U3413 ( .IN1(n4163), .IN2(n3391), .S(n4165), .Q(n4160) );
  NAND3X0 U3414 ( .IN1(n4166), .IN2(n4151), .IN3(n4167), .QN(n4157) );
  INVX0 U3415 ( .IN(n4168), .QN(n4167) );
  NAND2X0 U3416 ( .IN1(n4163), .IN2(n4165), .QN(n4166) );
  OAI22X1 U3417 ( .IN1(n1553), .IN2(n4169), .IN3(n4170), .IN4(n4171), .QN(
        n2786) );
  OA22X1 U3418 ( .IN1(n4172), .IN2(N3989), .IN3(n4095), .IN4(n4173), .Q(n4171)
         );
  OA22X1 U3419 ( .IN1(n4174), .IN2(n4175), .IN3(n4090), .IN4(n4176), .Q(n4172)
         );
  NOR4X0 U3420 ( .IN1(n4170), .IN2(n4177), .IN3(n4178), .IN4(n4168), .QN(n4169) );
  NAND2X0 U3421 ( .IN1(n4179), .IN2(n4152), .QN(n4168) );
  NAND2X0 U3422 ( .IN1(n1556), .IN2(n4089), .QN(n4152) );
  AO21X1 U3423 ( .IN1(n4095), .IN2(n4090), .IN3(N3991), .Q(n4179) );
  ISOLANDX1 U3424 ( .D(n4175), .ISO(n4174), .Q(n4178) );
  AO21X1 U3425 ( .IN1(n1472), .IN2(n4165), .IN3(n1554), .Q(n4175) );
  NAND2X0 U3426 ( .IN1(n1472), .IN2(N3991), .QN(n4165) );
  OA21X1 U3427 ( .IN1(n4089), .IN2(n4161), .IN3(n1554), .Q(n4177) );
  INVX0 U3428 ( .IN(n4151), .QN(n4170) );
  NAND3X0 U3429 ( .IN1(n4180), .IN2(n4147), .IN3(n4181), .QN(n4151) );
  NAND2X0 U3430 ( .IN1(n4133), .IN2(n2870), .QN(n4147) );
  NAND2X0 U3431 ( .IN1(N3494), .IN2(n4133), .QN(n4180) );
  INVX0 U3432 ( .IN(n4088), .QN(n4133) );
  NAND3X0 U3433 ( .IN1(n2865), .IN2(n2844), .IN3(n4116), .QN(n4088) );
  AO221X1 U3434 ( .IN1(n3080), .IN2(n4182), .IN3(n3101), .IN4(n4183), .IN5(
        n4184), .Q(n2785) );
  AO21X1 U3435 ( .IN1(n4185), .IN2(n4186), .IN3(n4187), .Q(n4184) );
  MUX21X1 U3436 ( .IN1(N2548), .IN2(n4188), .S(n4189), .Q(n4187) );
  AO221X1 U3437 ( .IN1(n3082), .IN2(n4182), .IN3(n3100), .IN4(n4183), .IN5(
        n4190), .Q(n2784) );
  AO21X1 U3438 ( .IN1(n4191), .IN2(n4186), .IN3(n4192), .Q(n4190) );
  MUX21X1 U3439 ( .IN1(N2549), .IN2(n4193), .S(n4189), .Q(n4192) );
  AO221X1 U3440 ( .IN1(n3084), .IN2(n4182), .IN3(n3099), .IN4(n4183), .IN5(
        n4194), .Q(n2783) );
  AO21X1 U3441 ( .IN1(n4195), .IN2(n4186), .IN3(n4196), .Q(n4194) );
  MUX21X1 U3442 ( .IN1(N2550), .IN2(n4197), .S(n4189), .Q(n4196) );
  AO221X1 U3443 ( .IN1(n3086), .IN2(n4182), .IN3(n3098), .IN4(n4183), .IN5(
        n4198), .Q(n2782) );
  AO21X1 U3444 ( .IN1(n4199), .IN2(n4186), .IN3(n4200), .Q(n4198) );
  MUX21X1 U3445 ( .IN1(N2551), .IN2(n4201), .S(n4189), .Q(n4200) );
  AO221X1 U3446 ( .IN1(n3088), .IN2(n4182), .IN3(n3097), .IN4(n4183), .IN5(
        n4202), .Q(n2781) );
  AO21X1 U3447 ( .IN1(n4203), .IN2(n4186), .IN3(n4204), .Q(n4202) );
  MUX21X1 U3448 ( .IN1(n4205), .IN2(N2552), .S(n4206), .Q(n4204) );
  AO221X1 U3449 ( .IN1(n3090), .IN2(n4182), .IN3(n3096), .IN4(n4183), .IN5(
        n4207), .Q(n2780) );
  AO21X1 U3450 ( .IN1(n4208), .IN2(n4186), .IN3(n4209), .Q(n4207) );
  MUX21X1 U3451 ( .IN1(n4210), .IN2(N2553), .S(n4206), .Q(n4209) );
  AO221X1 U3452 ( .IN1(n3092), .IN2(n4182), .IN3(n3095), .IN4(n4183), .IN5(
        n4211), .Q(n2779) );
  AO21X1 U3453 ( .IN1(n4212), .IN2(n4186), .IN3(n4213), .Q(n4211) );
  MUX21X1 U3454 ( .IN1(n4214), .IN2(N2554), .S(n4206), .Q(n4213) );
  AO221X1 U3455 ( .IN1(n3094), .IN2(n4182), .IN3(n2843), .IN4(n4183), .IN5(
        n4215), .Q(n2778) );
  AO21X1 U3456 ( .IN1(n4216), .IN2(n4186), .IN3(n4217), .Q(n4215) );
  MUX21X1 U3457 ( .IN1(n4218), .IN2(N2555), .S(n4206), .Q(n4217) );
  NOR4X0 U3458 ( .IN1(n4174), .IN2(n4206), .IN3(n4186), .IN4(n4219), .QN(n4182) );
  INVX0 U3459 ( .IN(n4189), .QN(n4206) );
  AO221X1 U3460 ( .IN1(n4220), .IN2(n4221), .IN3(n4222), .IN4(n4012), .IN5(
        n4223), .Q(n4189) );
  NAND2X0 U3461 ( .IN1(n4224), .IN2(n4225), .QN(n4223) );
  AO221X1 U3462 ( .IN1(n4226), .IN2(n3080), .IN3(n4227), .IN4(n3101), .IN5(
        n4228), .Q(n2777) );
  AO21X1 U3463 ( .IN1(n4185), .IN2(n4219), .IN3(n4229), .Q(n4228) );
  MUX21X1 U3464 ( .IN1(n4188), .IN2(test_so9), .S(n4231), .Q(n4229) );
  AO221X1 U3465 ( .IN1(n4226), .IN2(n3082), .IN3(n4227), .IN4(n3100), .IN5(
        n4232), .Q(n2776) );
  AO21X1 U3466 ( .IN1(n4191), .IN2(n4219), .IN3(n4233), .Q(n4232) );
  MUX21X1 U3467 ( .IN1(n4234), .IN2(n4193), .S(n4235), .Q(n4233) );
  AO221X1 U3468 ( .IN1(n4226), .IN2(n3084), .IN3(n4227), .IN4(n3099), .IN5(
        n4236), .Q(n2775) );
  AO21X1 U3469 ( .IN1(n4195), .IN2(n4219), .IN3(n4237), .Q(n4236) );
  MUX21X1 U3470 ( .IN1(n4238), .IN2(n4197), .S(n4235), .Q(n4237) );
  AO221X1 U3471 ( .IN1(n4226), .IN2(n3086), .IN3(n4227), .IN4(n3098), .IN5(
        n4239), .Q(n2774) );
  AO21X1 U3472 ( .IN1(n4199), .IN2(n4219), .IN3(n4240), .Q(n4239) );
  MUX21X1 U3473 ( .IN1(n4241), .IN2(n4201), .S(n4235), .Q(n4240) );
  AO221X1 U3474 ( .IN1(n4226), .IN2(n3088), .IN3(n4227), .IN4(n3097), .IN5(
        n4242), .Q(n2773) );
  AO21X1 U3475 ( .IN1(n4203), .IN2(n4219), .IN3(n4243), .Q(n4242) );
  MUX21X1 U3476 ( .IN1(n4205), .IN2(n4244), .S(n4231), .Q(n4243) );
  AO221X1 U3477 ( .IN1(n4226), .IN2(n3090), .IN3(n4227), .IN4(n3096), .IN5(
        n4245), .Q(n2772) );
  AO21X1 U3478 ( .IN1(n4208), .IN2(n4219), .IN3(n4246), .Q(n4245) );
  MUX21X1 U3479 ( .IN1(n4210), .IN2(n4247), .S(n4231), .Q(n4246) );
  AO221X1 U3480 ( .IN1(n4226), .IN2(n3092), .IN3(n4227), .IN4(n3095), .IN5(
        n4248), .Q(n2771) );
  AO21X1 U3481 ( .IN1(n4212), .IN2(n4219), .IN3(n4249), .Q(n4248) );
  MUX21X1 U3482 ( .IN1(n4214), .IN2(n4250), .S(n4231), .Q(n4249) );
  AO221X1 U3483 ( .IN1(n4226), .IN2(n3094), .IN3(n4227), .IN4(n2843), .IN5(
        n4251), .Q(n2770) );
  AO21X1 U3484 ( .IN1(n4216), .IN2(n4219), .IN3(n4252), .Q(n4251) );
  MUX21X1 U3485 ( .IN1(n4218), .IN2(n4253), .S(n4231), .Q(n4252) );
  INVX0 U3486 ( .IN(n4235), .QN(n4231) );
  AND4X1 U3487 ( .IN1(n4254), .IN2(n4235), .IN3(n4255), .IN4(n4256), .Q(n4226)
         );
  AO221X1 U3488 ( .IN1(n4220), .IN2(n4012), .IN3(n4257), .IN4(n4221), .IN5(
        n4258), .Q(n4235) );
  NAND2X0 U3489 ( .IN1(n4259), .IN2(n4225), .QN(n4258) );
  INVX0 U3490 ( .IN(n4183), .QN(n4225) );
  AO221X1 U3491 ( .IN1(n4260), .IN2(n3080), .IN3(n4261), .IN4(n3101), .IN5(
        n4262), .Q(n2769) );
  AO21X1 U3492 ( .IN1(n4185), .IN2(n4222), .IN3(n4263), .Q(n4262) );
  MUX21X1 U3493 ( .IN1(n2848), .IN2(n4188), .S(n4264), .Q(n4263) );
  AO221X1 U3494 ( .IN1(n4260), .IN2(n3082), .IN3(n4261), .IN4(n3100), .IN5(
        n4265), .Q(n2768) );
  AO21X1 U3495 ( .IN1(n4191), .IN2(n4222), .IN3(n4266), .Q(n4265) );
  MUX21X1 U3496 ( .IN1(n2861), .IN2(n4193), .S(n4264), .Q(n4266) );
  AO221X1 U3497 ( .IN1(n4260), .IN2(n3084), .IN3(n4261), .IN4(n3099), .IN5(
        n4267), .Q(n2767) );
  AO21X1 U3498 ( .IN1(n4195), .IN2(n4222), .IN3(n4268), .Q(n4267) );
  MUX21X1 U3499 ( .IN1(n2862), .IN2(n4197), .S(n4264), .Q(n4268) );
  AO221X1 U3500 ( .IN1(n4260), .IN2(n3086), .IN3(n4261), .IN4(n3098), .IN5(
        n4269), .Q(n2766) );
  AO21X1 U3501 ( .IN1(n4199), .IN2(n4222), .IN3(n4270), .Q(n4269) );
  MUX21X1 U3502 ( .IN1(n2863), .IN2(n4201), .S(n4264), .Q(n4270) );
  AO221X1 U3503 ( .IN1(n4260), .IN2(n3088), .IN3(n4261), .IN4(n3097), .IN5(
        n4271), .Q(n2765) );
  AO21X1 U3504 ( .IN1(n4203), .IN2(n4222), .IN3(n4272), .Q(n4271) );
  MUX21X1 U3505 ( .IN1(n4205), .IN2(n2857), .S(n4273), .Q(n4272) );
  AO221X1 U3506 ( .IN1(n4260), .IN2(n3090), .IN3(n4261), .IN4(n3096), .IN5(
        n4274), .Q(n2764) );
  AO21X1 U3507 ( .IN1(n4208), .IN2(n4222), .IN3(n4275), .Q(n4274) );
  MUX21X1 U3508 ( .IN1(n4210), .IN2(n2858), .S(n4273), .Q(n4275) );
  AO221X1 U3509 ( .IN1(n4260), .IN2(n3092), .IN3(n4261), .IN4(n3095), .IN5(
        n4276), .Q(n2763) );
  AO21X1 U3510 ( .IN1(n4212), .IN2(n4222), .IN3(n4277), .Q(n4276) );
  MUX21X1 U3511 ( .IN1(n4214), .IN2(n2859), .S(n4273), .Q(n4277) );
  AO221X1 U3512 ( .IN1(n4260), .IN2(n3094), .IN3(n4261), .IN4(n2843), .IN5(
        n4278), .Q(n2762) );
  AO21X1 U3513 ( .IN1(n4216), .IN2(n4222), .IN3(n4279), .Q(n4278) );
  MUX21X1 U3514 ( .IN1(n4218), .IN2(n2860), .S(n4273), .Q(n4279) );
  NOR4X0 U3515 ( .IN1(n4174), .IN2(n4273), .IN3(n4220), .IN4(n4222), .QN(n4260) );
  INVX0 U3516 ( .IN(n4264), .QN(n4273) );
  AO221X1 U3517 ( .IN1(n4257), .IN2(n4012), .IN3(n4280), .IN4(n4221), .IN5(
        n4281), .Q(n4264) );
  NAND2X0 U3518 ( .IN1(n4282), .IN2(n4259), .QN(n4281) );
  INVX0 U3519 ( .IN(n4227), .QN(n4259) );
  AO221X1 U3520 ( .IN1(n4283), .IN2(n3080), .IN3(n4185), .IN4(n4220), .IN5(
        n4284), .Q(n2761) );
  AO21X1 U3521 ( .IN1(n4285), .IN2(n3101), .IN3(n4286), .Q(n4284) );
  MUX21X1 U3522 ( .IN1(n4188), .IN2(n2916), .S(n4287), .Q(n4286) );
  AO221X1 U3523 ( .IN1(n4283), .IN2(n3082), .IN3(n4191), .IN4(n4220), .IN5(
        n4288), .Q(n2760) );
  AO21X1 U3524 ( .IN1(n4285), .IN2(n3100), .IN3(n4289), .Q(n4288) );
  MUX21X1 U3525 ( .IN1(n2931), .IN2(n4193), .S(n4290), .Q(n4289) );
  AO221X1 U3526 ( .IN1(n4283), .IN2(n3084), .IN3(n4195), .IN4(n4220), .IN5(
        n4291), .Q(n2759) );
  AO21X1 U3527 ( .IN1(n4285), .IN2(n3099), .IN3(n4292), .Q(n4291) );
  MUX21X1 U3528 ( .IN1(n2932), .IN2(n4197), .S(n4290), .Q(n4292) );
  AO221X1 U3529 ( .IN1(n4283), .IN2(n3086), .IN3(n4199), .IN4(n4220), .IN5(
        n4293), .Q(n2758) );
  AO21X1 U3530 ( .IN1(n4285), .IN2(n3098), .IN3(n4294), .Q(n4293) );
  MUX21X1 U3531 ( .IN1(n2933), .IN2(n4201), .S(n4290), .Q(n4294) );
  AO221X1 U3532 ( .IN1(n4283), .IN2(n3088), .IN3(n4203), .IN4(n4220), .IN5(
        n4295), .Q(n2757) );
  AO21X1 U3533 ( .IN1(n4285), .IN2(n3097), .IN3(n4296), .Q(n4295) );
  MUX21X1 U3534 ( .IN1(n4205), .IN2(n2917), .S(n4287), .Q(n4296) );
  AO221X1 U3535 ( .IN1(n4283), .IN2(n3090), .IN3(n4208), .IN4(n4220), .IN5(
        n4297), .Q(n2756) );
  AO21X1 U3536 ( .IN1(n4285), .IN2(n3096), .IN3(n4298), .Q(n4297) );
  MUX21X1 U3537 ( .IN1(n4210), .IN2(test_so10), .S(n4287), .Q(n4298) );
  AO221X1 U3538 ( .IN1(n4283), .IN2(n3092), .IN3(n4212), .IN4(n4220), .IN5(
        n4299), .Q(n2755) );
  AO21X1 U3539 ( .IN1(n4285), .IN2(n3095), .IN3(n4300), .Q(n4299) );
  MUX21X1 U3540 ( .IN1(n4214), .IN2(n2919), .S(n4287), .Q(n4300) );
  AO221X1 U3541 ( .IN1(n4283), .IN2(n3094), .IN3(n4216), .IN4(n4220), .IN5(
        n4301), .Q(n2754) );
  AO21X1 U3542 ( .IN1(n4285), .IN2(n2843), .IN3(n4302), .Q(n4301) );
  MUX21X1 U3543 ( .IN1(n4218), .IN2(n2920), .S(n4287), .Q(n4302) );
  INVX0 U3544 ( .IN(n4290), .QN(n4287) );
  AND4X1 U3545 ( .IN1(n4254), .IN2(n4290), .IN3(n4303), .IN4(n4304), .Q(n4283)
         );
  AO221X1 U3546 ( .IN1(n4280), .IN2(n4012), .IN3(n4305), .IN4(n4221), .IN5(
        n4306), .Q(n4290) );
  NAND2X0 U3547 ( .IN1(n4307), .IN2(n4282), .QN(n4306) );
  INVX0 U3548 ( .IN(n4261), .QN(n4282) );
  NAND3X0 U3549 ( .IN1(n1553), .IN2(n1554), .IN3(n4308), .QN(n4303) );
  AO221X1 U3550 ( .IN1(n4309), .IN2(n3080), .IN3(n4257), .IN4(n4185), .IN5(
        n4310), .Q(n2753) );
  AO21X1 U3551 ( .IN1(n4311), .IN2(n3101), .IN3(n4312), .Q(n4310) );
  MUX21X1 U3552 ( .IN1(n4313), .IN2(n4188), .S(n4314), .Q(n4312) );
  AO221X1 U3553 ( .IN1(n4309), .IN2(n3082), .IN3(n4257), .IN4(n4191), .IN5(
        n4315), .Q(n2752) );
  AO21X1 U3554 ( .IN1(n4311), .IN2(n3100), .IN3(n4316), .Q(n4315) );
  MUX21X1 U3555 ( .IN1(n4317), .IN2(n4193), .S(n4314), .Q(n4316) );
  AO221X1 U3556 ( .IN1(n4309), .IN2(n3084), .IN3(n4257), .IN4(n4195), .IN5(
        n4318), .Q(n2751) );
  AO21X1 U3557 ( .IN1(n4311), .IN2(n3099), .IN3(n4319), .Q(n4318) );
  MUX21X1 U3558 ( .IN1(n4320), .IN2(n4197), .S(n4314), .Q(n4319) );
  AO221X1 U3559 ( .IN1(n4309), .IN2(n3086), .IN3(n4257), .IN4(n4199), .IN5(
        n4321), .Q(n2750) );
  AO21X1 U3560 ( .IN1(n4311), .IN2(n3098), .IN3(n4322), .Q(n4321) );
  MUX21X1 U3561 ( .IN1(n4323), .IN2(n4201), .S(n4314), .Q(n4322) );
  AO221X1 U3562 ( .IN1(n4309), .IN2(n3088), .IN3(n4257), .IN4(n4203), .IN5(
        n4324), .Q(n2749) );
  AO21X1 U3563 ( .IN1(n4311), .IN2(n3097), .IN3(n4325), .Q(n4324) );
  MUX21X1 U3564 ( .IN1(n4205), .IN2(n4326), .S(n4327), .Q(n4325) );
  AO221X1 U3565 ( .IN1(n4309), .IN2(n3090), .IN3(n4257), .IN4(n4208), .IN5(
        n4328), .Q(n2748) );
  AO21X1 U3566 ( .IN1(n4311), .IN2(n3096), .IN3(n4329), .Q(n4328) );
  MUX21X1 U3567 ( .IN1(n4210), .IN2(n4330), .S(n4327), .Q(n4329) );
  AO221X1 U3568 ( .IN1(n4309), .IN2(n3092), .IN3(n4257), .IN4(n4212), .IN5(
        n4331), .Q(n2747) );
  AO21X1 U3569 ( .IN1(n4311), .IN2(n3095), .IN3(n4332), .Q(n4331) );
  MUX21X1 U3570 ( .IN1(n4214), .IN2(n4333), .S(n4327), .Q(n4332) );
  AO221X1 U3571 ( .IN1(n4309), .IN2(n3094), .IN3(n4257), .IN4(n4216), .IN5(
        n4334), .Q(n2746) );
  AO21X1 U3572 ( .IN1(n4311), .IN2(n2843), .IN3(n4335), .Q(n4334) );
  MUX21X1 U3573 ( .IN1(n4218), .IN2(n4336), .S(n4327), .Q(n4335) );
  NOR4X0 U3574 ( .IN1(n4174), .IN2(n4327), .IN3(n4257), .IN4(n4280), .QN(n4309) );
  INVX0 U3575 ( .IN(n4314), .QN(n4327) );
  AO221X1 U3576 ( .IN1(n4305), .IN2(n4012), .IN3(n4337), .IN4(n4221), .IN5(
        n4338), .Q(n4314) );
  NAND2X0 U3577 ( .IN1(n4339), .IN2(n4307), .QN(n4338) );
  INVX0 U3578 ( .IN(n4285), .QN(n4307) );
  NAND3X0 U3579 ( .IN1(n1553), .IN2(n1554), .IN3(n4340), .QN(n4304) );
  AO221X1 U3580 ( .IN1(n4341), .IN2(n3080), .IN3(n4280), .IN4(n4185), .IN5(
        n4342), .Q(n2745) );
  AO21X1 U3581 ( .IN1(n4343), .IN2(n3101), .IN3(n4344), .Q(n4342) );
  MUX21X1 U3582 ( .IN1(n4345), .IN2(n4188), .S(n4346), .Q(n4344) );
  AO221X1 U3583 ( .IN1(n4341), .IN2(n3082), .IN3(n4280), .IN4(n4191), .IN5(
        n4347), .Q(n2744) );
  AO21X1 U3584 ( .IN1(n4343), .IN2(n3100), .IN3(n4348), .Q(n4347) );
  MUX21X1 U3585 ( .IN1(n4349), .IN2(n4193), .S(n4346), .Q(n4348) );
  AO221X1 U3586 ( .IN1(n4341), .IN2(n3084), .IN3(n4280), .IN4(n4195), .IN5(
        n4350), .Q(n2743) );
  AO21X1 U3587 ( .IN1(n4343), .IN2(n3099), .IN3(n4351), .Q(n4350) );
  MUX21X1 U3588 ( .IN1(n4352), .IN2(n4197), .S(n4346), .Q(n4351) );
  AO221X1 U3589 ( .IN1(n4341), .IN2(n3086), .IN3(n4280), .IN4(n4199), .IN5(
        n4353), .Q(n2742) );
  AO21X1 U3590 ( .IN1(n4343), .IN2(n3098), .IN3(n4354), .Q(n4353) );
  MUX21X1 U3591 ( .IN1(n4201), .IN2(n4355), .S(n4356), .Q(n4354) );
  AO221X1 U3592 ( .IN1(n4341), .IN2(n3088), .IN3(n4280), .IN4(n4203), .IN5(
        n4357), .Q(n2741) );
  AO21X1 U3593 ( .IN1(n4343), .IN2(n3097), .IN3(n4358), .Q(n4357) );
  MUX21X1 U3594 ( .IN1(n4205), .IN2(n4359), .S(n4356), .Q(n4358) );
  AO221X1 U3595 ( .IN1(n4341), .IN2(n3090), .IN3(n4280), .IN4(n4208), .IN5(
        n4360), .Q(n2740) );
  AO21X1 U3596 ( .IN1(n4343), .IN2(n3096), .IN3(n4361), .Q(n4360) );
  MUX21X1 U3597 ( .IN1(n4210), .IN2(n4362), .S(n4356), .Q(n4361) );
  AO221X1 U3598 ( .IN1(n4341), .IN2(n3092), .IN3(n4280), .IN4(n4212), .IN5(
        n4363), .Q(n2739) );
  AO21X1 U3599 ( .IN1(n4343), .IN2(n3095), .IN3(n4364), .Q(n4363) );
  MUX21X1 U3600 ( .IN1(n4214), .IN2(n4365), .S(n4356), .Q(n4364) );
  AO221X1 U3601 ( .IN1(n4341), .IN2(n3094), .IN3(n4280), .IN4(n4216), .IN5(
        n4366), .Q(n2738) );
  AO21X1 U3602 ( .IN1(n4343), .IN2(n2843), .IN3(n4367), .Q(n4366) );
  MUX21X1 U3603 ( .IN1(n4218), .IN2(n4368), .S(n4356), .Q(n4367) );
  INVX0 U3604 ( .IN(n4346), .QN(n4356) );
  AND4X1 U3605 ( .IN1(n4254), .IN2(n4346), .IN3(n4369), .IN4(n4370), .Q(n4341)
         );
  AO221X1 U3606 ( .IN1(n4337), .IN2(n4012), .IN3(n4371), .IN4(n4221), .IN5(
        n4372), .Q(n4346) );
  NAND2X0 U3607 ( .IN1(n4373), .IN2(n4339), .QN(n4372) );
  INVX0 U3608 ( .IN(n4311), .QN(n4339) );
  NAND3X0 U3609 ( .IN1(n4162), .IN2(n1556), .IN3(n1553), .QN(n4369) );
  AO221X1 U3610 ( .IN1(n4374), .IN2(n3080), .IN3(n4305), .IN4(n4185), .IN5(
        n4375), .Q(n2737) );
  AO21X1 U3611 ( .IN1(n4376), .IN2(n3101), .IN3(n4377), .Q(n4375) );
  MUX21X1 U3612 ( .IN1(n2869), .IN2(n4188), .S(n4378), .Q(n4377) );
  AO221X1 U3613 ( .IN1(n4374), .IN2(n3082), .IN3(n4305), .IN4(n4191), .IN5(
        n4379), .Q(n2736) );
  AO21X1 U3614 ( .IN1(n4376), .IN2(n3100), .IN3(n4380), .Q(n4379) );
  MUX21X1 U3615 ( .IN1(n2884), .IN2(n4193), .S(n4378), .Q(n4380) );
  AO221X1 U3616 ( .IN1(n4374), .IN2(n3084), .IN3(n4305), .IN4(n4195), .IN5(
        n4381), .Q(n2735) );
  AO21X1 U3617 ( .IN1(n4376), .IN2(n3099), .IN3(n4382), .Q(n4381) );
  MUX21X1 U3618 ( .IN1(test_so11), .IN2(n4197), .S(n4378), .Q(n4382) );
  AO221X1 U3619 ( .IN1(n4374), .IN2(n3086), .IN3(n4305), .IN4(n4199), .IN5(
        n4383), .Q(n2734) );
  AO21X1 U3620 ( .IN1(n4376), .IN2(n3098), .IN3(n4384), .Q(n4383) );
  MUX21X1 U3621 ( .IN1(n2886), .IN2(n4201), .S(n4378), .Q(n4384) );
  AO221X1 U3622 ( .IN1(n4374), .IN2(n3088), .IN3(n4305), .IN4(n4203), .IN5(
        n4385), .Q(n2733) );
  AO21X1 U3623 ( .IN1(n4376), .IN2(n3097), .IN3(n4386), .Q(n4385) );
  MUX21X1 U3624 ( .IN1(n4205), .IN2(n2879), .S(n4387), .Q(n4386) );
  AO221X1 U3625 ( .IN1(n4374), .IN2(n3090), .IN3(n4305), .IN4(n4208), .IN5(
        n4388), .Q(n2732) );
  AO21X1 U3626 ( .IN1(n4376), .IN2(n3096), .IN3(n4389), .Q(n4388) );
  MUX21X1 U3627 ( .IN1(n4210), .IN2(n2880), .S(n4387), .Q(n4389) );
  AO221X1 U3628 ( .IN1(n4374), .IN2(n3092), .IN3(n4305), .IN4(n4212), .IN5(
        n4390), .Q(n2731) );
  AO21X1 U3629 ( .IN1(n4376), .IN2(n3095), .IN3(n4391), .Q(n4390) );
  MUX21X1 U3630 ( .IN1(n4214), .IN2(n2881), .S(n4387), .Q(n4391) );
  AO221X1 U3631 ( .IN1(n4374), .IN2(n3094), .IN3(n4305), .IN4(n4216), .IN5(
        n4392), .Q(n2730) );
  AO21X1 U3632 ( .IN1(n4376), .IN2(n2843), .IN3(n4393), .Q(n4392) );
  MUX21X1 U3633 ( .IN1(n4218), .IN2(n2882), .S(n4387), .Q(n4393) );
  NOR4X0 U3634 ( .IN1(n4174), .IN2(n4387), .IN3(n4305), .IN4(n4337), .QN(n4374) );
  INVX0 U3635 ( .IN(n4378), .QN(n4387) );
  AO221X1 U3636 ( .IN1(n4371), .IN2(n4012), .IN3(n4394), .IN4(n4221), .IN5(
        n4395), .Q(n4378) );
  NAND2X0 U3637 ( .IN1(n4396), .IN2(n4373), .QN(n4395) );
  INVX0 U3638 ( .IN(n4343), .QN(n4373) );
  NAND2X0 U3639 ( .IN1(n1553), .IN2(n4159), .QN(n4370) );
  AO221X1 U3640 ( .IN1(n4397), .IN2(n3080), .IN3(n4337), .IN4(n4185), .IN5(
        n4398), .Q(n2729) );
  AO21X1 U3641 ( .IN1(n4399), .IN2(n3101), .IN3(n4400), .Q(n4398) );
  MUX21X1 U3642 ( .IN1(n2921), .IN2(n4188), .S(n4401), .Q(n4400) );
  AO221X1 U3643 ( .IN1(n4397), .IN2(n3082), .IN3(n4337), .IN4(n4191), .IN5(
        n4402), .Q(n2728) );
  AO21X1 U3644 ( .IN1(n4399), .IN2(n3100), .IN3(n4403), .Q(n4402) );
  MUX21X1 U3645 ( .IN1(n2922), .IN2(n4193), .S(n4401), .Q(n4403) );
  AO221X1 U3646 ( .IN1(n4397), .IN2(n3084), .IN3(n4337), .IN4(n4195), .IN5(
        n4404), .Q(n2727) );
  AO21X1 U3647 ( .IN1(n4399), .IN2(n3099), .IN3(n4405), .Q(n4404) );
  MUX21X1 U3648 ( .IN1(n2923), .IN2(n4197), .S(n4401), .Q(n4405) );
  AO221X1 U3649 ( .IN1(n4397), .IN2(n3086), .IN3(n4337), .IN4(n4199), .IN5(
        n4406), .Q(n2726) );
  AO21X1 U3650 ( .IN1(n4399), .IN2(n3098), .IN3(n4407), .Q(n4406) );
  MUX21X1 U3651 ( .IN1(n4201), .IN2(n2902), .S(n4408), .Q(n4407) );
  AO221X1 U3652 ( .IN1(n4397), .IN2(n3088), .IN3(n4337), .IN4(n4203), .IN5(
        n4409), .Q(n2725) );
  AO21X1 U3653 ( .IN1(n4399), .IN2(n3097), .IN3(n4410), .Q(n4409) );
  MUX21X1 U3654 ( .IN1(n4205), .IN2(n2903), .S(n4408), .Q(n4410) );
  AO221X1 U3655 ( .IN1(n4397), .IN2(n3090), .IN3(n4337), .IN4(n4208), .IN5(
        n4411), .Q(n2724) );
  AO21X1 U3656 ( .IN1(n4399), .IN2(n3096), .IN3(n4412), .Q(n4411) );
  MUX21X1 U3657 ( .IN1(n4210), .IN2(n2904), .S(n4408), .Q(n4412) );
  AO221X1 U3658 ( .IN1(n4397), .IN2(n3092), .IN3(n4337), .IN4(n4212), .IN5(
        n4413), .Q(n2723) );
  AO21X1 U3659 ( .IN1(n4399), .IN2(n3095), .IN3(n4414), .Q(n4413) );
  MUX21X1 U3660 ( .IN1(n4214), .IN2(n2905), .S(n4408), .Q(n4414) );
  AO221X1 U3661 ( .IN1(n4397), .IN2(n3094), .IN3(n4337), .IN4(n4216), .IN5(
        n4415), .Q(n2722) );
  AO21X1 U3662 ( .IN1(n4399), .IN2(n2843), .IN3(n4416), .Q(n4415) );
  MUX21X1 U3663 ( .IN1(n4218), .IN2(n2906), .S(n4408), .Q(n4416) );
  INVX0 U3664 ( .IN(n4401), .QN(n4408) );
  AND4X1 U3665 ( .IN1(n4254), .IN2(n4401), .IN3(n4417), .IN4(n4418), .Q(n4397)
         );
  AO221X1 U3666 ( .IN1(n4394), .IN2(n4012), .IN3(n4419), .IN4(n4221), .IN5(
        n4420), .Q(n4401) );
  NAND2X0 U3667 ( .IN1(n4421), .IN2(n4396), .QN(n4420) );
  INVX0 U3668 ( .IN(n4376), .QN(n4396) );
  NAND3X0 U3669 ( .IN1(n1553), .IN2(N3990), .IN3(n4308), .QN(n4417) );
  AO221X1 U3670 ( .IN1(n4422), .IN2(n3080), .IN3(n4371), .IN4(n4185), .IN5(
        n4423), .Q(n2721) );
  AO21X1 U3671 ( .IN1(n4424), .IN2(n3101), .IN3(n4425), .Q(n4423) );
  MUX21X1 U3672 ( .IN1(n4426), .IN2(n4188), .S(n4427), .Q(n4425) );
  AO221X1 U3673 ( .IN1(n4422), .IN2(n3082), .IN3(n4371), .IN4(n4191), .IN5(
        n4428), .Q(n2720) );
  AO21X1 U3674 ( .IN1(n4424), .IN2(n3100), .IN3(n4429), .Q(n4428) );
  MUX21X1 U3675 ( .IN1(n4430), .IN2(n4193), .S(n4427), .Q(n4429) );
  AO221X1 U3676 ( .IN1(n4422), .IN2(n3084), .IN3(n4371), .IN4(n4195), .IN5(
        n4431), .Q(n2719) );
  AO21X1 U3677 ( .IN1(n4424), .IN2(n3099), .IN3(n4432), .Q(n4431) );
  MUX21X1 U3678 ( .IN1(n4433), .IN2(n4197), .S(n4427), .Q(n4432) );
  AO221X1 U3679 ( .IN1(n4422), .IN2(n3086), .IN3(n4371), .IN4(n4199), .IN5(
        n4434), .Q(n2718) );
  AO21X1 U3680 ( .IN1(n4424), .IN2(n3098), .IN3(n4435), .Q(n4434) );
  MUX21X1 U3681 ( .IN1(n4436), .IN2(n4201), .S(n4427), .Q(n4435) );
  AO221X1 U3682 ( .IN1(n4422), .IN2(n3088), .IN3(n4371), .IN4(n4203), .IN5(
        n4437), .Q(n2717) );
  AO21X1 U3683 ( .IN1(n4424), .IN2(n3097), .IN3(n4438), .Q(n4437) );
  MUX21X1 U3684 ( .IN1(n4205), .IN2(n4439), .S(n4440), .Q(n4438) );
  AO221X1 U3685 ( .IN1(n4422), .IN2(n3090), .IN3(n4371), .IN4(n4208), .IN5(
        n4441), .Q(n2716) );
  AO21X1 U3686 ( .IN1(n4424), .IN2(n3096), .IN3(n4442), .Q(n4441) );
  MUX21X1 U3687 ( .IN1(n4210), .IN2(n4443), .S(n4440), .Q(n4442) );
  AO221X1 U3688 ( .IN1(n4422), .IN2(n3092), .IN3(n4371), .IN4(n4212), .IN5(
        n4444), .Q(n2715) );
  AO21X1 U3689 ( .IN1(n4424), .IN2(n3095), .IN3(n4445), .Q(n4444) );
  MUX21X1 U3690 ( .IN1(n4214), .IN2(n4446), .S(n4440), .Q(n4445) );
  AO221X1 U3691 ( .IN1(n4422), .IN2(n3094), .IN3(n4371), .IN4(n4216), .IN5(
        n4447), .Q(n2714) );
  AO21X1 U3692 ( .IN1(n4424), .IN2(n2843), .IN3(n4448), .Q(n4447) );
  MUX21X1 U3693 ( .IN1(n4218), .IN2(test_so12), .S(n4440), .Q(n4448) );
  NOR4X0 U3694 ( .IN1(n4174), .IN2(n4440), .IN3(n4371), .IN4(n4394), .QN(n4422) );
  INVX0 U3695 ( .IN(n4427), .QN(n4440) );
  AO221X1 U3696 ( .IN1(n4419), .IN2(n4012), .IN3(n4450), .IN4(n4221), .IN5(
        n4451), .Q(n4427) );
  NAND2X0 U3697 ( .IN1(n4452), .IN2(n4421), .QN(n4451) );
  INVX0 U3698 ( .IN(n4399), .QN(n4421) );
  NAND3X0 U3699 ( .IN1(n1553), .IN2(N3990), .IN3(n4340), .QN(n4418) );
  AO221X1 U3700 ( .IN1(n4453), .IN2(n3080), .IN3(n4394), .IN4(n4185), .IN5(
        n4454), .Q(n2713) );
  AO21X1 U3701 ( .IN1(n4455), .IN2(n3101), .IN3(n4456), .Q(n4454) );
  MUX21X1 U3702 ( .IN1(n4457), .IN2(n4188), .S(n4458), .Q(n4456) );
  AO221X1 U3703 ( .IN1(n4453), .IN2(n3082), .IN3(n4394), .IN4(n4191), .IN5(
        n4459), .Q(n2712) );
  AO21X1 U3704 ( .IN1(n4455), .IN2(n3100), .IN3(n4460), .Q(n4459) );
  MUX21X1 U3705 ( .IN1(n4461), .IN2(n4193), .S(n4458), .Q(n4460) );
  AO221X1 U3706 ( .IN1(n4453), .IN2(n3084), .IN3(n4394), .IN4(n4195), .IN5(
        n4462), .Q(n2711) );
  AO21X1 U3707 ( .IN1(n4455), .IN2(n3099), .IN3(n4463), .Q(n4462) );
  MUX21X1 U3708 ( .IN1(n4464), .IN2(n4197), .S(n4458), .Q(n4463) );
  AO221X1 U3709 ( .IN1(n4453), .IN2(n3086), .IN3(n4394), .IN4(n4199), .IN5(
        n4465), .Q(n2710) );
  AO21X1 U3710 ( .IN1(n4455), .IN2(n3098), .IN3(n4466), .Q(n4465) );
  MUX21X1 U3711 ( .IN1(n4201), .IN2(n4467), .S(n4468), .Q(n4466) );
  AO221X1 U3712 ( .IN1(n4453), .IN2(n3088), .IN3(n4394), .IN4(n4203), .IN5(
        n4469), .Q(n2709) );
  AO21X1 U3713 ( .IN1(n4455), .IN2(n3097), .IN3(n4470), .Q(n4469) );
  MUX21X1 U3714 ( .IN1(n4205), .IN2(n4471), .S(n4468), .Q(n4470) );
  AO221X1 U3715 ( .IN1(n4453), .IN2(n3090), .IN3(n4394), .IN4(n4208), .IN5(
        n4472), .Q(n2708) );
  AO21X1 U3716 ( .IN1(n4455), .IN2(n3096), .IN3(n4473), .Q(n4472) );
  MUX21X1 U3717 ( .IN1(n4210), .IN2(n4474), .S(n4468), .Q(n4473) );
  AO221X1 U3718 ( .IN1(n4453), .IN2(n3092), .IN3(n4394), .IN4(n4212), .IN5(
        n4475), .Q(n2707) );
  AO21X1 U3719 ( .IN1(n4455), .IN2(n3095), .IN3(n4476), .Q(n4475) );
  MUX21X1 U3720 ( .IN1(n4214), .IN2(n4477), .S(n4468), .Q(n4476) );
  AO221X1 U3721 ( .IN1(n4453), .IN2(n3094), .IN3(n4394), .IN4(n4216), .IN5(
        n4478), .Q(n2706) );
  AO21X1 U3722 ( .IN1(n4455), .IN2(n2843), .IN3(n4479), .Q(n4478) );
  MUX21X1 U3723 ( .IN1(n4218), .IN2(n4480), .S(n4468), .Q(n4479) );
  INVX0 U3724 ( .IN(n4458), .QN(n4468) );
  INVX0 U3725 ( .IN(n4481), .QN(n4455) );
  AND4X1 U3726 ( .IN1(n4254), .IN2(n4458), .IN3(n4482), .IN4(n4173), .Q(n4453)
         );
  AO221X1 U3727 ( .IN1(n4450), .IN2(n4012), .IN3(n4483), .IN4(n4221), .IN5(
        n4484), .Q(n4458) );
  NAND2X0 U3728 ( .IN1(n4481), .IN2(n4452), .QN(n4484) );
  INVX0 U3729 ( .IN(n4424), .QN(n4452) );
  NAND3X0 U3730 ( .IN1(n4485), .IN2(n1556), .IN3(n1553), .QN(n4482) );
  AO221X1 U3731 ( .IN1(n4486), .IN2(n3080), .IN3(n4185), .IN4(n4419), .IN5(
        n4487), .Q(n2705) );
  AO21X1 U3732 ( .IN1(n4488), .IN2(n3101), .IN3(n4489), .Q(n4487) );
  MUX21X1 U3733 ( .IN1(n2854), .IN2(n4188), .S(n4490), .Q(n4489) );
  AO221X1 U3734 ( .IN1(n4486), .IN2(n3082), .IN3(n4191), .IN4(n4419), .IN5(
        n4491), .Q(n2704) );
  AO21X1 U3735 ( .IN1(n4488), .IN2(n3100), .IN3(n4492), .Q(n4491) );
  MUX21X1 U3736 ( .IN1(n2855), .IN2(n4193), .S(n4490), .Q(n4492) );
  AO221X1 U3737 ( .IN1(n4486), .IN2(n3084), .IN3(n4195), .IN4(n4419), .IN5(
        n4493), .Q(n2703) );
  AO21X1 U3738 ( .IN1(n4488), .IN2(n3099), .IN3(n4494), .Q(n4493) );
  MUX21X1 U3739 ( .IN1(n2856), .IN2(n4197), .S(n4490), .Q(n4494) );
  AO221X1 U3740 ( .IN1(n4486), .IN2(n3086), .IN3(n4199), .IN4(n4419), .IN5(
        n4495), .Q(n2702) );
  AO21X1 U3741 ( .IN1(n4488), .IN2(n3098), .IN3(n4496), .Q(n4495) );
  MUX21X1 U3742 ( .IN1(n4201), .IN2(n2849), .S(n4497), .Q(n4496) );
  AO221X1 U3743 ( .IN1(n4486), .IN2(n3088), .IN3(n4203), .IN4(n4419), .IN5(
        n4498), .Q(n2701) );
  AO21X1 U3744 ( .IN1(n4488), .IN2(n3097), .IN3(n4499), .Q(n4498) );
  MUX21X1 U3745 ( .IN1(n4205), .IN2(n2850), .S(n4497), .Q(n4499) );
  AO221X1 U3746 ( .IN1(n4486), .IN2(n3090), .IN3(n4208), .IN4(n4419), .IN5(
        n4500), .Q(n2700) );
  AO21X1 U3747 ( .IN1(n4488), .IN2(n3096), .IN3(n4501), .Q(n4500) );
  MUX21X1 U3748 ( .IN1(n4210), .IN2(n2851), .S(n4497), .Q(n4501) );
  AO221X1 U3749 ( .IN1(n4486), .IN2(n3092), .IN3(n4212), .IN4(n4419), .IN5(
        n4502), .Q(n2699) );
  AO21X1 U3750 ( .IN1(n4488), .IN2(n3095), .IN3(n4503), .Q(n4502) );
  MUX21X1 U3751 ( .IN1(n4214), .IN2(n2852), .S(n4497), .Q(n4503) );
  AO221X1 U3752 ( .IN1(n4486), .IN2(n3094), .IN3(n4216), .IN4(n4419), .IN5(
        n4504), .Q(n2698) );
  AO21X1 U3753 ( .IN1(n4488), .IN2(n2843), .IN3(n4505), .Q(n4504) );
  MUX21X1 U3754 ( .IN1(n4218), .IN2(n2853), .S(n4497), .Q(n4505) );
  INVX0 U3755 ( .IN(n4490), .QN(n4497) );
  AND4X1 U3756 ( .IN1(n4254), .IN2(n4490), .IN3(n4173), .IN4(n4506), .Q(n4486)
         );
  AO221X1 U3757 ( .IN1(n4483), .IN2(n4012), .IN3(n4507), .IN4(n4221), .IN5(
        n4508), .Q(n4490) );
  NAND2X0 U3758 ( .IN1(n4509), .IN2(n4481), .QN(n4508) );
  NAND2X0 U3759 ( .IN1(n3392), .IN2(n4419), .QN(n4481) );
  NAND3X0 U3760 ( .IN1(n4485), .IN2(N1239), .IN3(n1553), .QN(n4173) );
  AO221X1 U3761 ( .IN1(n4510), .IN2(n3080), .IN3(n4450), .IN4(n4185), .IN5(
        n4511), .Q(n2697) );
  AO21X1 U3762 ( .IN1(n4512), .IN2(n3101), .IN3(n4513), .Q(n4511) );
  MUX21X1 U3763 ( .IN1(n2924), .IN2(n4188), .S(n4514), .Q(n4513) );
  AO221X1 U3764 ( .IN1(n4510), .IN2(n3082), .IN3(n4450), .IN4(n4191), .IN5(
        n4515), .Q(n2696) );
  AO21X1 U3765 ( .IN1(n4512), .IN2(n3100), .IN3(n4516), .Q(n4515) );
  MUX21X1 U3766 ( .IN1(n2925), .IN2(n4193), .S(n4514), .Q(n4516) );
  AO221X1 U3767 ( .IN1(n4510), .IN2(n3084), .IN3(n4450), .IN4(n4195), .IN5(
        n4517), .Q(n2695) );
  AO21X1 U3768 ( .IN1(n4512), .IN2(n3099), .IN3(n4518), .Q(n4517) );
  MUX21X1 U3769 ( .IN1(n2926), .IN2(n4197), .S(n4514), .Q(n4518) );
  AO221X1 U3770 ( .IN1(n4510), .IN2(n3086), .IN3(n4450), .IN4(n4199), .IN5(
        n4519), .Q(n2694) );
  AO21X1 U3771 ( .IN1(n4512), .IN2(n3098), .IN3(n4520), .Q(n4519) );
  MUX21X1 U3772 ( .IN1(n2927), .IN2(n4201), .S(n4514), .Q(n4520) );
  AO221X1 U3773 ( .IN1(n4510), .IN2(n3088), .IN3(n4450), .IN4(n4203), .IN5(
        n4521), .Q(n2693) );
  AO21X1 U3774 ( .IN1(n4512), .IN2(n3097), .IN3(n4522), .Q(n4521) );
  MUX21X1 U3775 ( .IN1(n4205), .IN2(test_so13), .S(n4523), .Q(n4522) );
  AO221X1 U3776 ( .IN1(n4510), .IN2(n3090), .IN3(n4450), .IN4(n4208), .IN5(
        n4524), .Q(n2692) );
  AO21X1 U3777 ( .IN1(n4512), .IN2(n3096), .IN3(n4525), .Q(n4524) );
  MUX21X1 U3778 ( .IN1(n4210), .IN2(n2908), .S(n4523), .Q(n4525) );
  AO221X1 U3779 ( .IN1(n4510), .IN2(n3092), .IN3(n4450), .IN4(n4212), .IN5(
        n4526), .Q(n2691) );
  AO21X1 U3780 ( .IN1(n4512), .IN2(n3095), .IN3(n4527), .Q(n4526) );
  MUX21X1 U3781 ( .IN1(n4214), .IN2(n2909), .S(n4523), .Q(n4527) );
  AO221X1 U3782 ( .IN1(n4510), .IN2(n3094), .IN3(n4450), .IN4(n4216), .IN5(
        n4528), .Q(n2690) );
  AO21X1 U3783 ( .IN1(n4512), .IN2(n2843), .IN3(n4529), .Q(n4528) );
  MUX21X1 U3784 ( .IN1(n4218), .IN2(n2910), .S(n4523), .Q(n4529) );
  NOR4X0 U3785 ( .IN1(n4174), .IN2(n4523), .IN3(n4450), .IN4(n4483), .QN(n4510) );
  INVX0 U3786 ( .IN(n4514), .QN(n4523) );
  AO221X1 U3787 ( .IN1(n4507), .IN2(n4012), .IN3(n4530), .IN4(n4221), .IN5(
        n4531), .Q(n4514) );
  NAND2X0 U3788 ( .IN1(n4532), .IN2(n4509), .QN(n4531) );
  INVX0 U3789 ( .IN(n4488), .QN(n4509) );
  NAND3X0 U3790 ( .IN1(n1554), .IN2(N3989), .IN3(n4308), .QN(n4506) );
  AO221X1 U3791 ( .IN1(n4533), .IN2(n3080), .IN3(n4483), .IN4(n4185), .IN5(
        n4534), .Q(n2689) );
  AO21X1 U3792 ( .IN1(n4535), .IN2(n3101), .IN3(n4536), .Q(n4534) );
  MUX21X1 U3793 ( .IN1(n4537), .IN2(n4188), .S(n4538), .Q(n4536) );
  AO221X1 U3794 ( .IN1(n4533), .IN2(n3082), .IN3(n4483), .IN4(n4191), .IN5(
        n4539), .Q(n2688) );
  AO21X1 U3795 ( .IN1(n4535), .IN2(n3100), .IN3(n4540), .Q(n4539) );
  MUX21X1 U3796 ( .IN1(n4541), .IN2(n4193), .S(n4538), .Q(n4540) );
  AO221X1 U3797 ( .IN1(n4533), .IN2(n3084), .IN3(n4483), .IN4(n4195), .IN5(
        n4542), .Q(n2687) );
  AO21X1 U3798 ( .IN1(n4535), .IN2(n3099), .IN3(n4543), .Q(n4542) );
  MUX21X1 U3799 ( .IN1(n4544), .IN2(n4197), .S(n4538), .Q(n4543) );
  AO221X1 U3800 ( .IN1(n4533), .IN2(n3086), .IN3(n4483), .IN4(n4199), .IN5(
        n4545), .Q(n2686) );
  AO21X1 U3801 ( .IN1(n4535), .IN2(n3098), .IN3(n4546), .Q(n4545) );
  MUX21X1 U3802 ( .IN1(n4201), .IN2(n4547), .S(n4548), .Q(n4546) );
  AO221X1 U3803 ( .IN1(n4533), .IN2(n3088), .IN3(n4483), .IN4(n4203), .IN5(
        n4549), .Q(n2685) );
  AO21X1 U3804 ( .IN1(n4535), .IN2(n3097), .IN3(n4550), .Q(n4549) );
  MUX21X1 U3805 ( .IN1(n4205), .IN2(n4551), .S(n4548), .Q(n4550) );
  AO221X1 U3806 ( .IN1(n4533), .IN2(n3090), .IN3(n4483), .IN4(n4208), .IN5(
        n4552), .Q(n2684) );
  AO21X1 U3807 ( .IN1(n4535), .IN2(n3096), .IN3(n4553), .Q(n4552) );
  MUX21X1 U3808 ( .IN1(n4210), .IN2(n4554), .S(n4548), .Q(n4553) );
  AO221X1 U3809 ( .IN1(n4533), .IN2(n3092), .IN3(n4483), .IN4(n4212), .IN5(
        n4555), .Q(n2683) );
  AO21X1 U3810 ( .IN1(n4535), .IN2(n3095), .IN3(n4556), .Q(n4555) );
  MUX21X1 U3811 ( .IN1(n4214), .IN2(n4557), .S(n4548), .Q(n4556) );
  AO221X1 U3812 ( .IN1(n4533), .IN2(n3094), .IN3(n4483), .IN4(n4216), .IN5(
        n4558), .Q(n2682) );
  AO21X1 U3813 ( .IN1(n4535), .IN2(n2843), .IN3(n4559), .Q(n4558) );
  MUX21X1 U3814 ( .IN1(n4218), .IN2(n4560), .S(n4548), .Q(n4559) );
  INVX0 U3815 ( .IN(n4538), .QN(n4548) );
  AND4X1 U3816 ( .IN1(n4254), .IN2(n4538), .IN3(n4561), .IN4(n4562), .Q(n4533)
         );
  AO221X1 U3817 ( .IN1(n4530), .IN2(n4012), .IN3(n4563), .IN4(n4221), .IN5(
        n4564), .Q(n4538) );
  NAND2X0 U3818 ( .IN1(n4565), .IN2(n4532), .QN(n4564) );
  INVX0 U3819 ( .IN(n4512), .QN(n4532) );
  NAND3X0 U3820 ( .IN1(n1554), .IN2(N3989), .IN3(n4340), .QN(n4561) );
  AO221X1 U3821 ( .IN1(n4566), .IN2(n3080), .IN3(n4507), .IN4(n4185), .IN5(
        n4567), .Q(n2681) );
  AO21X1 U3822 ( .IN1(n4568), .IN2(n3101), .IN3(n4569), .Q(n4567) );
  MUX21X1 U3823 ( .IN1(n4570), .IN2(n4188), .S(n4571), .Q(n4569) );
  AO221X1 U3824 ( .IN1(n4566), .IN2(n3082), .IN3(n4507), .IN4(n4191), .IN5(
        n4572), .Q(n2680) );
  AO21X1 U3825 ( .IN1(n4568), .IN2(n3100), .IN3(n4573), .Q(n4572) );
  MUX21X1 U3826 ( .IN1(n4574), .IN2(n4193), .S(n4571), .Q(n4573) );
  AO221X1 U3827 ( .IN1(n4566), .IN2(n3084), .IN3(n4507), .IN4(n4195), .IN5(
        n4575), .Q(n2679) );
  AO21X1 U3828 ( .IN1(n4568), .IN2(n3099), .IN3(n4576), .Q(n4575) );
  MUX21X1 U3829 ( .IN1(n4577), .IN2(n4197), .S(n4571), .Q(n4576) );
  AO221X1 U3830 ( .IN1(n4566), .IN2(n3086), .IN3(n4507), .IN4(n4199), .IN5(
        n4578), .Q(n2678) );
  AO21X1 U3831 ( .IN1(n4568), .IN2(n3098), .IN3(n4579), .Q(n4578) );
  MUX21X1 U3832 ( .IN1(n4201), .IN2(n4580), .S(n4581), .Q(n4579) );
  AO221X1 U3833 ( .IN1(n4566), .IN2(n3088), .IN3(n4507), .IN4(n4203), .IN5(
        n4582), .Q(n2677) );
  AO21X1 U3834 ( .IN1(n4568), .IN2(n3097), .IN3(n4583), .Q(n4582) );
  MUX21X1 U3835 ( .IN1(n4205), .IN2(n4584), .S(n4581), .Q(n4583) );
  AO221X1 U3836 ( .IN1(n4566), .IN2(n3090), .IN3(n4507), .IN4(n4208), .IN5(
        n4585), .Q(n2676) );
  AO21X1 U3837 ( .IN1(n4568), .IN2(n3096), .IN3(n4586), .Q(n4585) );
  MUX21X1 U3838 ( .IN1(n4210), .IN2(n4587), .S(n4581), .Q(n4586) );
  AO221X1 U3839 ( .IN1(n4566), .IN2(n3092), .IN3(n4507), .IN4(n4212), .IN5(
        n4588), .Q(n2675) );
  AO21X1 U3840 ( .IN1(n4568), .IN2(n3095), .IN3(n4589), .Q(n4588) );
  MUX21X1 U3841 ( .IN1(n4214), .IN2(n4590), .S(n4581), .Q(n4589) );
  AO221X1 U3842 ( .IN1(n4566), .IN2(n3094), .IN3(n4507), .IN4(n4216), .IN5(
        n4591), .Q(n2674) );
  AO21X1 U3843 ( .IN1(n4568), .IN2(n2843), .IN3(n4592), .Q(n4591) );
  MUX21X1 U3844 ( .IN1(n4218), .IN2(n4593), .S(n4581), .Q(n4592) );
  INVX0 U3845 ( .IN(n4571), .QN(n4581) );
  AND4X1 U3846 ( .IN1(n4254), .IN2(n4571), .IN3(n4562), .IN4(n4594), .Q(n4566)
         );
  AO221X1 U3847 ( .IN1(n4186), .IN2(n4221), .IN3(n4563), .IN4(n4012), .IN5(
        n4595), .Q(n4571) );
  NAND2X0 U3848 ( .IN1(n4596), .IN2(n4565), .QN(n4595) );
  INVX0 U3849 ( .IN(n4535), .QN(n4565) );
  NAND3X0 U3850 ( .IN1(n1556), .IN2(N3989), .IN3(n4162), .QN(n4562) );
  AO221X1 U3851 ( .IN1(n4597), .IN2(n3080), .IN3(n4530), .IN4(n4185), .IN5(
        n4598), .Q(n2673) );
  AO21X1 U3852 ( .IN1(n4599), .IN2(n3101), .IN3(n4600), .Q(n4598) );
  MUX21X1 U3853 ( .IN1(n2876), .IN2(n4188), .S(n4601), .Q(n4600) );
  AO221X1 U3854 ( .IN1(n4597), .IN2(n3082), .IN3(n4530), .IN4(n4191), .IN5(
        n4602), .Q(n2672) );
  AO21X1 U3855 ( .IN1(n4599), .IN2(n3100), .IN3(n4603), .Q(n4602) );
  MUX21X1 U3856 ( .IN1(test_so14), .IN2(n4193), .S(n4601), .Q(n4603) );
  AO221X1 U3857 ( .IN1(n4597), .IN2(n3084), .IN3(n4530), .IN4(n4195), .IN5(
        n4604), .Q(n2671) );
  AO21X1 U3858 ( .IN1(n4599), .IN2(n3099), .IN3(n4605), .Q(n4604) );
  MUX21X1 U3859 ( .IN1(n2878), .IN2(n4197), .S(n4601), .Q(n4605) );
  AO221X1 U3860 ( .IN1(n4597), .IN2(n3086), .IN3(n4530), .IN4(n4199), .IN5(
        n4606), .Q(n2670) );
  AO21X1 U3861 ( .IN1(n4599), .IN2(n3098), .IN3(n4607), .Q(n4606) );
  MUX21X1 U3862 ( .IN1(n4201), .IN2(n2871), .S(n4608), .Q(n4607) );
  AO221X1 U3863 ( .IN1(n4597), .IN2(n3088), .IN3(n4530), .IN4(n4203), .IN5(
        n4609), .Q(n2669) );
  AO21X1 U3864 ( .IN1(n4599), .IN2(n3097), .IN3(n4610), .Q(n4609) );
  MUX21X1 U3865 ( .IN1(n4205), .IN2(n2872), .S(n4608), .Q(n4610) );
  AO221X1 U3866 ( .IN1(n4597), .IN2(n3090), .IN3(n4530), .IN4(n4208), .IN5(
        n4611), .Q(n2668) );
  AO21X1 U3867 ( .IN1(n4599), .IN2(n3096), .IN3(n4612), .Q(n4611) );
  MUX21X1 U3868 ( .IN1(n4210), .IN2(n2873), .S(n4608), .Q(n4612) );
  AO221X1 U3869 ( .IN1(n4597), .IN2(n3092), .IN3(n4530), .IN4(n4212), .IN5(
        n4613), .Q(n2667) );
  AO21X1 U3870 ( .IN1(n4599), .IN2(n3095), .IN3(n4614), .Q(n4613) );
  MUX21X1 U3871 ( .IN1(n4214), .IN2(n2874), .S(n4608), .Q(n4614) );
  AO221X1 U3872 ( .IN1(n4597), .IN2(n3094), .IN3(n4530), .IN4(n4216), .IN5(
        n4615), .Q(n2666) );
  AO21X1 U3873 ( .IN1(n4599), .IN2(n2843), .IN3(n4616), .Q(n4615) );
  MUX21X1 U3874 ( .IN1(n4218), .IN2(n2875), .S(n4608), .Q(n4616) );
  INVX0 U3875 ( .IN(n4601), .QN(n4608) );
  AND4X1 U3876 ( .IN1(n4254), .IN2(n4601), .IN3(n4594), .IN4(n4617), .Q(n4597)
         );
  AO221X1 U3877 ( .IN1(n4186), .IN2(n4012), .IN3(n4219), .IN4(n4221), .IN5(
        n4618), .Q(n4601) );
  NAND2X0 U3878 ( .IN1(n4619), .IN2(n4596), .QN(n4618) );
  INVX0 U3879 ( .IN(n4568), .QN(n4596) );
  NAND2X0 U3880 ( .IN1(n4159), .IN2(N3989), .QN(n4594) );
  AND2X1 U3881 ( .IN1(n4162), .IN2(N1239), .Q(n4159) );
  NOR2X0 U3882 ( .IN1(N3990), .IN2(n1555), .QN(n4162) );
  AO221X1 U3883 ( .IN1(n4563), .IN2(n4185), .IN3(n4621), .IN4(n3080), .IN5(
        n4622), .Q(n2665) );
  AO21X1 U3884 ( .IN1(n4623), .IN2(n3101), .IN3(n4624), .Q(n4622) );
  MUX21X1 U3885 ( .IN1(n2928), .IN2(n4188), .S(n4625), .Q(n4624) );
  AO221X1 U3886 ( .IN1(n4563), .IN2(n4191), .IN3(n4621), .IN4(n3082), .IN5(
        n4626), .Q(n2664) );
  AO21X1 U3887 ( .IN1(n4623), .IN2(n3100), .IN3(n4627), .Q(n4626) );
  MUX21X1 U3888 ( .IN1(n2929), .IN2(n4193), .S(n4625), .Q(n4627) );
  AO221X1 U3889 ( .IN1(n4563), .IN2(n4195), .IN3(n4621), .IN4(n3084), .IN5(
        n4629), .Q(n2663) );
  AO21X1 U3890 ( .IN1(n4623), .IN2(n3099), .IN3(n4630), .Q(n4629) );
  MUX21X1 U3891 ( .IN1(n2930), .IN2(n4197), .S(n4625), .Q(n4630) );
  AO221X1 U3892 ( .IN1(n4563), .IN2(n4199), .IN3(n4621), .IN4(n3086), .IN5(
        n4632), .Q(n2662) );
  AO21X1 U3893 ( .IN1(n4623), .IN2(n3098), .IN3(n4633), .Q(n4632) );
  MUX21X1 U3894 ( .IN1(n4201), .IN2(n2911), .S(n4634), .Q(n4633) );
  AO221X1 U3895 ( .IN1(n4563), .IN2(n4203), .IN3(n4621), .IN4(n3088), .IN5(
        n4636), .Q(n2661) );
  AO21X1 U3896 ( .IN1(n4623), .IN2(n3097), .IN3(n4637), .Q(n4636) );
  MUX21X1 U3897 ( .IN1(n4205), .IN2(n2912), .S(n4634), .Q(n4637) );
  AO221X1 U3898 ( .IN1(n4563), .IN2(n4208), .IN3(n4621), .IN4(n3090), .IN5(
        n4639), .Q(n2660) );
  AO21X1 U3899 ( .IN1(n4623), .IN2(n3096), .IN3(n4640), .Q(n4639) );
  MUX21X1 U3900 ( .IN1(n4210), .IN2(n2913), .S(n4634), .Q(n4640) );
  AO221X1 U3901 ( .IN1(n4563), .IN2(n4212), .IN3(n4621), .IN4(n3092), .IN5(
        n4642), .Q(n2659) );
  AO21X1 U3902 ( .IN1(n4623), .IN2(n3095), .IN3(n4643), .Q(n4642) );
  MUX21X1 U3903 ( .IN1(n4214), .IN2(n2914), .S(n4634), .Q(n4643) );
  AO221X1 U3904 ( .IN1(n4621), .IN2(n3094), .IN3(n4563), .IN4(n4216), .IN5(
        n4645), .Q(n2658) );
  AO21X1 U3905 ( .IN1(n4623), .IN2(n2843), .IN3(n4646), .Q(n4645) );
  MUX21X1 U3906 ( .IN1(n4218), .IN2(n2915), .S(n4634), .Q(n4646) );
  INVX0 U3907 ( .IN(n4625), .QN(n4634) );
  AND4X1 U3908 ( .IN1(n4254), .IN2(n4625), .IN3(n4620), .IN4(n4617), .Q(n4621)
         );
  AO221X1 U3909 ( .IN1(n4222), .IN2(n4221), .IN3(n4219), .IN4(n4012), .IN5(
        n4648), .Q(n4625) );
  NAND2X0 U3910 ( .IN1(n4619), .IN2(n4224), .QN(n4648) );
  INVX0 U3911 ( .IN(n4623), .QN(n4224) );
  NAND3X0 U3912 ( .IN1(N3989), .IN2(N3990), .IN3(n4340), .QN(n4620) );
  NOR2X0 U3913 ( .IN1(N3991), .IN2(n1556), .QN(n4340) );
  INVX0 U3914 ( .IN(n4599), .QN(n4619) );
  NAND3X0 U3915 ( .IN1(N3989), .IN2(N3990), .IN3(n4308), .QN(n4617) );
  NOR2X0 U3916 ( .IN1(N3991), .IN2(N1239), .QN(n4308) );
  NAND3X0 U3917 ( .IN1(n1556), .IN2(N3989), .IN3(n4485), .QN(n4256) );
  NOR2X0 U3918 ( .IN1(n4012), .IN2(n4081), .QN(n4181) );
  NOR2X0 U3919 ( .IN1(InstQueueRd_Addr[4]), .IN2(n4095), .QN(n4081) );
  NAND3X0 U3920 ( .IN1(n1492), .IN2(n4097), .IN3(n4649), .QN(n4095) );
  NAND3X0 U3921 ( .IN1(N3989), .IN2(N1239), .IN3(n4485), .QN(n4255) );
  INVX0 U3922 ( .IN(n4176), .QN(n4485) );
  NAND2X0 U3923 ( .IN1(N3990), .IN2(N3991), .QN(n4176) );
  INVX0 U3924 ( .IN(n4650), .QN(n2657) );
  MUX21X1 U3925 ( .IN1(n3873), .IN2(n4108), .S(n4131), .Q(n4650) );
  ISOLANDX1 U3926 ( .D(n4110), .ISO(n4091), .Q(n4131) );
  NAND4X0 U3927 ( .IN1(n4651), .IN2(n4652), .IN3(n4653), .IN4(n4654), .QN(
        n4110) );
  NOR3X0 U3928 ( .IN1(n4655), .IN2(n4656), .IN3(n4657), .QN(n4654) );
  INVX0 U3929 ( .IN(n4658), .QN(n4653) );
  NAND2X0 U3930 ( .IN1(n4659), .IN2(n2948), .QN(n4652) );
  AOI222X1 U3931 ( .IN1(n4660), .IN2(n4661), .IN3(n4662), .IN4(n4123), .IN5(
        n4657), .IN6(n4663), .QN(n4108) );
  NAND4X0 U3932 ( .IN1(n4664), .IN2(n4665), .IN3(n4666), .IN4(n4667), .QN(
        n2656) );
  AOI221X1 U3933 ( .IN1(N1769), .IN2(n3233), .IN3(N1956), .IN4(n3250), .IN5(
        n4668), .QN(n4667) );
  AO22X1 U3934 ( .IN1(n3230), .IN2(EBX_0_), .IN3(n1552), .IN4(n4669), .Q(n4668) );
  OA22X1 U3935 ( .IN1(n3103), .IN2(n2845), .IN3(n1589), .IN4(n3105), .Q(n4666)
         );
  NAND2X0 U3936 ( .IN1(N997), .IN2(n3241), .QN(n4665) );
  NAND2X0 U3937 ( .IN1(N1031), .IN2(n3220), .QN(n4664) );
  NAND4X0 U3938 ( .IN1(n4670), .IN2(n4671), .IN3(n4672), .IN4(n4673), .QN(
        n2655) );
  AOI221X1 U3939 ( .IN1(N1770), .IN2(n3233), .IN3(N1957), .IN4(n3250), .IN5(
        n4674), .QN(n4673) );
  AO22X1 U3940 ( .IN1(n3230), .IN2(EBX_1_), .IN3(N2700), .IN4(n4669), .Q(n4674) );
  OA22X1 U3941 ( .IN1(n3103), .IN2(n2888), .IN3(n1588), .IN4(n3105), .Q(n4672)
         );
  NAND2X0 U3942 ( .IN1(N998), .IN2(n3241), .QN(n4671) );
  NAND2X0 U3943 ( .IN1(N1032), .IN2(n3220), .QN(n4670) );
  NAND4X0 U3944 ( .IN1(n4675), .IN2(n4676), .IN3(n4677), .IN4(n4678), .QN(
        n2654) );
  AOI221X1 U3945 ( .IN1(N1771), .IN2(n3234), .IN3(N1958), .IN4(n3250), .IN5(
        n4679), .QN(n4678) );
  AO22X1 U3946 ( .IN1(n3230), .IN2(EBX_2_), .IN3(N2701), .IN4(n4669), .Q(n4679) );
  OA22X1 U3947 ( .IN1(n3102), .IN2(n4680), .IN3(n1587), .IN4(n3104), .Q(n4677)
         );
  NAND2X0 U3948 ( .IN1(N999), .IN2(n3242), .QN(n4676) );
  NAND2X0 U3949 ( .IN1(N1033), .IN2(n3221), .QN(n4675) );
  NAND4X0 U3950 ( .IN1(n4681), .IN2(n4682), .IN3(n4683), .IN4(n4684), .QN(
        n2653) );
  AOI221X1 U3951 ( .IN1(N1772), .IN2(n3233), .IN3(N1959), .IN4(n3250), .IN5(
        n4685), .QN(n4684) );
  AO22X1 U3952 ( .IN1(n3230), .IN2(EBX_3_), .IN3(N2702), .IN4(n4669), .Q(n4685) );
  OA22X1 U3953 ( .IN1(n3103), .IN2(n4686), .IN3(n1586), .IN4(n3105), .Q(n4683)
         );
  NAND2X0 U3954 ( .IN1(N1000), .IN2(n3241), .QN(n4682) );
  NAND2X0 U3955 ( .IN1(N1034), .IN2(n3220), .QN(n4681) );
  NAND4X0 U3956 ( .IN1(n4687), .IN2(n4688), .IN3(n4689), .IN4(n4690), .QN(
        n2652) );
  AOI221X1 U3957 ( .IN1(N1773), .IN2(n3234), .IN3(N1960), .IN4(n3250), .IN5(
        n4691), .QN(n4690) );
  AO221X1 U3958 ( .IN1(N2703), .IN2(n4669), .IN3(n3227), .IN4(EBX_4_), .IN5(
        n3204), .Q(n4691) );
  OA22X1 U3959 ( .IN1(n3102), .IN2(n4692), .IN3(n1585), .IN4(n3104), .Q(n4689)
         );
  NAND2X0 U3960 ( .IN1(N1001), .IN2(n3242), .QN(n4688) );
  NAND2X0 U3961 ( .IN1(N1035), .IN2(n3221), .QN(n4687) );
  NAND4X0 U3962 ( .IN1(n4693), .IN2(n4694), .IN3(n4695), .IN4(n4696), .QN(
        n2651) );
  AOI221X1 U3963 ( .IN1(N1774), .IN2(n3234), .IN3(N1961), .IN4(n3251), .IN5(
        n4697), .QN(n4696) );
  AO221X1 U3964 ( .IN1(N2704), .IN2(n4669), .IN3(n3227), .IN4(EBX_5_), .IN5(
        n3195), .Q(n4697) );
  ISOLANDX1 U3965 ( .D(n4698), .ISO(n4699), .Q(n4669) );
  OA22X1 U3966 ( .IN1(n3102), .IN2(n4700), .IN3(n1584), .IN4(n3105), .Q(n4695)
         );
  NAND2X0 U3967 ( .IN1(N1002), .IN2(n3241), .QN(n4694) );
  NAND2X0 U3968 ( .IN1(N1036), .IN2(n3221), .QN(n4693) );
  NAND4X0 U3969 ( .IN1(n4701), .IN2(n3185), .IN3(n4702), .IN4(n4703), .QN(
        n2650) );
  OA221X1 U3970 ( .IN1(n1583), .IN2(n3105), .IN3(n3102), .IN4(n4704), .IN5(
        n4705), .Q(n4703) );
  AOI22X1 U3971 ( .IN1(N1003), .IN2(n3245), .IN3(N1037), .IN4(n3223), .QN(
        n4705) );
  AOI22X1 U3972 ( .IN1(N1775), .IN2(n3236), .IN3(N1962), .IN4(n3256), .QN(
        n4702) );
  NAND2X0 U3973 ( .IN1(n3229), .IN2(EBX_6_), .QN(n4701) );
  NAND4X0 U3974 ( .IN1(n4706), .IN2(n3185), .IN3(n4707), .IN4(n4708), .QN(
        n2649) );
  OA221X1 U3975 ( .IN1(n1582), .IN2(n3105), .IN3(n3102), .IN4(n4709), .IN5(
        n4710), .Q(n4708) );
  AOI22X1 U3976 ( .IN1(N1004), .IN2(n3245), .IN3(N1038), .IN4(n3223), .QN(
        n4710) );
  AOI22X1 U3977 ( .IN1(N1776), .IN2(n3236), .IN3(N1963), .IN4(n3256), .QN(
        n4707) );
  NAND2X0 U3978 ( .IN1(n3228), .IN2(EBX_7_), .QN(n4706) );
  NAND4X0 U3979 ( .IN1(n4711), .IN2(n3186), .IN3(n4712), .IN4(n4713), .QN(
        n2648) );
  OA221X1 U3980 ( .IN1(n1581), .IN2(n3104), .IN3(n3102), .IN4(n4714), .IN5(
        n4715), .Q(n4713) );
  AOI22X1 U3981 ( .IN1(N1005), .IN2(n3245), .IN3(N1039), .IN4(n3224), .QN(
        n4715) );
  AOI22X1 U3982 ( .IN1(N1777), .IN2(n3237), .IN3(N1964), .IN4(n3255), .QN(
        n4712) );
  NAND2X0 U3983 ( .IN1(n3229), .IN2(EBX_8_), .QN(n4711) );
  NAND4X0 U3984 ( .IN1(n4716), .IN2(n3186), .IN3(n4717), .IN4(n4718), .QN(
        n2647) );
  OA221X1 U3985 ( .IN1(n1580), .IN2(n3105), .IN3(n3102), .IN4(n4719), .IN5(
        n4720), .Q(n4718) );
  AOI22X1 U3986 ( .IN1(N1006), .IN2(n3244), .IN3(N1040), .IN4(n3223), .QN(
        n4720) );
  AOI22X1 U3987 ( .IN1(N1778), .IN2(n3236), .IN3(N1965), .IN4(n3255), .QN(
        n4717) );
  NAND2X0 U3988 ( .IN1(n3229), .IN2(EBX_9_), .QN(n4716) );
  NAND4X0 U3989 ( .IN1(n4721), .IN2(n3186), .IN3(n4722), .IN4(n4723), .QN(
        n2646) );
  OA221X1 U3990 ( .IN1(n1579), .IN2(n3105), .IN3(n3103), .IN4(n4724), .IN5(
        n4725), .Q(n4723) );
  AOI22X1 U3991 ( .IN1(N1007), .IN2(n3245), .IN3(N1041), .IN4(n3224), .QN(
        n4725) );
  AOI22X1 U3992 ( .IN1(N1779), .IN2(n3237), .IN3(N1966), .IN4(n3255), .QN(
        n4722) );
  NAND2X0 U3993 ( .IN1(n3229), .IN2(EBX_10_), .QN(n4721) );
  NAND4X0 U3994 ( .IN1(n4726), .IN2(n3186), .IN3(n4727), .IN4(n4728), .QN(
        n2645) );
  OA221X1 U3995 ( .IN1(n1578), .IN2(n3105), .IN3(n3102), .IN4(n4729), .IN5(
        n4730), .Q(n4728) );
  AOI22X1 U3996 ( .IN1(N1008), .IN2(n3244), .IN3(N1042), .IN4(n3223), .QN(
        n4730) );
  AOI22X1 U3997 ( .IN1(N1780), .IN2(n3236), .IN3(N1967), .IN4(n3255), .QN(
        n4727) );
  NAND2X0 U3998 ( .IN1(n3229), .IN2(EBX_11_), .QN(n4726) );
  NAND4X0 U3999 ( .IN1(n4731), .IN2(n3186), .IN3(n4732), .IN4(n4733), .QN(
        n2644) );
  OA221X1 U4000 ( .IN1(n1577), .IN2(n3105), .IN3(n3102), .IN4(n4734), .IN5(
        n4735), .Q(n4733) );
  AOI22X1 U4001 ( .IN1(N1009), .IN2(n3243), .IN3(N1043), .IN4(n3222), .QN(
        n4735) );
  AOI22X1 U4002 ( .IN1(N1781), .IN2(n3235), .IN3(N1968), .IN4(n3255), .QN(
        n4732) );
  NAND2X0 U4003 ( .IN1(n3229), .IN2(EBX_12_), .QN(n4731) );
  NAND4X0 U4004 ( .IN1(n4736), .IN2(n3187), .IN3(n4737), .IN4(n4738), .QN(
        n2643) );
  OA221X1 U4005 ( .IN1(n1576), .IN2(n3105), .IN3(n3103), .IN4(n4739), .IN5(
        n4740), .Q(n4738) );
  AOI22X1 U4006 ( .IN1(N1010), .IN2(n3242), .IN3(N1044), .IN4(n3221), .QN(
        n4740) );
  AOI22X1 U4007 ( .IN1(N1782), .IN2(n3234), .IN3(N1969), .IN4(n3254), .QN(
        n4737) );
  NAND2X0 U4008 ( .IN1(n3228), .IN2(EBX_13_), .QN(n4736) );
  NAND4X0 U4009 ( .IN1(n4741), .IN2(n3187), .IN3(n4742), .IN4(n4743), .QN(
        n2642) );
  OA221X1 U4010 ( .IN1(n1575), .IN2(n3105), .IN3(n3103), .IN4(n4744), .IN5(
        n4745), .Q(n4743) );
  AOI22X1 U4011 ( .IN1(N1011), .IN2(n3244), .IN3(N1045), .IN4(n3223), .QN(
        n4745) );
  AOI22X1 U4012 ( .IN1(N1783), .IN2(n3236), .IN3(N1970), .IN4(n3254), .QN(
        n4742) );
  NAND2X0 U4013 ( .IN1(n3228), .IN2(EBX_14_), .QN(n4741) );
  NAND4X0 U4014 ( .IN1(n4746), .IN2(n3187), .IN3(n4747), .IN4(n4748), .QN(
        n2641) );
  OA221X1 U4015 ( .IN1(n1574), .IN2(n3105), .IN3(n3102), .IN4(n4749), .IN5(
        n4750), .Q(n4748) );
  AOI22X1 U4016 ( .IN1(N1012), .IN2(n3243), .IN3(N1046), .IN4(n3222), .QN(
        n4750) );
  AOI22X1 U4017 ( .IN1(N1784), .IN2(n3235), .IN3(N1971), .IN4(n3254), .QN(
        n4747) );
  NAND2X0 U4018 ( .IN1(n3228), .IN2(EBX_15_), .QN(n4746) );
  NAND4X0 U4019 ( .IN1(n4751), .IN2(n3187), .IN3(n4752), .IN4(n4753), .QN(
        n2640) );
  OA221X1 U4020 ( .IN1(n1573), .IN2(n3105), .IN3(n3102), .IN4(n4754), .IN5(
        n4755), .Q(n4753) );
  AOI22X1 U4021 ( .IN1(N1013), .IN2(n3242), .IN3(N1047), .IN4(n3221), .QN(
        n4755) );
  AOI22X1 U4022 ( .IN1(N1785), .IN2(n3234), .IN3(N1972), .IN4(n3254), .QN(
        n4752) );
  NAND2X0 U4023 ( .IN1(n3228), .IN2(EBX_16_), .QN(n4751) );
  NAND4X0 U4024 ( .IN1(n4756), .IN2(n3188), .IN3(n4757), .IN4(n4758), .QN(
        n2639) );
  OA221X1 U4025 ( .IN1(n1572), .IN2(n3105), .IN3(n3102), .IN4(n4759), .IN5(
        n4760), .Q(n4758) );
  AOI22X1 U4026 ( .IN1(N1014), .IN2(n3243), .IN3(N1048), .IN4(n3222), .QN(
        n4760) );
  AOI22X1 U4027 ( .IN1(N1786), .IN2(n3235), .IN3(N1973), .IN4(n3253), .QN(
        n4757) );
  NAND2X0 U4028 ( .IN1(n3228), .IN2(EBX_17_), .QN(n4756) );
  NAND4X0 U4029 ( .IN1(n4761), .IN2(n3187), .IN3(n4762), .IN4(n4763), .QN(
        n2638) );
  OA221X1 U4030 ( .IN1(n1571), .IN2(n3104), .IN3(n3103), .IN4(n4764), .IN5(
        n4765), .Q(n4763) );
  AOI22X1 U4031 ( .IN1(N1015), .IN2(n3244), .IN3(N1049), .IN4(n3222), .QN(
        n4765) );
  AOI22X1 U4032 ( .IN1(N1787), .IN2(n3235), .IN3(N1974), .IN4(n3253), .QN(
        n4762) );
  NAND2X0 U4033 ( .IN1(n3227), .IN2(EBX_18_), .QN(n4761) );
  NAND4X0 U4034 ( .IN1(n4766), .IN2(n3188), .IN3(n4767), .IN4(n4768), .QN(
        n2637) );
  OA221X1 U4035 ( .IN1(n1570), .IN2(n3104), .IN3(n3102), .IN4(n4769), .IN5(
        n4770), .Q(n4768) );
  AOI22X1 U4036 ( .IN1(N1016), .IN2(n3243), .IN3(N1050), .IN4(n3222), .QN(
        n4770) );
  AOI22X1 U4037 ( .IN1(N1788), .IN2(n3235), .IN3(N1975), .IN4(n3254), .QN(
        n4767) );
  NAND2X0 U4038 ( .IN1(n3227), .IN2(test_so6), .QN(n4766) );
  OR2X1 U4039 ( .IN1(n4771), .IN2(n4772), .Q(n2636) );
  AO222X1 U4040 ( .IN1(rEIP_20_), .IN2(n2952), .IN3(N1051), .IN4(n3220), .IN5(
        n2956), .IN6(PhyAddrPointer_20_), .Q(n4772) );
  AO221X1 U4041 ( .IN1(n3227), .IN2(EBX_20_), .IN3(N1789), .IN4(n3233), .IN5(
        n4773), .Q(n4771) );
  AO22X1 U4042 ( .IN1(N1017), .IN2(n3240), .IN3(N1976), .IN4(n3253), .Q(n4773)
         );
  OR2X1 U4043 ( .IN1(n4774), .IN2(n4775), .Q(n2635) );
  AO222X1 U4044 ( .IN1(rEIP_21_), .IN2(n2951), .IN3(N1052), .IN4(n3220), .IN5(
        n2956), .IN6(PhyAddrPointer_21_), .Q(n4775) );
  AO221X1 U4045 ( .IN1(n3227), .IN2(EBX_21_), .IN3(N1790), .IN4(n3233), .IN5(
        n4776), .Q(n4774) );
  AO22X1 U4046 ( .IN1(N1018), .IN2(n3240), .IN3(N1977), .IN4(n3253), .Q(n4776)
         );
  OR2X1 U4047 ( .IN1(n4777), .IN2(n4778), .Q(n2634) );
  AO222X1 U4048 ( .IN1(rEIP_22_), .IN2(n2952), .IN3(N1053), .IN4(n3219), .IN5(
        n2956), .IN6(PhyAddrPointer_22_), .Q(n4778) );
  AO221X1 U4049 ( .IN1(n3226), .IN2(EBX_22_), .IN3(N1791), .IN4(n3232), .IN5(
        n4779), .Q(n4777) );
  AO22X1 U4050 ( .IN1(N1019), .IN2(n3240), .IN3(N1978), .IN4(n3252), .Q(n4779)
         );
  OR2X1 U4051 ( .IN1(n4780), .IN2(n4781), .Q(n2633) );
  AO222X1 U4052 ( .IN1(rEIP_23_), .IN2(n2950), .IN3(N1054), .IN4(n3219), .IN5(
        n2956), .IN6(PhyAddrPointer_23_), .Q(n4781) );
  AO221X1 U4053 ( .IN1(n3226), .IN2(EBX_23_), .IN3(N1792), .IN4(n3232), .IN5(
        n4782), .Q(n4780) );
  AO22X1 U4054 ( .IN1(N1020), .IN2(n3240), .IN3(N1979), .IN4(n3252), .Q(n4782)
         );
  OR2X1 U4055 ( .IN1(n4783), .IN2(n4784), .Q(n2632) );
  AO222X1 U4056 ( .IN1(rEIP_24_), .IN2(n2951), .IN3(N1055), .IN4(n3219), .IN5(
        n2956), .IN6(test_so16), .Q(n4784) );
  AO221X1 U4057 ( .IN1(n3226), .IN2(EBX_24_), .IN3(N1793), .IN4(n3232), .IN5(
        n4785), .Q(n4783) );
  AO22X1 U4058 ( .IN1(N1021), .IN2(n3239), .IN3(N1980), .IN4(n3252), .Q(n4785)
         );
  OR2X1 U4059 ( .IN1(n4786), .IN2(n4787), .Q(n2631) );
  AO222X1 U4060 ( .IN1(rEIP_25_), .IN2(n2950), .IN3(N1056), .IN4(n3219), .IN5(
        n2956), .IN6(PhyAddrPointer_25_), .Q(n4787) );
  AO221X1 U4061 ( .IN1(n3226), .IN2(EBX_25_), .IN3(N1794), .IN4(n3232), .IN5(
        n4788), .Q(n4786) );
  AO22X1 U4062 ( .IN1(N1022), .IN2(n3239), .IN3(N1981), .IN4(n3252), .Q(n4788)
         );
  OR2X1 U4063 ( .IN1(n4789), .IN2(n4790), .Q(n2630) );
  AO222X1 U4064 ( .IN1(test_so19), .IN2(n2951), .IN3(N1057), .IN4(n3219), 
        .IN5(n2956), .IN6(PhyAddrPointer_26_), .Q(n4790) );
  AO221X1 U4065 ( .IN1(n3225), .IN2(EBX_26_), .IN3(N1795), .IN4(n3232), .IN5(
        n4791), .Q(n4789) );
  AO22X1 U4066 ( .IN1(N1023), .IN2(n3239), .IN3(N1982), .IN4(n3252), .Q(n4791)
         );
  OR2X1 U4067 ( .IN1(n4792), .IN2(n4793), .Q(n2629) );
  AO222X1 U4068 ( .IN1(rEIP_27_), .IN2(n2950), .IN3(N1058), .IN4(n3218), .IN5(
        n2956), .IN6(PhyAddrPointer_27_), .Q(n4793) );
  AO221X1 U4069 ( .IN1(n3225), .IN2(EBX_27_), .IN3(N1796), .IN4(n3231), .IN5(
        n4794), .Q(n4792) );
  AO22X1 U4070 ( .IN1(N1024), .IN2(n3239), .IN3(N1983), .IN4(n3251), .Q(n4794)
         );
  OR2X1 U4071 ( .IN1(n4795), .IN2(n4796), .Q(n2628) );
  AO222X1 U4072 ( .IN1(rEIP_28_), .IN2(n2951), .IN3(N1059), .IN4(n3218), .IN5(
        n2956), .IN6(PhyAddrPointer_28_), .Q(n4796) );
  AO221X1 U4073 ( .IN1(n3225), .IN2(EBX_28_), .IN3(N1797), .IN4(n3231), .IN5(
        n4797), .Q(n4795) );
  AO22X1 U4074 ( .IN1(N1025), .IN2(n3238), .IN3(N1984), .IN4(n3251), .Q(n4797)
         );
  OR2X1 U4075 ( .IN1(n4798), .IN2(n4799), .Q(n2627) );
  AO222X1 U4076 ( .IN1(rEIP_29_), .IN2(n2951), .IN3(N1060), .IN4(n3218), .IN5(
        n2956), .IN6(PhyAddrPointer_29_), .Q(n4799) );
  AO221X1 U4077 ( .IN1(n3225), .IN2(EBX_29_), .IN3(N1798), .IN4(n3231), .IN5(
        n4800), .Q(n4798) );
  AO22X1 U4078 ( .IN1(N1026), .IN2(n3238), .IN3(N1985), .IN4(n3251), .Q(n4800)
         );
  OR2X1 U4079 ( .IN1(n4801), .IN2(n4802), .Q(n2626) );
  AO222X1 U4080 ( .IN1(rEIP_30_), .IN2(n2951), .IN3(N1061), .IN4(n3218), .IN5(
        n2956), .IN6(PhyAddrPointer_30_), .Q(n4802) );
  AND3X1 U4081 ( .IN1(n4254), .IN2(n3103), .IN3(N1029), .Q(n4058) );
  AO221X1 U4082 ( .IN1(n3226), .IN2(EBX_30_), .IN3(N1799), .IN4(n3231), .IN5(
        n4803), .Q(n4801) );
  AO22X1 U4083 ( .IN1(N1027), .IN2(n3238), .IN3(N1986), .IN4(n3253), .Q(n4803)
         );
  AND4X1 U4084 ( .IN1(N1954), .IN2(n4804), .IN3(n4805), .IN4(n4806), .Q(n4063)
         );
  NOR3X0 U4085 ( .IN1(n2950), .IN2(N1029), .IN3(n4174), .QN(n4062) );
  AOI21X1 U4086 ( .IN1(n4102), .IN2(n4807), .IN3(n4699), .QN(n4060) );
  NAND2X0 U4087 ( .IN1(n4808), .IN2(n4805), .QN(n4807) );
  NAND3X0 U4088 ( .IN1(mult_add_463_aco_A_0_), .IN2(n4019), .IN3(n4808), .QN(
        n4102) );
  AOI21X1 U4089 ( .IN1(n4809), .IN2(n4810), .IN3(n4699), .QN(n4059) );
  INVX0 U4090 ( .IN(n4804), .QN(n4699) );
  NOR2X0 U4091 ( .IN1(n4091), .IN2(n2952), .QN(n4804) );
  OR3X1 U4092 ( .IN1(n4808), .IN2(N1954), .IN3(n4812), .Q(n4810) );
  AO21X1 U4093 ( .IN1(n4808), .IN2(n4019), .IN3(n4021), .Q(n4809) );
  INVX0 U4094 ( .IN(n4806), .QN(n4808) );
  NAND2X0 U4095 ( .IN1(n1472), .IN2(n2948), .QN(n4806) );
  AO222X1 U4096 ( .IN1(N499), .IN2(n3399), .IN3(n3211), .IN4(Address[0]), 
        .IN5(N426), .IN6(n3212), .Q(n2625) );
  AO222X1 U4097 ( .IN1(N500), .IN2(n3399), .IN3(n3210), .IN4(Address[1]), 
        .IN5(N427), .IN6(n3212), .Q(n2624) );
  AO222X1 U4098 ( .IN1(N501), .IN2(n3399), .IN3(n3210), .IN4(Address[2]), 
        .IN5(N428), .IN6(n3212), .Q(n2623) );
  AO222X1 U4099 ( .IN1(N502), .IN2(n3399), .IN3(n3210), .IN4(Address[3]), 
        .IN5(N429), .IN6(n3212), .Q(n2622) );
  AO222X1 U4100 ( .IN1(N503), .IN2(n3399), .IN3(n3210), .IN4(Address[4]), 
        .IN5(N430), .IN6(n3213), .Q(n2621) );
  AO222X1 U4101 ( .IN1(N504), .IN2(n3400), .IN3(n3210), .IN4(Address[5]), 
        .IN5(N431), .IN6(n3213), .Q(n2620) );
  AO222X1 U4102 ( .IN1(N505), .IN2(n3400), .IN3(n3208), .IN4(Address[6]), 
        .IN5(N432), .IN6(n3213), .Q(n2619) );
  AO222X1 U4103 ( .IN1(N506), .IN2(n3400), .IN3(n3210), .IN4(Address[7]), 
        .IN5(N433), .IN6(n3213), .Q(n2618) );
  AO222X1 U4104 ( .IN1(N507), .IN2(n3400), .IN3(n3209), .IN4(Address[8]), 
        .IN5(N434), .IN6(n3213), .Q(n2617) );
  AO222X1 U4105 ( .IN1(N508), .IN2(n3400), .IN3(n3209), .IN4(Address[9]), 
        .IN5(N435), .IN6(n3214), .Q(n2616) );
  AO222X1 U4106 ( .IN1(N509), .IN2(n3401), .IN3(n3209), .IN4(Address[10]), 
        .IN5(N436), .IN6(n3214), .Q(n2615) );
  AO222X1 U4107 ( .IN1(N510), .IN2(n3401), .IN3(n3209), .IN4(Address[11]), 
        .IN5(N437), .IN6(n3214), .Q(n2614) );
  AO222X1 U4108 ( .IN1(N511), .IN2(n3401), .IN3(n3209), .IN4(Address[12]), 
        .IN5(N438), .IN6(n3214), .Q(n2613) );
  AO222X1 U4109 ( .IN1(N512), .IN2(n3401), .IN3(n3209), .IN4(Address[13]), 
        .IN5(N439), .IN6(n3214), .Q(n2612) );
  AO222X1 U4110 ( .IN1(N513), .IN2(n3401), .IN3(n3208), .IN4(Address[14]), 
        .IN5(N440), .IN6(n3215), .Q(n2611) );
  AO222X1 U4111 ( .IN1(N514), .IN2(n3402), .IN3(n3208), .IN4(Address[15]), 
        .IN5(N441), .IN6(n3215), .Q(n2610) );
  AO222X1 U4112 ( .IN1(N515), .IN2(n3402), .IN3(n3208), .IN4(Address[16]), 
        .IN5(N442), .IN6(n3215), .Q(n2609) );
  AO222X1 U4113 ( .IN1(N516), .IN2(n3402), .IN3(n3208), .IN4(Address[17]), 
        .IN5(N443), .IN6(n3215), .Q(n2608) );
  AO222X1 U4114 ( .IN1(N517), .IN2(n3402), .IN3(n3208), .IN4(Address[18]), 
        .IN5(N444), .IN6(n3215), .Q(n2607) );
  AO222X1 U4115 ( .IN1(N518), .IN2(n3402), .IN3(n3207), .IN4(Address[19]), 
        .IN5(N445), .IN6(n3216), .Q(n2606) );
  AO222X1 U4116 ( .IN1(N519), .IN2(n3403), .IN3(n3207), .IN4(Address[20]), 
        .IN5(N446), .IN6(n3216), .Q(n2605) );
  AO222X1 U4117 ( .IN1(N520), .IN2(n3403), .IN3(n3207), .IN4(Address[21]), 
        .IN5(N447), .IN6(n3216), .Q(n2604) );
  AO222X1 U4118 ( .IN1(N521), .IN2(n3403), .IN3(n3207), .IN4(Address[22]), 
        .IN5(N448), .IN6(n3216), .Q(n2603) );
  AO222X1 U4119 ( .IN1(N522), .IN2(n3403), .IN3(n3207), .IN4(Address[23]), 
        .IN5(N449), .IN6(n3216), .Q(n2602) );
  AO222X1 U4120 ( .IN1(N523), .IN2(n3403), .IN3(n3207), .IN4(Address[24]), 
        .IN5(N450), .IN6(n3217), .Q(n2601) );
  AO222X1 U4121 ( .IN1(N524), .IN2(n3404), .IN3(n3206), .IN4(Address[25]), 
        .IN5(N451), .IN6(n3217), .Q(n2600) );
  AO222X1 U4122 ( .IN1(N525), .IN2(n3404), .IN3(n3206), .IN4(Address[26]), 
        .IN5(N452), .IN6(n3217), .Q(n2599) );
  AO222X1 U4123 ( .IN1(N526), .IN2(n3404), .IN3(n3206), .IN4(Address[27]), 
        .IN5(N453), .IN6(n3217), .Q(n2598) );
  AO222X1 U4124 ( .IN1(N527), .IN2(n3404), .IN3(n3206), .IN4(Address[28]), 
        .IN5(N454), .IN6(n3217), .Q(n2597) );
  AO222X1 U4125 ( .IN1(N528), .IN2(n3404), .IN3(n3205), .IN4(Address[29]), 
        .IN5(N455), .IN6(n3217), .Q(n2596) );
  INVX0 U4126 ( .IN(n4814), .QN(n4049) );
  INVX0 U4127 ( .IN(n4030), .QN(n4813) );
  MUX21X1 U4128 ( .IN1(n4815), .IN2(n4816), .S(n4817), .Q(n2595) );
  NAND2X0 U4129 ( .IN1(n4818), .IN2(n4148), .QN(n4815) );
  MUX21X1 U4130 ( .IN1(n1595), .IN2(W_R_n), .S(n3206), .Q(n2594) );
  MUX21X1 U4131 ( .IN1(n4819), .IN2(n4820), .S(n4817), .Q(n2593) );
  INVX0 U4132 ( .IN(n4011), .QN(n4817) );
  NAND3X0 U4133 ( .IN1(n4115), .IN2(n3185), .IN3(n4811), .QN(n4011) );
  NAND2X0 U4134 ( .IN1(n4818), .IN2(n4021), .QN(n4819) );
  NOR3X0 U4135 ( .IN1(n4112), .IN2(n3196), .IN3(n4805), .QN(n4818) );
  MUX21X1 U4136 ( .IN1(n4820), .IN2(M_IO_n), .S(n3205), .Q(n2592) );
  AO21X1 U4137 ( .IN1(n4811), .IN2(n4821), .IN3(n4112), .Q(n2591) );
  INVX0 U4138 ( .IN(n4115), .QN(n4112) );
  NAND2X0 U4139 ( .IN1(n4116), .IN2(n4649), .QN(n4115) );
  NAND3X0 U4140 ( .IN1(n4017), .IN2(n4660), .IN3(n4651), .QN(n4811) );
  OR3X1 U4141 ( .IN1(n4805), .IN2(mult_add_463_aco_A_0_), .IN3(n4698), .Q(
        n4660) );
  NAND2X0 U4142 ( .IN1(n4822), .IN2(n4148), .QN(n4698) );
  NAND2X0 U4143 ( .IN1(n4823), .IN2(n4044), .QN(n2590) );
  NAND3X0 U4144 ( .IN1(n1436), .IN2(n1434), .IN3(n1435), .QN(n4044) );
  MUX21X1 U4145 ( .IN1(n4821), .IN2(n3872), .S(n3205), .Q(n4823) );
  AO222X1 U4146 ( .IN1(Datai[15]), .IN2(n3408), .IN3(n3411), .IN4(N3361), 
        .IN5(n3417), .IN6(N3449), .Q(n2589) );
  AO221X1 U4147 ( .IN1(N1551), .IN2(n3424), .IN3(n3434), .IN4(N3346), .IN5(
        n4829), .Q(n2588) );
  AO222X1 U4148 ( .IN1(N2385), .IN2(n3441), .IN3(N2103), .IN4(n3453), .IN5(
        n3465), .IN6(n3080), .Q(n4829) );
  AO221X1 U4149 ( .IN1(N1552), .IN2(n3424), .IN3(n3437), .IN4(N3347), .IN5(
        n4833), .Q(n2587) );
  AO222X1 U4150 ( .IN1(N2386), .IN2(n3441), .IN3(N2104), .IN4(n3453), .IN5(
        n3465), .IN6(Datai[1]), .Q(n4833) );
  AO221X1 U4151 ( .IN1(N1553), .IN2(n3424), .IN3(n3436), .IN4(N3348), .IN5(
        n4834), .Q(n2586) );
  AO222X1 U4152 ( .IN1(N2387), .IN2(n3441), .IN3(N2105), .IN4(n3453), .IN5(
        n3465), .IN6(n3084), .Q(n4834) );
  AO221X1 U4153 ( .IN1(N1554), .IN2(n3424), .IN3(n3436), .IN4(N3349), .IN5(
        n4835), .Q(n2585) );
  AO222X1 U4154 ( .IN1(N2388), .IN2(n3441), .IN3(N2106), .IN4(n3453), .IN5(
        n3465), .IN6(Datai[3]), .Q(n4835) );
  AO221X1 U4155 ( .IN1(N1555), .IN2(n3424), .IN3(n3436), .IN4(N3350), .IN5(
        n4836), .Q(n2584) );
  AO222X1 U4156 ( .IN1(N2389), .IN2(n3441), .IN3(N2107), .IN4(n3453), .IN5(
        n3466), .IN6(Datai[4]), .Q(n4836) );
  AO221X1 U4157 ( .IN1(N1556), .IN2(n3425), .IN3(n3436), .IN4(N3351), .IN5(
        n4837), .Q(n2583) );
  AO222X1 U4158 ( .IN1(N2390), .IN2(n3442), .IN3(N2108), .IN4(n3454), .IN5(
        n3466), .IN6(Datai[5]), .Q(n4837) );
  AO221X1 U4159 ( .IN1(N1557), .IN2(n3425), .IN3(n3436), .IN4(N3352), .IN5(
        n4838), .Q(n2582) );
  AO222X1 U4160 ( .IN1(N2391), .IN2(n3442), .IN3(N2109), .IN4(n3454), .IN5(
        n3466), .IN6(n3092), .Q(n4838) );
  AO221X1 U4161 ( .IN1(N1558), .IN2(n3425), .IN3(n3435), .IN4(N3353), .IN5(
        n4839), .Q(n2581) );
  AO222X1 U4162 ( .IN1(N2392), .IN2(n3442), .IN3(N2110), .IN4(n3454), .IN5(
        n3466), .IN6(n3094), .Q(n4839) );
  AO221X1 U4163 ( .IN1(N1559), .IN2(n3425), .IN3(n3435), .IN4(N3354), .IN5(
        n4840), .Q(n2580) );
  AO222X1 U4164 ( .IN1(N2393), .IN2(n3442), .IN3(N2111), .IN4(n3454), .IN5(
        n2941), .IN6(n3467), .Q(n4840) );
  AO221X1 U4165 ( .IN1(N1560), .IN2(n3425), .IN3(n3435), .IN4(test_so4), .IN5(
        n4841), .Q(n2579) );
  AO222X1 U4166 ( .IN1(N2394), .IN2(n3442), .IN3(N2112), .IN4(n3454), .IN5(
        n2945), .IN6(n3471), .Q(n4841) );
  AO221X1 U4167 ( .IN1(N1561), .IN2(n3426), .IN3(n3435), .IN4(N3356), .IN5(
        n4842), .Q(n2578) );
  AO222X1 U4168 ( .IN1(N2395), .IN2(n3443), .IN3(N2113), .IN4(n3455), .IN5(
        n2937), .IN6(n3471), .Q(n4842) );
  AO221X1 U4169 ( .IN1(N1562), .IN2(n3426), .IN3(n3435), .IN4(N3357), .IN5(
        n4843), .Q(n2577) );
  AO222X1 U4170 ( .IN1(N2396), .IN2(n3443), .IN3(N2114), .IN4(n3455), .IN5(
        n2943), .IN6(n3470), .Q(n4843) );
  AO221X1 U4171 ( .IN1(N1563), .IN2(n3426), .IN3(n3434), .IN4(N3358), .IN5(
        n4844), .Q(n2576) );
  AO222X1 U4172 ( .IN1(N2397), .IN2(n3443), .IN3(N2115), .IN4(n3455), .IN5(
        n2947), .IN6(n3470), .Q(n4844) );
  AO221X1 U4173 ( .IN1(N1564), .IN2(n3426), .IN3(n3434), .IN4(N3359), .IN5(
        n4845), .Q(n2575) );
  AO222X1 U4174 ( .IN1(N2398), .IN2(n3443), .IN3(N2116), .IN4(n3455), .IN5(
        n2935), .IN6(n3470), .Q(n4845) );
  AO221X1 U4175 ( .IN1(N1565), .IN2(n3426), .IN3(n3434), .IN4(N3360), .IN5(
        n4846), .Q(n2574) );
  AO222X1 U4176 ( .IN1(N2399), .IN2(n3443), .IN3(N2117), .IN4(n3455), .IN5(
        n2939), .IN6(n3470), .Q(n4846) );
  AO221X1 U4177 ( .IN1(N1566), .IN2(n3427), .IN3(n3434), .IN4(N3361), .IN5(
        n4847), .Q(n2573) );
  AO222X1 U4178 ( .IN1(N2400), .IN2(n3444), .IN3(N2118), .IN4(n3456), .IN5(
        n3466), .IN6(Datai[15]), .Q(n4847) );
  AO222X1 U4179 ( .IN1(n3405), .IN2(n3080), .IN3(n3411), .IN4(N3346), .IN5(
        n3417), .IN6(N3434), .Q(n2572) );
  AO222X1 U4180 ( .IN1(n3405), .IN2(n3082), .IN3(n3411), .IN4(N3347), .IN5(
        n3417), .IN6(N3435), .Q(n2571) );
  AO222X1 U4181 ( .IN1(n3405), .IN2(n3084), .IN3(n3411), .IN4(N3348), .IN5(
        n3417), .IN6(test_so17), .Q(n2570) );
  AO222X1 U4182 ( .IN1(n3405), .IN2(n3086), .IN3(n3411), .IN4(N3349), .IN5(
        n3417), .IN6(N3437), .Q(n2569) );
  AO222X1 U4183 ( .IN1(n3405), .IN2(n3088), .IN3(n3412), .IN4(N3350), .IN5(
        n3418), .IN6(N3438), .Q(n2568) );
  AO222X1 U4184 ( .IN1(n3406), .IN2(n3090), .IN3(n3412), .IN4(N3351), .IN5(
        n3418), .IN6(N3439), .Q(n2567) );
  AO222X1 U4185 ( .IN1(n3406), .IN2(n3092), .IN3(n3412), .IN4(N3352), .IN5(
        n3418), .IN6(N3440), .Q(n2566) );
  AO222X1 U4186 ( .IN1(n3406), .IN2(n3094), .IN3(n3412), .IN4(N3353), .IN5(
        n3418), .IN6(N3441), .Q(n2565) );
  AO222X1 U4187 ( .IN1(n2941), .IN2(n3409), .IN3(n3412), .IN4(N3354), .IN5(
        n3418), .IN6(N3442), .Q(n2564) );
  AO222X1 U4188 ( .IN1(n2945), .IN2(n3410), .IN3(n3413), .IN4(test_so4), .IN5(
        n3419), .IN6(N3443), .Q(n2563) );
  AO222X1 U4189 ( .IN1(n2937), .IN2(n3410), .IN3(n3413), .IN4(N3356), .IN5(
        n3419), .IN6(N3444), .Q(n2562) );
  AO222X1 U4190 ( .IN1(n2943), .IN2(n3410), .IN3(n3413), .IN4(N3357), .IN5(
        n3419), .IN6(N3445), .Q(n2561) );
  AO222X1 U4191 ( .IN1(n2947), .IN2(n3410), .IN3(n3413), .IN4(N3358), .IN5(
        n3419), .IN6(N3446), .Q(n2560) );
  AO222X1 U4192 ( .IN1(n2935), .IN2(n3410), .IN3(n3413), .IN4(N3359), .IN5(
        n3419), .IN6(N3447), .Q(n2559) );
  AO222X1 U4193 ( .IN1(n2939), .IN2(n3409), .IN3(n3414), .IN4(N3360), .IN5(
        n3420), .IN6(N3448), .Q(n2558) );
  AO221X1 U4194 ( .IN1(N1567), .IN2(n3427), .IN3(n3433), .IN4(EAX_16_), .IN5(
        n4848), .Q(n2557) );
  AO222X1 U4195 ( .IN1(N2401), .IN2(n3444), .IN3(Datai[0]), .IN4(n3456), .IN5(
        Datai[16]), .IN6(n3470), .Q(n4848) );
  AO221X1 U4196 ( .IN1(N1568), .IN2(n3427), .IN3(n3433), .IN4(EAX_17_), .IN5(
        n4849), .Q(n2556) );
  AO222X1 U4197 ( .IN1(N2402), .IN2(n3444), .IN3(n3082), .IN4(n3456), .IN5(
        Datai[17]), .IN6(n3469), .Q(n4849) );
  AO221X1 U4198 ( .IN1(N1569), .IN2(n3427), .IN3(n3433), .IN4(EAX_18_), .IN5(
        n4850), .Q(n2555) );
  AO222X1 U4199 ( .IN1(N2403), .IN2(n3444), .IN3(Datai[2]), .IN4(n3456), .IN5(
        Datai[18]), .IN6(n3469), .Q(n4850) );
  AO221X1 U4200 ( .IN1(N1570), .IN2(n3427), .IN3(n3433), .IN4(EAX_19_), .IN5(
        n4851), .Q(n2554) );
  AO222X1 U4201 ( .IN1(N2404), .IN2(n3444), .IN3(Datai[3]), .IN4(n3456), .IN5(
        Datai[19]), .IN6(n3469), .Q(n4851) );
  AO221X1 U4202 ( .IN1(N1571), .IN2(n3428), .IN3(n3433), .IN4(EAX_20_), .IN5(
        n4852), .Q(n2553) );
  AO222X1 U4203 ( .IN1(N2405), .IN2(n3445), .IN3(Datai[4]), .IN4(n3457), .IN5(
        Datai[20]), .IN6(n3469), .Q(n4852) );
  AO221X1 U4204 ( .IN1(N1572), .IN2(n3428), .IN3(n3432), .IN4(EAX_21_), .IN5(
        n4853), .Q(n2552) );
  AO222X1 U4205 ( .IN1(N2406), .IN2(n3445), .IN3(n3090), .IN4(n3457), .IN5(
        Datai[21]), .IN6(n3468), .Q(n4853) );
  AO221X1 U4206 ( .IN1(N1573), .IN2(n3428), .IN3(n3432), .IN4(EAX_22_), .IN5(
        n4854), .Q(n2551) );
  AO222X1 U4207 ( .IN1(N2407), .IN2(n3445), .IN3(Datai[6]), .IN4(n3457), .IN5(
        Datai[22]), .IN6(n3468), .Q(n4854) );
  AO221X1 U4208 ( .IN1(N1574), .IN2(n3428), .IN3(n3432), .IN4(EAX_23_), .IN5(
        n4855), .Q(n2550) );
  AO222X1 U4209 ( .IN1(N2408), .IN2(n3445), .IN3(Datai[7]), .IN4(n3457), .IN5(
        Datai[23]), .IN6(n3469), .Q(n4855) );
  AO221X1 U4210 ( .IN1(N1575), .IN2(n3428), .IN3(n3432), .IN4(EAX_24_), .IN5(
        n4856), .Q(n2549) );
  AO222X1 U4211 ( .IN1(N2409), .IN2(n3445), .IN3(n2941), .IN4(n3457), .IN5(
        Datai[24]), .IN6(n3468), .Q(n4856) );
  AO221X1 U4212 ( .IN1(N1576), .IN2(n3429), .IN3(n3432), .IN4(EAX_25_), .IN5(
        n4857), .Q(n2548) );
  AO222X1 U4213 ( .IN1(N2410), .IN2(n3446), .IN3(n2945), .IN4(n3458), .IN5(
        Datai[25]), .IN6(n3468), .Q(n4857) );
  AO221X1 U4214 ( .IN1(N1577), .IN2(n3429), .IN3(n3431), .IN4(EAX_26_), .IN5(
        n4858), .Q(n2547) );
  AO222X1 U4215 ( .IN1(N2411), .IN2(n3446), .IN3(n2937), .IN4(n3458), .IN5(
        Datai[26]), .IN6(n3468), .Q(n4858) );
  AO221X1 U4216 ( .IN1(N1578), .IN2(n3429), .IN3(n3431), .IN4(EAX_27_), .IN5(
        n4859), .Q(n2546) );
  AO222X1 U4217 ( .IN1(N2412), .IN2(n3446), .IN3(n2943), .IN4(n3458), .IN5(
        Datai[27]), .IN6(n3467), .Q(n4859) );
  AO221X1 U4218 ( .IN1(N1579), .IN2(n3429), .IN3(n3431), .IN4(EAX_28_), .IN5(
        n4860), .Q(n2545) );
  AO222X1 U4219 ( .IN1(N2413), .IN2(n3446), .IN3(n2947), .IN4(n3458), .IN5(
        Datai[28]), .IN6(n3467), .Q(n4860) );
  AO221X1 U4220 ( .IN1(N1580), .IN2(n3429), .IN3(n3431), .IN4(EAX_29_), .IN5(
        n4861), .Q(n2544) );
  AO222X1 U4221 ( .IN1(N2414), .IN2(n3446), .IN3(n2935), .IN4(n3458), .IN5(
        Datai[29]), .IN6(n3467), .Q(n4861) );
  AO221X1 U4222 ( .IN1(N1581), .IN2(n3430), .IN3(n3431), .IN4(test_so5), .IN5(
        n4862), .Q(n2543) );
  AO222X1 U4223 ( .IN1(N2415), .IN2(n3447), .IN3(n2939), .IN4(n3459), .IN5(
        Datai[30]), .IN6(n3467), .Q(n4862) );
  NOR2X0 U4224 ( .IN1(n3437), .IN2(n4812), .QN(n4831) );
  NOR2X0 U4225 ( .IN1(n3437), .IN2(n4863), .QN(n4830) );
  AO222X1 U4226 ( .IN1(N1582), .IN2(n3430), .IN3(n3465), .IN4(Datai[31]), 
        .IN5(n3437), .IN6(EAX_31_), .Q(n2542) );
  NOR2X0 U4227 ( .IN1(n3437), .IN2(n4148), .QN(n4832) );
  ISOLANDX1 U4228 ( .D(n4864), .ISO(n3439), .Q(n4827) );
  NAND2X0 U4229 ( .IN1(n4017), .IN2(n4865), .QN(n4828) );
  AO221X1 U4230 ( .IN1(n4866), .IN2(n4651), .IN3(n4867), .IN4(n4868), .IN5(
        n4864), .Q(n4865) );
  INVX0 U4231 ( .IN(n4863), .QN(n4867) );
  ISOLANDX1 U4232 ( .D(n4869), .ISO(n2949), .Q(n4866) );
  AND4X1 U4233 ( .IN1(n4870), .IN2(n4125), .IN3(n4124), .IN4(n4871), .Q(n4864)
         );
  NOR2X0 U4234 ( .IN1(n4628), .IN2(n4129), .QN(n4871) );
  AO222X1 U4235 ( .IN1(n3407), .IN2(n3080), .IN3(N1750), .IN4(n3414), .IN5(
        N3450), .IN6(n3421), .Q(n2541) );
  AO222X1 U4236 ( .IN1(n3407), .IN2(n3082), .IN3(N1751), .IN4(n3414), .IN5(
        N3451), .IN6(n3423), .Q(n2540) );
  AO222X1 U4237 ( .IN1(n3406), .IN2(n3084), .IN3(N1752), .IN4(n3414), .IN5(
        N3452), .IN6(n3423), .Q(n2539) );
  AO222X1 U4238 ( .IN1(n3407), .IN2(n3086), .IN3(N1753), .IN4(n3414), .IN5(
        N3453), .IN6(n3423), .Q(n2538) );
  AO222X1 U4239 ( .IN1(n3407), .IN2(n3088), .IN3(N1754), .IN4(n3415), .IN5(
        N3454), .IN6(n3422), .Q(n2537) );
  AO222X1 U4240 ( .IN1(n3408), .IN2(n3090), .IN3(N1755), .IN4(n3415), .IN5(
        N3455), .IN6(n3422), .Q(n2536) );
  AO222X1 U4241 ( .IN1(n3406), .IN2(n3092), .IN3(N1756), .IN4(n3415), .IN5(
        N3456), .IN6(n3422), .Q(n2535) );
  AO222X1 U4242 ( .IN1(n3407), .IN2(n3094), .IN3(N1757), .IN4(n3415), .IN5(
        N3457), .IN6(n3422), .Q(n2534) );
  AO222X1 U4243 ( .IN1(n2941), .IN2(n3409), .IN3(N1758), .IN4(n3415), .IN5(
        N3458), .IN6(n3422), .Q(n2533) );
  AO222X1 U4244 ( .IN1(n2945), .IN2(n3408), .IN3(N1759), .IN4(n3416), .IN5(
        N3459), .IN6(n3421), .Q(n2532) );
  AO222X1 U4245 ( .IN1(n2937), .IN2(n3409), .IN3(N1760), .IN4(n3416), .IN5(
        N3460), .IN6(n3421), .Q(n2531) );
  AO222X1 U4246 ( .IN1(n2943), .IN2(n3408), .IN3(N1761), .IN4(n3416), .IN5(
        N3461), .IN6(n3421), .Q(n2530) );
  AO222X1 U4247 ( .IN1(n2947), .IN2(n3409), .IN3(N1762), .IN4(n3416), .IN5(
        N3462), .IN6(n3421), .Q(n2529) );
  AO222X1 U4248 ( .IN1(n2935), .IN2(n3408), .IN3(N1763), .IN4(n3416), .IN5(
        N3463), .IN6(n3420), .Q(n2528) );
  AO222X1 U4249 ( .IN1(n2939), .IN2(n3409), .IN3(N1764), .IN4(n3413), .IN5(
        test_so20), .IN6(n3420), .Q(n2527) );
  NOR2X0 U4250 ( .IN1(n3420), .IN2(n4021), .QN(n4825) );
  NOR2X0 U4251 ( .IN1(n3420), .IN2(n4812), .QN(n4824) );
  NAND3X0 U4252 ( .IN1(n4017), .IN2(n4872), .IN3(n4651), .QN(n4826) );
  AO21X1 U4253 ( .IN1(n4805), .IN2(n2948), .IN3(mult_add_463_aco_A_0_), .Q(
        n4872) );
  INVX0 U4254 ( .IN(n4812), .QN(n4805) );
  NAND4X0 U4255 ( .IN1(n4873), .IN2(n4874), .IN3(n4875), .IN4(n4876), .QN(
        n2526) );
  OA22X1 U4256 ( .IN1(n3257), .IN2(n4877), .IN3(n3264), .IN4(n4878), .Q(n4876)
         );
  AOI22X1 U4257 ( .IN1(N1479), .IN2(n3276), .IN3(n65), .IN4(n3288), .QN(n4875)
         );
  AOI22X1 U4258 ( .IN1(N2856), .IN2(n3300), .IN3(N2416), .IN4(n3312), .QN(
        n4874) );
  OA22X1 U4259 ( .IN1(n1557), .IN2(n3331), .IN3(n3188), .IN4(n2845), .Q(n4873)
         );
  NAND4X0 U4260 ( .IN1(n4879), .IN2(n4880), .IN3(n4881), .IN4(n4882), .QN(
        n2525) );
  OA22X1 U4261 ( .IN1(n3257), .IN2(n4883), .IN3(n3264), .IN4(n4884), .Q(n4882)
         );
  AOI22X1 U4262 ( .IN1(N1480), .IN2(n3276), .IN3(n64), .IN4(n3288), .QN(n4881)
         );
  AOI22X1 U4263 ( .IN1(N2857), .IN2(n3300), .IN3(N2417), .IN4(n3312), .QN(
        n4880) );
  OA22X1 U4264 ( .IN1(n3867), .IN2(n3331), .IN3(n3188), .IN4(n2888), .Q(n4879)
         );
  NAND4X0 U4265 ( .IN1(n4885), .IN2(n4886), .IN3(n4887), .IN4(n4888), .QN(
        n2524) );
  OA22X1 U4266 ( .IN1(n3257), .IN2(n4889), .IN3(n3264), .IN4(n4890), .Q(n4888)
         );
  AOI22X1 U4267 ( .IN1(N1481), .IN2(n3276), .IN3(n63), .IN4(n3288), .QN(n4887)
         );
  AOI22X1 U4268 ( .IN1(N2858), .IN2(n3300), .IN3(N2418), .IN4(n3312), .QN(
        n4886) );
  OA22X1 U4269 ( .IN1(n3866), .IN2(n3331), .IN3(n3188), .IN4(n4680), .Q(n4885)
         );
  NAND4X0 U4270 ( .IN1(n4891), .IN2(n4892), .IN3(n4893), .IN4(n4894), .QN(
        n2523) );
  OA22X1 U4271 ( .IN1(n3257), .IN2(n4895), .IN3(n3265), .IN4(n4896), .Q(n4894)
         );
  AOI22X1 U4272 ( .IN1(N1482), .IN2(n3277), .IN3(n62), .IN4(n3289), .QN(n4893)
         );
  AOI22X1 U4273 ( .IN1(N2859), .IN2(n3301), .IN3(N2419), .IN4(n3313), .QN(
        n4892) );
  OA22X1 U4274 ( .IN1(n3865), .IN2(n3331), .IN3(n3189), .IN4(n4686), .Q(n4891)
         );
  NAND4X0 U4275 ( .IN1(n4897), .IN2(n4898), .IN3(n4899), .IN4(n4900), .QN(
        n2522) );
  OA22X1 U4276 ( .IN1(n3258), .IN2(n4901), .IN3(n3265), .IN4(n4902), .Q(n4900)
         );
  AOI22X1 U4277 ( .IN1(N1483), .IN2(n3277), .IN3(n61), .IN4(n3289), .QN(n4899)
         );
  AOI22X1 U4278 ( .IN1(N2860), .IN2(n3301), .IN3(N2420), .IN4(n3313), .QN(
        n4898) );
  OA22X1 U4279 ( .IN1(n3864), .IN2(n3330), .IN3(n3189), .IN4(n4692), .Q(n4897)
         );
  NAND4X0 U4280 ( .IN1(n4903), .IN2(n4904), .IN3(n4905), .IN4(n4906), .QN(
        n2521) );
  OA22X1 U4281 ( .IN1(n3258), .IN2(n4907), .IN3(n3265), .IN4(n4908), .Q(n4906)
         );
  AOI22X1 U4282 ( .IN1(N1484), .IN2(n3277), .IN3(n60), .IN4(n3289), .QN(n4905)
         );
  AOI22X1 U4283 ( .IN1(N2861), .IN2(n3301), .IN3(N2421), .IN4(n3313), .QN(
        n4904) );
  OA22X1 U4284 ( .IN1(n3870), .IN2(n3330), .IN3(n3189), .IN4(n4700), .Q(n4903)
         );
  NAND4X0 U4285 ( .IN1(n4909), .IN2(n4910), .IN3(n4911), .IN4(n4912), .QN(
        n2520) );
  OA22X1 U4286 ( .IN1(n3258), .IN2(n4913), .IN3(n3265), .IN4(n4914), .Q(n4912)
         );
  AOI22X1 U4287 ( .IN1(N1485), .IN2(n3277), .IN3(n59), .IN4(n3289), .QN(n4911)
         );
  AOI22X1 U4288 ( .IN1(N2862), .IN2(n3301), .IN3(N2422), .IN4(n3313), .QN(
        n4910) );
  OA22X1 U4289 ( .IN1(n3863), .IN2(n3330), .IN3(n3189), .IN4(n4704), .Q(n4909)
         );
  NAND4X0 U4290 ( .IN1(n4915), .IN2(n4916), .IN3(n4917), .IN4(n4918), .QN(
        n2519) );
  OA22X1 U4291 ( .IN1(n3258), .IN2(n4919), .IN3(n3266), .IN4(n4920), .Q(n4918)
         );
  AOI22X1 U4292 ( .IN1(N1486), .IN2(n3278), .IN3(n58), .IN4(n3290), .QN(n4917)
         );
  AOI22X1 U4293 ( .IN1(N2863), .IN2(n3302), .IN3(N2423), .IN4(n3314), .QN(
        n4916) );
  OA22X1 U4294 ( .IN1(n3862), .IN2(n3330), .IN3(n3190), .IN4(n4709), .Q(n4915)
         );
  NAND4X0 U4295 ( .IN1(n4921), .IN2(n4922), .IN3(n4923), .IN4(n4924), .QN(
        n2518) );
  OA22X1 U4296 ( .IN1(n3258), .IN2(n4925), .IN3(n3266), .IN4(n4926), .Q(n4924)
         );
  AOI22X1 U4297 ( .IN1(N1487), .IN2(n3278), .IN3(n57), .IN4(n3290), .QN(n4923)
         );
  AOI22X1 U4298 ( .IN1(N2864), .IN2(n3302), .IN3(N2424), .IN4(n3314), .QN(
        n4922) );
  OA22X1 U4299 ( .IN1(n3861), .IN2(n3329), .IN3(n3190), .IN4(n4714), .Q(n4921)
         );
  NAND4X0 U4300 ( .IN1(n4927), .IN2(n4928), .IN3(n4929), .IN4(n4930), .QN(
        n2517) );
  OA22X1 U4301 ( .IN1(n3259), .IN2(n4931), .IN3(n3266), .IN4(n4932), .Q(n4930)
         );
  AOI22X1 U4302 ( .IN1(N1488), .IN2(n3278), .IN3(n56), .IN4(n3290), .QN(n4929)
         );
  AOI22X1 U4303 ( .IN1(N2865), .IN2(n3302), .IN3(N2425), .IN4(n3314), .QN(
        n4928) );
  OA22X1 U4304 ( .IN1(n3860), .IN2(n3329), .IN3(n3190), .IN4(n4719), .Q(n4927)
         );
  NAND4X0 U4305 ( .IN1(n4933), .IN2(n4934), .IN3(n4935), .IN4(n4936), .QN(
        n2516) );
  OA22X1 U4306 ( .IN1(n3259), .IN2(n4937), .IN3(n3266), .IN4(n4938), .Q(n4936)
         );
  AOI22X1 U4307 ( .IN1(N1489), .IN2(n3278), .IN3(n55), .IN4(n3290), .QN(n4935)
         );
  AOI22X1 U4308 ( .IN1(N2866), .IN2(n3302), .IN3(N2426), .IN4(n3314), .QN(
        n4934) );
  OA22X1 U4309 ( .IN1(n3859), .IN2(n3329), .IN3(n3190), .IN4(n4724), .Q(n4933)
         );
  NAND4X0 U4310 ( .IN1(n4939), .IN2(n4940), .IN3(n4941), .IN4(n4942), .QN(
        n2515) );
  OA22X1 U4311 ( .IN1(n3259), .IN2(n4943), .IN3(n3267), .IN4(n4944), .Q(n4942)
         );
  AOI22X1 U4312 ( .IN1(N1490), .IN2(n3279), .IN3(n54), .IN4(n3291), .QN(n4941)
         );
  AOI22X1 U4313 ( .IN1(N2867), .IN2(n3303), .IN3(N2427), .IN4(n3315), .QN(
        n4940) );
  OA22X1 U4314 ( .IN1(n3858), .IN2(n3329), .IN3(n3190), .IN4(n4729), .Q(n4939)
         );
  NAND4X0 U4315 ( .IN1(n4945), .IN2(n4946), .IN3(n4947), .IN4(n4948), .QN(
        n2514) );
  OA22X1 U4316 ( .IN1(n3259), .IN2(n4949), .IN3(n3267), .IN4(n4950), .Q(n4948)
         );
  AOI22X1 U4317 ( .IN1(N1491), .IN2(n3279), .IN3(n53), .IN4(n3291), .QN(n4947)
         );
  AOI22X1 U4318 ( .IN1(N2868), .IN2(n3303), .IN3(N2428), .IN4(n3315), .QN(
        n4946) );
  OA22X1 U4319 ( .IN1(n3857), .IN2(n3328), .IN3(n3191), .IN4(n4734), .Q(n4945)
         );
  NAND4X0 U4320 ( .IN1(n4951), .IN2(n4952), .IN3(n4953), .IN4(n4954), .QN(
        n2513) );
  OA22X1 U4321 ( .IN1(n3259), .IN2(n4955), .IN3(n3267), .IN4(n4956), .Q(n4954)
         );
  AOI22X1 U4322 ( .IN1(N1492), .IN2(n3279), .IN3(n52), .IN4(n3291), .QN(n4953)
         );
  AOI22X1 U4323 ( .IN1(N2869), .IN2(n3303), .IN3(N2429), .IN4(n3315), .QN(
        n4952) );
  OA22X1 U4324 ( .IN1(n3856), .IN2(n3328), .IN3(n3191), .IN4(n4739), .Q(n4951)
         );
  NAND4X0 U4325 ( .IN1(n4957), .IN2(n4958), .IN3(n4959), .IN4(n4960), .QN(
        n2512) );
  OA22X1 U4326 ( .IN1(n3260), .IN2(n4961), .IN3(n3267), .IN4(n4962), .Q(n4960)
         );
  AOI22X1 U4327 ( .IN1(N1493), .IN2(n3279), .IN3(n51), .IN4(n3291), .QN(n4959)
         );
  AOI22X1 U4328 ( .IN1(N2870), .IN2(n3303), .IN3(N2430), .IN4(n3315), .QN(
        n4958) );
  OA22X1 U4329 ( .IN1(n3855), .IN2(n3328), .IN3(n3191), .IN4(n4744), .Q(n4957)
         );
  NAND4X0 U4330 ( .IN1(n4963), .IN2(n4964), .IN3(n4965), .IN4(n4966), .QN(
        n2511) );
  OA22X1 U4331 ( .IN1(n3260), .IN2(n4967), .IN3(n3268), .IN4(n4968), .Q(n4966)
         );
  AOI22X1 U4332 ( .IN1(N1494), .IN2(n3280), .IN3(n50), .IN4(n3292), .QN(n4965)
         );
  AOI22X1 U4333 ( .IN1(N2871), .IN2(n3304), .IN3(N2431), .IN4(n3316), .QN(
        n4964) );
  OA22X1 U4334 ( .IN1(n3854), .IN2(n3327), .IN3(n3191), .IN4(n4749), .Q(n4963)
         );
  NAND4X0 U4335 ( .IN1(n4969), .IN2(n4970), .IN3(n4971), .IN4(n4972), .QN(
        n2510) );
  OA22X1 U4336 ( .IN1(n3260), .IN2(n4973), .IN3(n3268), .IN4(n4974), .Q(n4972)
         );
  AOI22X1 U4337 ( .IN1(N1495), .IN2(n3280), .IN3(n49), .IN4(n3292), .QN(n4971)
         );
  AOI22X1 U4338 ( .IN1(N2872), .IN2(n3304), .IN3(N2432), .IN4(n3316), .QN(
        n4970) );
  OA22X1 U4339 ( .IN1(n3853), .IN2(n3327), .IN3(n3191), .IN4(n4754), .Q(n4969)
         );
  NAND4X0 U4340 ( .IN1(n4975), .IN2(n4976), .IN3(n4977), .IN4(n4978), .QN(
        n2509) );
  OA22X1 U4341 ( .IN1(n3260), .IN2(n4979), .IN3(n3268), .IN4(n4980), .Q(n4978)
         );
  AOI22X1 U4342 ( .IN1(N1496), .IN2(n3280), .IN3(n48), .IN4(n3292), .QN(n4977)
         );
  AOI22X1 U4343 ( .IN1(N2873), .IN2(n3304), .IN3(N2433), .IN4(n3316), .QN(
        n4976) );
  OA22X1 U4344 ( .IN1(n3852), .IN2(n3327), .IN3(n3192), .IN4(n4759), .Q(n4975)
         );
  NAND4X0 U4345 ( .IN1(n4981), .IN2(n4982), .IN3(n4983), .IN4(n4984), .QN(
        n2508) );
  OA22X1 U4346 ( .IN1(n3260), .IN2(n4985), .IN3(n3268), .IN4(n4986), .Q(n4984)
         );
  AOI22X1 U4347 ( .IN1(N1497), .IN2(n3280), .IN3(n47), .IN4(n3292), .QN(n4983)
         );
  AOI22X1 U4348 ( .IN1(N2874), .IN2(n3304), .IN3(N2434), .IN4(n3316), .QN(
        n4982) );
  OA22X1 U4349 ( .IN1(n3851), .IN2(n3327), .IN3(n3192), .IN4(n4764), .Q(n4981)
         );
  NAND4X0 U4350 ( .IN1(n4987), .IN2(n4988), .IN3(n4989), .IN4(n4990), .QN(
        n2507) );
  OA22X1 U4351 ( .IN1(n3261), .IN2(n4991), .IN3(n3269), .IN4(n4992), .Q(n4990)
         );
  AOI22X1 U4352 ( .IN1(N1498), .IN2(n3281), .IN3(n46), .IN4(n3293), .QN(n4989)
         );
  AOI22X1 U4353 ( .IN1(N2875), .IN2(n3305), .IN3(N2435), .IN4(n3317), .QN(
        n4988) );
  OA22X1 U4354 ( .IN1(n3850), .IN2(n3326), .IN3(n3189), .IN4(n4769), .Q(n4987)
         );
  NAND4X0 U4355 ( .IN1(n4993), .IN2(n4994), .IN3(n4995), .IN4(n4996), .QN(
        n2506) );
  OA22X1 U4356 ( .IN1(n3261), .IN2(n4997), .IN3(n3269), .IN4(n4998), .Q(n4996)
         );
  AOI22X1 U4357 ( .IN1(N1499), .IN2(n3281), .IN3(n45), .IN4(n3293), .QN(n4995)
         );
  AOI22X1 U4358 ( .IN1(N2876), .IN2(n3305), .IN3(N2436), .IN4(n3317), .QN(
        n4994) );
  OA22X1 U4359 ( .IN1(n3849), .IN2(n3326), .IN3(n3192), .IN4(n2891), .Q(n4993)
         );
  NAND4X0 U4360 ( .IN1(n4999), .IN2(n5000), .IN3(n5001), .IN4(n5002), .QN(
        n2505) );
  OA22X1 U4361 ( .IN1(n3261), .IN2(n5003), .IN3(n3269), .IN4(n5004), .Q(n5002)
         );
  AOI22X1 U4362 ( .IN1(N1500), .IN2(n3281), .IN3(n44), .IN4(n3293), .QN(n5001)
         );
  AOI22X1 U4363 ( .IN1(N2877), .IN2(n3305), .IN3(N2437), .IN4(n3317), .QN(
        n5000) );
  OA22X1 U4364 ( .IN1(n3848), .IN2(n3326), .IN3(n3192), .IN4(n2892), .Q(n4999)
         );
  NAND4X0 U4365 ( .IN1(n5005), .IN2(n5006), .IN3(n5007), .IN4(n5008), .QN(
        n2504) );
  OA22X1 U4366 ( .IN1(n3261), .IN2(n5009), .IN3(n3269), .IN4(n5010), .Q(n5008)
         );
  AOI22X1 U4367 ( .IN1(N1501), .IN2(n3281), .IN3(n43), .IN4(n3293), .QN(n5007)
         );
  AOI22X1 U4368 ( .IN1(N2878), .IN2(n3305), .IN3(N2438), .IN4(n3317), .QN(
        n5006) );
  OA22X1 U4369 ( .IN1(n3847), .IN2(n3326), .IN3(n3192), .IN4(n2893), .Q(n5005)
         );
  NAND4X0 U4370 ( .IN1(n5011), .IN2(n5012), .IN3(n5013), .IN4(n5014), .QN(
        n2503) );
  OA22X1 U4371 ( .IN1(n3261), .IN2(n5015), .IN3(n3270), .IN4(n5016), .Q(n5014)
         );
  AOI22X1 U4372 ( .IN1(N1502), .IN2(n3282), .IN3(n42), .IN4(n3294), .QN(n5013)
         );
  AOI22X1 U4373 ( .IN1(N2879), .IN2(n3306), .IN3(N2439), .IN4(n3318), .QN(
        n5012) );
  OA22X1 U4374 ( .IN1(n3846), .IN2(n3325), .IN3(n3193), .IN4(n2894), .Q(n5011)
         );
  NAND4X0 U4375 ( .IN1(n5017), .IN2(n5018), .IN3(n5019), .IN4(n5020), .QN(
        n2502) );
  OA22X1 U4376 ( .IN1(n3262), .IN2(n5021), .IN3(n3270), .IN4(n5022), .Q(n5020)
         );
  AOI22X1 U4377 ( .IN1(N1503), .IN2(n3282), .IN3(n41), .IN4(n3294), .QN(n5019)
         );
  AOI22X1 U4378 ( .IN1(N2880), .IN2(n3306), .IN3(N2440), .IN4(n3318), .QN(
        n5018) );
  OA22X1 U4379 ( .IN1(n3845), .IN2(n3325), .IN3(n3193), .IN4(n2895), .Q(n5017)
         );
  NAND4X0 U4380 ( .IN1(n5023), .IN2(n5024), .IN3(n5025), .IN4(n5026), .QN(
        n2501) );
  OA22X1 U4381 ( .IN1(n3262), .IN2(n5027), .IN3(n3270), .IN4(n5028), .Q(n5026)
         );
  AOI22X1 U4382 ( .IN1(N1504), .IN2(n3282), .IN3(n40), .IN4(n3294), .QN(n5025)
         );
  AOI22X1 U4383 ( .IN1(N2881), .IN2(n3306), .IN3(N2441), .IN4(n3318), .QN(
        n5024) );
  OA22X1 U4384 ( .IN1(n3844), .IN2(n3325), .IN3(n3193), .IN4(n2896), .Q(n5023)
         );
  NAND4X0 U4385 ( .IN1(n5029), .IN2(n5030), .IN3(n5031), .IN4(n5032), .QN(
        n2500) );
  OA22X1 U4386 ( .IN1(n3262), .IN2(n5033), .IN3(n3270), .IN4(n5034), .Q(n5032)
         );
  AOI22X1 U4387 ( .IN1(N1505), .IN2(n3282), .IN3(n39), .IN4(n3294), .QN(n5031)
         );
  AOI22X1 U4388 ( .IN1(N2882), .IN2(n3306), .IN3(N2442), .IN4(n3318), .QN(
        n5030) );
  OA22X1 U4389 ( .IN1(n3843), .IN2(n3325), .IN3(n3193), .IN4(n2897), .Q(n5029)
         );
  NAND4X0 U4390 ( .IN1(n5035), .IN2(n5036), .IN3(n5037), .IN4(n5038), .QN(
        n2499) );
  OA22X1 U4391 ( .IN1(n3262), .IN2(n5039), .IN3(n3271), .IN4(n5040), .Q(n5038)
         );
  AOI22X1 U4392 ( .IN1(N1506), .IN2(n3283), .IN3(n38), .IN4(n3295), .QN(n5037)
         );
  AOI22X1 U4393 ( .IN1(N2883), .IN2(n3307), .IN3(N2443), .IN4(n3319), .QN(
        n5036) );
  OA22X1 U4394 ( .IN1(n3842), .IN2(n3324), .IN3(n3193), .IN4(n2898), .Q(n5035)
         );
  NAND4X0 U4395 ( .IN1(n5041), .IN2(n5042), .IN3(n5043), .IN4(n5044), .QN(
        n2498) );
  OA22X1 U4396 ( .IN1(n3262), .IN2(n5045), .IN3(n3271), .IN4(n5046), .Q(n5044)
         );
  AOI22X1 U4397 ( .IN1(N1507), .IN2(n3283), .IN3(n37), .IN4(n3295), .QN(n5043)
         );
  AOI22X1 U4398 ( .IN1(N2884), .IN2(n3307), .IN3(N2444), .IN4(n3319), .QN(
        n5042) );
  OA22X1 U4399 ( .IN1(n3841), .IN2(n3324), .IN3(n3194), .IN4(n2899), .Q(n5041)
         );
  NAND4X0 U4400 ( .IN1(n5047), .IN2(n5048), .IN3(n5049), .IN4(n5050), .QN(
        n2497) );
  OA22X1 U4401 ( .IN1(n3263), .IN2(n5051), .IN3(n3271), .IN4(n5052), .Q(n5050)
         );
  AOI22X1 U4402 ( .IN1(N1508), .IN2(n3283), .IN3(n36), .IN4(n3295), .QN(n5049)
         );
  AOI22X1 U4403 ( .IN1(N2885), .IN2(n3307), .IN3(N2445), .IN4(n3319), .QN(
        n5048) );
  OA22X1 U4404 ( .IN1(n3840), .IN2(n3324), .IN3(n3194), .IN4(n2900), .Q(n5047)
         );
  NAND4X0 U4405 ( .IN1(n5053), .IN2(n5054), .IN3(n5055), .IN4(n5056), .QN(
        n2496) );
  OA22X1 U4406 ( .IN1(n3263), .IN2(n5057), .IN3(n3271), .IN4(n5058), .Q(n5056)
         );
  NAND2X0 U4407 ( .IN1(n5059), .IN2(n5060), .QN(n4070) );
  NAND3X0 U4408 ( .IN1(n5060), .IN2(n4657), .IN3(N2392), .QN(n4068) );
  AOI22X1 U4409 ( .IN1(N1509), .IN2(n3283), .IN3(n35), .IN4(n3295), .QN(n5055)
         );
  ISOLANDX1 U4410 ( .D(n5060), .ISO(n5061), .Q(n4073) );
  ISOLANDX1 U4411 ( .D(n5060), .ISO(n5062), .Q(n4072) );
  AOI22X1 U4412 ( .IN1(N2886), .IN2(n3307), .IN3(N2446), .IN4(n3319), .QN(
        n5054) );
  ISOLANDX1 U4413 ( .D(n5060), .ISO(n5063), .Q(n4075) );
  ISOLANDX1 U4414 ( .D(n5060), .ISO(n5064), .Q(n4074) );
  OA22X1 U4415 ( .IN1(n3868), .IN2(n3328), .IN3(n3194), .IN4(n2901), .Q(n5053)
         );
  NAND2X0 U4416 ( .IN1(n5065), .IN2(n4146), .QN(n4076) );
  NAND2X0 U4417 ( .IN1(n4017), .IN2(n5066), .QN(n4146) );
  NAND3X0 U4418 ( .IN1(n5067), .IN2(n5068), .IN3(n5069), .QN(n2495) );
  AOI222X1 U4419 ( .IN1(N997), .IN2(n3383), .IN3(rEIP_0_), .IN4(n3196), .IN5(
        N964), .IN6(n3391), .QN(n5069) );
  OA22X1 U4420 ( .IN1(n5070), .IN2(n3478), .IN3(n4877), .IN4(n3490), .Q(n5068)
         );
  INVX0 U4421 ( .IN(N2995), .QN(n4877) );
  INVX0 U4422 ( .IN(N2856), .QN(n5070) );
  OA22X1 U4423 ( .IN1(n4878), .IN2(n3502), .IN3(n1589), .IN4(n3514), .Q(n5067)
         );
  INVX0 U4424 ( .IN(N3067), .QN(n4878) );
  NAND3X0 U4425 ( .IN1(n5075), .IN2(n5076), .IN3(n5077), .QN(n2494) );
  AOI222X1 U4426 ( .IN1(N998), .IN2(n3383), .IN3(rEIP_1_), .IN4(n3201), .IN5(
        N965), .IN6(n3390), .QN(n5077) );
  OA22X1 U4427 ( .IN1(n5078), .IN2(n3478), .IN3(n4883), .IN4(n3490), .Q(n5076)
         );
  INVX0 U4428 ( .IN(N2996), .QN(n4883) );
  INVX0 U4429 ( .IN(N2857), .QN(n5078) );
  OA22X1 U4430 ( .IN1(n4884), .IN2(n3502), .IN3(n1588), .IN4(n3520), .Q(n5075)
         );
  INVX0 U4431 ( .IN(N3068), .QN(n4884) );
  NAND3X0 U4432 ( .IN1(n5079), .IN2(n5080), .IN3(n5081), .QN(n2493) );
  AOI222X1 U4433 ( .IN1(N999), .IN2(n3382), .IN3(rEIP_2_), .IN4(n3201), .IN5(
        N966), .IN6(n3390), .QN(n5081) );
  OA22X1 U4434 ( .IN1(n5082), .IN2(n3478), .IN3(n4889), .IN4(n3490), .Q(n5080)
         );
  INVX0 U4435 ( .IN(N2997), .QN(n4889) );
  INVX0 U4436 ( .IN(N2858), .QN(n5082) );
  OA22X1 U4437 ( .IN1(n4890), .IN2(n3502), .IN3(n1587), .IN4(n3520), .Q(n5079)
         );
  INVX0 U4438 ( .IN(N3069), .QN(n4890) );
  NAND3X0 U4439 ( .IN1(n5083), .IN2(n5084), .IN3(n5085), .QN(n2492) );
  AOI222X1 U4440 ( .IN1(N1000), .IN2(n3382), .IN3(rEIP_3_), .IN4(n3200), .IN5(
        N967), .IN6(n3390), .QN(n5085) );
  OA22X1 U4441 ( .IN1(n5086), .IN2(n3478), .IN3(n4895), .IN4(n3490), .Q(n5084)
         );
  INVX0 U4442 ( .IN(N2998), .QN(n4895) );
  INVX0 U4443 ( .IN(N2859), .QN(n5086) );
  OA22X1 U4444 ( .IN1(n4896), .IN2(n3502), .IN3(n1586), .IN4(n3520), .Q(n5083)
         );
  INVX0 U4445 ( .IN(N3070), .QN(n4896) );
  NAND3X0 U4446 ( .IN1(n5087), .IN2(n5088), .IN3(n5089), .QN(n2491) );
  AOI222X1 U4447 ( .IN1(N1001), .IN2(n3382), .IN3(rEIP_4_), .IN4(n3200), .IN5(
        N968), .IN6(n3391), .QN(n5089) );
  OA22X1 U4448 ( .IN1(n5090), .IN2(n3479), .IN3(n4901), .IN4(n3491), .Q(n5088)
         );
  INVX0 U4449 ( .IN(N2999), .QN(n4901) );
  INVX0 U4450 ( .IN(N2860), .QN(n5090) );
  OA22X1 U4451 ( .IN1(n4902), .IN2(n3503), .IN3(n1585), .IN4(n3520), .Q(n5087)
         );
  INVX0 U4452 ( .IN(N3071), .QN(n4902) );
  NAND3X0 U4453 ( .IN1(n5091), .IN2(n5092), .IN3(n5093), .QN(n2490) );
  AOI222X1 U4454 ( .IN1(N1002), .IN2(n3382), .IN3(rEIP_5_), .IN4(n3200), .IN5(
        N969), .IN6(n3391), .QN(n5093) );
  OA22X1 U4455 ( .IN1(n5094), .IN2(n3479), .IN3(n4907), .IN4(n3491), .Q(n5092)
         );
  INVX0 U4456 ( .IN(N3000), .QN(n4907) );
  INVX0 U4457 ( .IN(N2861), .QN(n5094) );
  OA22X1 U4458 ( .IN1(n4908), .IN2(n3503), .IN3(n1584), .IN4(n3520), .Q(n5091)
         );
  INVX0 U4459 ( .IN(N3072), .QN(n4908) );
  NAND3X0 U4460 ( .IN1(n5095), .IN2(n5096), .IN3(n5097), .QN(n2489) );
  AOI222X1 U4461 ( .IN1(N1003), .IN2(n3382), .IN3(test_so18), .IN4(n3203), 
        .IN5(N970), .IN6(n3390), .QN(n5097) );
  OA22X1 U4462 ( .IN1(n5098), .IN2(n3479), .IN3(n4913), .IN4(n3491), .Q(n5096)
         );
  INVX0 U4463 ( .IN(N3001), .QN(n4913) );
  INVX0 U4464 ( .IN(N2862), .QN(n5098) );
  OA22X1 U4465 ( .IN1(n4914), .IN2(n3503), .IN3(n1583), .IN4(n3519), .Q(n5095)
         );
  INVX0 U4466 ( .IN(N3073), .QN(n4914) );
  NAND3X0 U4467 ( .IN1(n5099), .IN2(n5100), .IN3(n5101), .QN(n2488) );
  AOI222X1 U4468 ( .IN1(N1004), .IN2(n3381), .IN3(rEIP_7_), .IN4(n3202), .IN5(
        N971), .IN6(n3390), .QN(n5101) );
  OA22X1 U4469 ( .IN1(n5102), .IN2(n3479), .IN3(n4919), .IN4(n3491), .Q(n5100)
         );
  INVX0 U4470 ( .IN(N3002), .QN(n4919) );
  INVX0 U4471 ( .IN(N2863), .QN(n5102) );
  OA22X1 U4472 ( .IN1(n4920), .IN2(n3503), .IN3(n1582), .IN4(n3519), .Q(n5099)
         );
  INVX0 U4473 ( .IN(N3074), .QN(n4920) );
  NAND3X0 U4474 ( .IN1(n5103), .IN2(n5104), .IN3(n5105), .QN(n2487) );
  AOI222X1 U4475 ( .IN1(N1005), .IN2(n3381), .IN3(rEIP_8_), .IN4(n3202), .IN5(
        N972), .IN6(n3390), .QN(n5105) );
  OA22X1 U4476 ( .IN1(n5106), .IN2(n3480), .IN3(n4925), .IN4(n3492), .Q(n5104)
         );
  INVX0 U4477 ( .IN(N3003), .QN(n4925) );
  INVX0 U4478 ( .IN(N2864), .QN(n5106) );
  OA22X1 U4479 ( .IN1(n4926), .IN2(n3504), .IN3(n1581), .IN4(n3519), .Q(n5103)
         );
  INVX0 U4480 ( .IN(N3075), .QN(n4926) );
  NAND3X0 U4481 ( .IN1(n5107), .IN2(n5108), .IN3(n5109), .QN(n2486) );
  AOI222X1 U4482 ( .IN1(N1006), .IN2(n3381), .IN3(rEIP_9_), .IN4(n3202), .IN5(
        N973), .IN6(n3390), .QN(n5109) );
  OA22X1 U4483 ( .IN1(n5110), .IN2(n3480), .IN3(n4931), .IN4(n3492), .Q(n5108)
         );
  INVX0 U4484 ( .IN(N3004), .QN(n4931) );
  INVX0 U4485 ( .IN(N2865), .QN(n5110) );
  OA22X1 U4486 ( .IN1(n4932), .IN2(n3504), .IN3(n1580), .IN4(n3519), .Q(n5107)
         );
  INVX0 U4487 ( .IN(N3076), .QN(n4932) );
  NAND3X0 U4488 ( .IN1(n5111), .IN2(n5112), .IN3(n5113), .QN(n2485) );
  AOI222X1 U4489 ( .IN1(N1007), .IN2(n3381), .IN3(rEIP_10_), .IN4(n3201), 
        .IN5(N974), .IN6(n3391), .QN(n5113) );
  OA22X1 U4490 ( .IN1(n5114), .IN2(n3480), .IN3(n4937), .IN4(n3492), .Q(n5112)
         );
  INVX0 U4491 ( .IN(N3005), .QN(n4937) );
  INVX0 U4492 ( .IN(N2866), .QN(n5114) );
  OA22X1 U4493 ( .IN1(n4938), .IN2(n3504), .IN3(n1579), .IN4(n3519), .Q(n5111)
         );
  INVX0 U4494 ( .IN(N3077), .QN(n4938) );
  NAND3X0 U4495 ( .IN1(n5115), .IN2(n5116), .IN3(n5117), .QN(n2484) );
  AOI222X1 U4496 ( .IN1(N1008), .IN2(n3381), .IN3(rEIP_11_), .IN4(n3199), 
        .IN5(N975), .IN6(n3390), .QN(n5117) );
  OA22X1 U4497 ( .IN1(n5118), .IN2(n3480), .IN3(n4943), .IN4(n3492), .Q(n5116)
         );
  INVX0 U4498 ( .IN(N3006), .QN(n4943) );
  INVX0 U4499 ( .IN(N2867), .QN(n5118) );
  OA22X1 U4500 ( .IN1(n4944), .IN2(n3504), .IN3(n1578), .IN4(n3518), .Q(n5115)
         );
  INVX0 U4501 ( .IN(N3078), .QN(n4944) );
  NAND3X0 U4502 ( .IN1(n5119), .IN2(n5120), .IN3(n5121), .QN(n2483) );
  AOI222X1 U4503 ( .IN1(N1009), .IN2(n3380), .IN3(rEIP_12_), .IN4(n3198), 
        .IN5(N976), .IN6(n3391), .QN(n5121) );
  OA22X1 U4504 ( .IN1(n5122), .IN2(n3481), .IN3(n4949), .IN4(n3493), .Q(n5120)
         );
  INVX0 U4505 ( .IN(N3007), .QN(n4949) );
  INVX0 U4506 ( .IN(N2868), .QN(n5122) );
  OA22X1 U4507 ( .IN1(n4950), .IN2(n3505), .IN3(n1577), .IN4(n3518), .Q(n5119)
         );
  INVX0 U4508 ( .IN(N3079), .QN(n4950) );
  NAND3X0 U4509 ( .IN1(n5123), .IN2(n5124), .IN3(n5125), .QN(n2482) );
  AOI222X1 U4510 ( .IN1(N1010), .IN2(n3380), .IN3(rEIP_13_), .IN4(n3198), 
        .IN5(N977), .IN6(n3390), .QN(n5125) );
  OA22X1 U4511 ( .IN1(n5126), .IN2(n3481), .IN3(n4955), .IN4(n3493), .Q(n5124)
         );
  INVX0 U4512 ( .IN(N3008), .QN(n4955) );
  INVX0 U4513 ( .IN(N2869), .QN(n5126) );
  OA22X1 U4514 ( .IN1(n4956), .IN2(n3505), .IN3(n1576), .IN4(n3518), .Q(n5123)
         );
  INVX0 U4515 ( .IN(N3080), .QN(n4956) );
  NAND3X0 U4516 ( .IN1(n5127), .IN2(n5128), .IN3(n5129), .QN(n2481) );
  AOI222X1 U4517 ( .IN1(N1011), .IN2(n3380), .IN3(rEIP_14_), .IN4(n3198), 
        .IN5(N978), .IN6(n3390), .QN(n5129) );
  OA22X1 U4518 ( .IN1(n5130), .IN2(n3481), .IN3(n4961), .IN4(n3493), .Q(n5128)
         );
  INVX0 U4519 ( .IN(N3009), .QN(n4961) );
  INVX0 U4520 ( .IN(N2870), .QN(n5130) );
  OA22X1 U4521 ( .IN1(n4962), .IN2(n3505), .IN3(n1575), .IN4(n3518), .Q(n5127)
         );
  INVX0 U4522 ( .IN(N3081), .QN(n4962) );
  NAND3X0 U4523 ( .IN1(n5131), .IN2(n5132), .IN3(n5133), .QN(n2480) );
  AOI222X1 U4524 ( .IN1(N1012), .IN2(n3380), .IN3(rEIP_15_), .IN4(n3197), 
        .IN5(N979), .IN6(n3390), .QN(n5133) );
  OA22X1 U4525 ( .IN1(n5134), .IN2(n3481), .IN3(n4967), .IN4(n3493), .Q(n5132)
         );
  INVX0 U4526 ( .IN(N3010), .QN(n4967) );
  INVX0 U4527 ( .IN(N2871), .QN(n5134) );
  OA22X1 U4528 ( .IN1(n4968), .IN2(n3505), .IN3(n1574), .IN4(n3518), .Q(n5131)
         );
  INVX0 U4529 ( .IN(N3082), .QN(n4968) );
  NAND3X0 U4530 ( .IN1(n5135), .IN2(n5136), .IN3(n5137), .QN(n2479) );
  AOI222X1 U4531 ( .IN1(N1013), .IN2(n3380), .IN3(rEIP_16_), .IN4(n3200), 
        .IN5(N980), .IN6(n3390), .QN(n5137) );
  OA22X1 U4532 ( .IN1(n5138), .IN2(n3482), .IN3(n4973), .IN4(n3494), .Q(n5136)
         );
  INVX0 U4533 ( .IN(N3011), .QN(n4973) );
  INVX0 U4534 ( .IN(N2872), .QN(n5138) );
  OA22X1 U4535 ( .IN1(n4974), .IN2(n3506), .IN3(n1573), .IN4(n3517), .Q(n5135)
         );
  INVX0 U4536 ( .IN(N3083), .QN(n4974) );
  NAND3X0 U4537 ( .IN1(n5139), .IN2(n5140), .IN3(n5141), .QN(n2478) );
  AOI222X1 U4538 ( .IN1(N1014), .IN2(n3379), .IN3(rEIP_17_), .IN4(n3202), 
        .IN5(N981), .IN6(n3390), .QN(n5141) );
  OA22X1 U4539 ( .IN1(n5142), .IN2(n3482), .IN3(n4979), .IN4(n3494), .Q(n5140)
         );
  INVX0 U4540 ( .IN(N3012), .QN(n4979) );
  INVX0 U4541 ( .IN(N2873), .QN(n5142) );
  OA22X1 U4542 ( .IN1(n4980), .IN2(n3506), .IN3(n1572), .IN4(n3517), .Q(n5139)
         );
  INVX0 U4543 ( .IN(N3084), .QN(n4980) );
  NAND3X0 U4544 ( .IN1(n5143), .IN2(n5144), .IN3(n5145), .QN(n2477) );
  AOI222X1 U4545 ( .IN1(N1015), .IN2(n3379), .IN3(rEIP_18_), .IN4(n3199), 
        .IN5(N982), .IN6(n3391), .QN(n5145) );
  OA22X1 U4546 ( .IN1(n5146), .IN2(n3482), .IN3(n4985), .IN4(n3494), .Q(n5144)
         );
  INVX0 U4547 ( .IN(N3013), .QN(n4985) );
  INVX0 U4548 ( .IN(N2874), .QN(n5146) );
  OA22X1 U4549 ( .IN1(n4986), .IN2(n3506), .IN3(n1571), .IN4(n3517), .Q(n5143)
         );
  INVX0 U4550 ( .IN(N3085), .QN(n4986) );
  NAND3X0 U4551 ( .IN1(n5147), .IN2(n5148), .IN3(n5149), .QN(n2476) );
  AOI222X1 U4552 ( .IN1(N1016), .IN2(n3379), .IN3(rEIP_19_), .IN4(n3199), 
        .IN5(N983), .IN6(n3391), .QN(n5149) );
  OA22X1 U4553 ( .IN1(n5150), .IN2(n3482), .IN3(n4991), .IN4(n3494), .Q(n5148)
         );
  INVX0 U4554 ( .IN(N3014), .QN(n4991) );
  INVX0 U4555 ( .IN(N2875), .QN(n5150) );
  OA22X1 U4556 ( .IN1(n4992), .IN2(n3506), .IN3(n1570), .IN4(n3517), .Q(n5147)
         );
  INVX0 U4557 ( .IN(N3086), .QN(n4992) );
  NAND3X0 U4558 ( .IN1(n5151), .IN2(n5152), .IN3(n5153), .QN(n2475) );
  AOI222X1 U4559 ( .IN1(N1017), .IN2(n3379), .IN3(rEIP_20_), .IN4(n3200), 
        .IN5(N984), .IN6(n3391), .QN(n5153) );
  OA22X1 U4560 ( .IN1(n5154), .IN2(n3483), .IN3(n4997), .IN4(n3495), .Q(n5152)
         );
  INVX0 U4561 ( .IN(N3015), .QN(n4997) );
  INVX0 U4562 ( .IN(N2876), .QN(n5154) );
  OA22X1 U4563 ( .IN1(n4998), .IN2(n3507), .IN3(n1569), .IN4(n3516), .Q(n5151)
         );
  INVX0 U4564 ( .IN(N3087), .QN(n4998) );
  NAND3X0 U4565 ( .IN1(n5155), .IN2(n5156), .IN3(n5157), .QN(n2474) );
  AOI222X1 U4566 ( .IN1(N1018), .IN2(n3379), .IN3(rEIP_21_), .IN4(n3202), 
        .IN5(N985), .IN6(n3391), .QN(n5157) );
  OA22X1 U4567 ( .IN1(n5158), .IN2(n3483), .IN3(n5003), .IN4(n3495), .Q(n5156)
         );
  INVX0 U4568 ( .IN(N3016), .QN(n5003) );
  INVX0 U4569 ( .IN(N2877), .QN(n5158) );
  OA22X1 U4570 ( .IN1(n5004), .IN2(n3507), .IN3(n1568), .IN4(n3516), .Q(n5155)
         );
  INVX0 U4571 ( .IN(N3088), .QN(n5004) );
  NAND3X0 U4572 ( .IN1(n5159), .IN2(n5160), .IN3(n5161), .QN(n2473) );
  AOI222X1 U4573 ( .IN1(N1019), .IN2(n3378), .IN3(rEIP_22_), .IN4(n3201), 
        .IN5(N986), .IN6(n3391), .QN(n5161) );
  OA22X1 U4574 ( .IN1(n5162), .IN2(n3483), .IN3(n5009), .IN4(n3495), .Q(n5160)
         );
  INVX0 U4575 ( .IN(N3017), .QN(n5009) );
  INVX0 U4576 ( .IN(N2878), .QN(n5162) );
  OA22X1 U4577 ( .IN1(n5010), .IN2(n3507), .IN3(n1567), .IN4(n3516), .Q(n5159)
         );
  INVX0 U4578 ( .IN(N3089), .QN(n5010) );
  NAND3X0 U4579 ( .IN1(n5163), .IN2(n5164), .IN3(n5165), .QN(n2472) );
  AOI222X1 U4580 ( .IN1(N1020), .IN2(n3378), .IN3(rEIP_23_), .IN4(n3201), 
        .IN5(N987), .IN6(n3391), .QN(n5165) );
  OA22X1 U4581 ( .IN1(n5166), .IN2(n3483), .IN3(n5015), .IN4(n3495), .Q(n5164)
         );
  INVX0 U4582 ( .IN(N3018), .QN(n5015) );
  INVX0 U4583 ( .IN(N2879), .QN(n5166) );
  OA22X1 U4584 ( .IN1(n5016), .IN2(n3507), .IN3(n1566), .IN4(n3516), .Q(n5163)
         );
  INVX0 U4585 ( .IN(N3090), .QN(n5016) );
  NAND3X0 U4586 ( .IN1(n5167), .IN2(n5168), .IN3(n5169), .QN(n2471) );
  AOI222X1 U4587 ( .IN1(N1021), .IN2(n3378), .IN3(rEIP_24_), .IN4(n3196), 
        .IN5(N988), .IN6(n3390), .QN(n5169) );
  OA22X1 U4588 ( .IN1(n5170), .IN2(n3484), .IN3(n5021), .IN4(n3496), .Q(n5168)
         );
  INVX0 U4589 ( .IN(N3019), .QN(n5021) );
  INVX0 U4590 ( .IN(N2880), .QN(n5170) );
  OA22X1 U4591 ( .IN1(n5022), .IN2(n3508), .IN3(n1565), .IN4(n3516), .Q(n5167)
         );
  INVX0 U4592 ( .IN(N3091), .QN(n5022) );
  NAND3X0 U4593 ( .IN1(n5171), .IN2(n5172), .IN3(n5173), .QN(n2470) );
  AOI222X1 U4594 ( .IN1(N1022), .IN2(n3378), .IN3(rEIP_25_), .IN4(n3196), 
        .IN5(N989), .IN6(n3390), .QN(n5173) );
  OA22X1 U4595 ( .IN1(n5174), .IN2(n3484), .IN3(n5027), .IN4(n3496), .Q(n5172)
         );
  INVX0 U4596 ( .IN(N3020), .QN(n5027) );
  INVX0 U4597 ( .IN(N2881), .QN(n5174) );
  OA22X1 U4598 ( .IN1(n5028), .IN2(n3508), .IN3(n1564), .IN4(n3515), .Q(n5171)
         );
  INVX0 U4599 ( .IN(N3092), .QN(n5028) );
  NAND3X0 U4600 ( .IN1(n5175), .IN2(n5176), .IN3(n5177), .QN(n2469) );
  AOI222X1 U4601 ( .IN1(N1023), .IN2(n3378), .IN3(test_so19), .IN4(n3197), 
        .IN5(N990), .IN6(n3391), .QN(n5177) );
  OA22X1 U4602 ( .IN1(n5178), .IN2(n3484), .IN3(n5033), .IN4(n3496), .Q(n5176)
         );
  INVX0 U4603 ( .IN(N3021), .QN(n5033) );
  INVX0 U4604 ( .IN(N2882), .QN(n5178) );
  OA22X1 U4605 ( .IN1(n5034), .IN2(n3508), .IN3(n1563), .IN4(n3517), .Q(n5175)
         );
  INVX0 U4606 ( .IN(N3093), .QN(n5034) );
  NAND3X0 U4607 ( .IN1(n5179), .IN2(n5180), .IN3(n5181), .QN(n2468) );
  AOI222X1 U4608 ( .IN1(N1024), .IN2(n3377), .IN3(rEIP_27_), .IN4(n3197), 
        .IN5(N991), .IN6(n3390), .QN(n5181) );
  OA22X1 U4609 ( .IN1(n5182), .IN2(n3484), .IN3(n5039), .IN4(n3496), .Q(n5180)
         );
  INVX0 U4610 ( .IN(N3022), .QN(n5039) );
  INVX0 U4611 ( .IN(N2883), .QN(n5182) );
  OA22X1 U4612 ( .IN1(n5040), .IN2(n3508), .IN3(n1562), .IN4(n3515), .Q(n5179)
         );
  INVX0 U4613 ( .IN(N3094), .QN(n5040) );
  NAND3X0 U4614 ( .IN1(n5183), .IN2(n5184), .IN3(n5185), .QN(n2467) );
  AOI222X1 U4615 ( .IN1(N1025), .IN2(n3377), .IN3(rEIP_28_), .IN4(n3197), 
        .IN5(N992), .IN6(n3392), .QN(n5185) );
  OA22X1 U4616 ( .IN1(n5186), .IN2(n3485), .IN3(n5045), .IN4(n3497), .Q(n5184)
         );
  INVX0 U4617 ( .IN(N3023), .QN(n5045) );
  INVX0 U4618 ( .IN(N2884), .QN(n5186) );
  OA22X1 U4619 ( .IN1(n5046), .IN2(n3509), .IN3(n1561), .IN4(n3515), .Q(n5183)
         );
  INVX0 U4620 ( .IN(N3095), .QN(n5046) );
  NAND3X0 U4621 ( .IN1(n5187), .IN2(n5188), .IN3(n5189), .QN(n2466) );
  AOI222X1 U4622 ( .IN1(N1026), .IN2(n3377), .IN3(rEIP_29_), .IN4(n3198), 
        .IN5(N993), .IN6(n3392), .QN(n5189) );
  OA22X1 U4623 ( .IN1(n5190), .IN2(n3485), .IN3(n5051), .IN4(n3497), .Q(n5188)
         );
  INVX0 U4624 ( .IN(N3024), .QN(n5051) );
  INVX0 U4625 ( .IN(N2885), .QN(n5190) );
  OA22X1 U4626 ( .IN1(n5052), .IN2(n3509), .IN3(n1560), .IN4(n3515), .Q(n5187)
         );
  INVX0 U4627 ( .IN(N3096), .QN(n5052) );
  NAND3X0 U4628 ( .IN1(n5191), .IN2(n5192), .IN3(n5193), .QN(n2465) );
  AOI222X1 U4629 ( .IN1(N1027), .IN2(n3377), .IN3(rEIP_30_), .IN4(n3199), 
        .IN5(N994), .IN6(n3392), .QN(n5193) );
  OA22X1 U4630 ( .IN1(n5194), .IN2(n3485), .IN3(n5057), .IN4(n3497), .Q(n5192)
         );
  INVX0 U4631 ( .IN(N3025), .QN(n5057) );
  INVX0 U4632 ( .IN(N2886), .QN(n5194) );
  OA22X1 U4633 ( .IN1(n5058), .IN2(n3509), .IN3(n1559), .IN4(n3515), .Q(n5191)
         );
  INVX0 U4634 ( .IN(N3097), .QN(n5058) );
  NAND3X0 U4635 ( .IN1(n5195), .IN2(n5196), .IN3(n5197), .QN(n2464) );
  AOI222X1 U4636 ( .IN1(N1029), .IN2(n3377), .IN3(n3195), .IN4(rEIP_31_), 
        .IN5(N995), .IN6(n3391), .QN(n5197) );
  NOR2X0 U4637 ( .IN1(n4174), .IN2(n1472), .QN(n4164) );
  NAND2X0 U4638 ( .IN1(n4090), .IN2(n4113), .QN(n4156) );
  INVX0 U4639 ( .IN(n4163), .QN(n4113) );
  NOR2X0 U4640 ( .IN1(n4174), .IN2(n2868), .QN(n4163) );
  OA22X1 U4641 ( .IN1(n5198), .IN2(n3485), .IN3(n4069), .IN4(n3497), .Q(n5196)
         );
  NAND4X0 U4642 ( .IN1(N2392), .IN2(n4657), .IN3(n4017), .IN4(n3514), .QN(
        n5072) );
  INVX0 U4643 ( .IN(n5199), .QN(n4657) );
  INVX0 U4644 ( .IN(N3026), .QN(n4069) );
  NAND3X0 U4645 ( .IN1(n4017), .IN2(n3514), .IN3(n4655), .QN(n5071) );
  INVX0 U4646 ( .IN(n5064), .QN(n4655) );
  INVX0 U4647 ( .IN(N2887), .QN(n5198) );
  OA22X1 U4648 ( .IN1(n4071), .IN2(n3509), .IN3(n1558), .IN4(n3514), .Q(n5195)
         );
  NAND3X0 U4649 ( .IN1(n4017), .IN2(n3514), .IN3(n5059), .QN(n5073) );
  NOR2X0 U4650 ( .IN1(n5199), .IN2(N2392), .QN(n5059) );
  NAND2X0 U4651 ( .IN1(n5065), .IN2(n4103), .QN(n5074) );
  NOR2X0 U4652 ( .IN1(n4161), .IN2(n4254), .QN(n4103) );
  INVX0 U4653 ( .IN(n4090), .QN(n4161) );
  NAND3X0 U4654 ( .IN1(n5200), .IN2(n2865), .IN3(n1491), .QN(n4090) );
  OA21X1 U4655 ( .IN1(n4091), .IN2(n4106), .IN3(n3194), .Q(n5065) );
  NAND2X0 U4656 ( .IN1(n4649), .IN2(n5200), .QN(n4015) );
  NOR2X0 U4657 ( .IN1(n2844), .IN2(n2865), .QN(n4649) );
  OA22X1 U4658 ( .IN1(n5064), .IN2(n4123), .IN3(n4663), .IN4(n5199), .Q(n4106)
         );
  AO21X1 U4659 ( .IN1(n5201), .IN2(n5202), .IN3(n2955), .Q(n4663) );
  NAND2X0 U4660 ( .IN1(r680_B_1_), .IN2(gte_355_B_0_), .QN(n5202) );
  INVX0 U4661 ( .IN(n4868), .QN(n4123) );
  INVX0 U4662 ( .IN(N3098), .QN(n4071) );
  AO222X1 U4663 ( .IN1(n3531), .IN2(Datao[0]), .IN3(N3346), .IN4(n3532), .IN5(
        N3434), .IN6(n3344), .Q(n2463) );
  AO222X1 U4664 ( .IN1(n3531), .IN2(Datao[1]), .IN3(N3347), .IN4(n3532), .IN5(
        N3435), .IN6(n3344), .Q(n2462) );
  AO222X1 U4665 ( .IN1(n3530), .IN2(Datao[2]), .IN3(N3348), .IN4(n3532), .IN5(
        test_so17), .IN6(n3344), .Q(n2461) );
  AO222X1 U4666 ( .IN1(n3530), .IN2(Datao[3]), .IN3(N3349), .IN4(n3532), .IN5(
        N3437), .IN6(n3343), .Q(n2460) );
  AO222X1 U4667 ( .IN1(n3530), .IN2(Datao[4]), .IN3(N3350), .IN4(n3532), .IN5(
        N3438), .IN6(n3343), .Q(n2459) );
  AO222X1 U4668 ( .IN1(n3530), .IN2(Datao[5]), .IN3(N3351), .IN4(n3533), .IN5(
        N3439), .IN6(n3343), .Q(n2458) );
  AO222X1 U4669 ( .IN1(n3530), .IN2(Datao[6]), .IN3(N3352), .IN4(n3533), .IN5(
        N3440), .IN6(n3343), .Q(n2457) );
  AO222X1 U4670 ( .IN1(n3529), .IN2(Datao[7]), .IN3(N3353), .IN4(n3533), .IN5(
        N3441), .IN6(n3342), .Q(n2456) );
  AO222X1 U4671 ( .IN1(n3529), .IN2(Datao[8]), .IN3(N3354), .IN4(n3533), .IN5(
        N3442), .IN6(n3342), .Q(n2455) );
  AO222X1 U4672 ( .IN1(n3529), .IN2(Datao[9]), .IN3(test_so4), .IN4(n3533), 
        .IN5(N3443), .IN6(n3342), .Q(n2454) );
  AO222X1 U4673 ( .IN1(n3529), .IN2(Datao[10]), .IN3(N3356), .IN4(n3534), 
        .IN5(N3444), .IN6(n3342), .Q(n2453) );
  AO222X1 U4674 ( .IN1(n3529), .IN2(Datao[11]), .IN3(N3357), .IN4(n3534), 
        .IN5(N3445), .IN6(n3341), .Q(n2452) );
  AO222X1 U4675 ( .IN1(n3528), .IN2(Datao[12]), .IN3(N3358), .IN4(n3534), 
        .IN5(N3446), .IN6(n3341), .Q(n2451) );
  AO222X1 U4676 ( .IN1(n3528), .IN2(Datao[13]), .IN3(N3359), .IN4(n3534), 
        .IN5(N3447), .IN6(n3341), .Q(n2450) );
  AO222X1 U4677 ( .IN1(n3528), .IN2(Datao[14]), .IN3(N3360), .IN4(n3534), 
        .IN5(N3448), .IN6(n3341), .Q(n2449) );
  AO222X1 U4678 ( .IN1(n3528), .IN2(Datao[15]), .IN3(N3361), .IN4(n3535), 
        .IN5(N3449), .IN6(n3340), .Q(n2448) );
  AO222X1 U4679 ( .IN1(n3528), .IN2(Datao[16]), .IN3(n2970), .IN4(n3535), 
        .IN5(N3450), .IN6(n3340), .Q(n2447) );
  AO222X1 U4680 ( .IN1(n3527), .IN2(Datao[17]), .IN3(n2969), .IN4(n3535), 
        .IN5(N3451), .IN6(n3340), .Q(n2446) );
  AO222X1 U4681 ( .IN1(n3527), .IN2(Datao[18]), .IN3(n2968), .IN4(n3535), 
        .IN5(N3452), .IN6(n3340), .Q(n2445) );
  AO222X1 U4682 ( .IN1(n3527), .IN2(Datao[19]), .IN3(n2967), .IN4(n3535), 
        .IN5(N3453), .IN6(n3339), .Q(n2444) );
  AO222X1 U4683 ( .IN1(n3527), .IN2(Datao[20]), .IN3(n2966), .IN4(n3536), 
        .IN5(N3454), .IN6(n3339), .Q(n2443) );
  AO222X1 U4684 ( .IN1(n3527), .IN2(Datao[21]), .IN3(n2965), .IN4(n3536), 
        .IN5(N3455), .IN6(n3339), .Q(n2442) );
  AO222X1 U4685 ( .IN1(n3526), .IN2(Datao[22]), .IN3(n2964), .IN4(n3536), 
        .IN5(N3456), .IN6(n3339), .Q(n2441) );
  AO222X1 U4686 ( .IN1(n3526), .IN2(Datao[23]), .IN3(n2963), .IN4(n3536), 
        .IN5(N3457), .IN6(n3338), .Q(n2440) );
  AO222X1 U4687 ( .IN1(n3526), .IN2(Datao[24]), .IN3(n2962), .IN4(n3536), 
        .IN5(N3458), .IN6(n3338), .Q(n2439) );
  AO222X1 U4688 ( .IN1(n3526), .IN2(Datao[25]), .IN3(n2961), .IN4(n3537), 
        .IN5(N3459), .IN6(n3338), .Q(n2438) );
  AO222X1 U4689 ( .IN1(n3526), .IN2(Datao[26]), .IN3(n2960), .IN4(n3537), 
        .IN5(N3460), .IN6(n3338), .Q(n2437) );
  AO222X1 U4690 ( .IN1(n3525), .IN2(Datao[27]), .IN3(n2959), .IN4(n3537), 
        .IN5(N3461), .IN6(n3337), .Q(n2436) );
  AO222X1 U4691 ( .IN1(n3525), .IN2(Datao[28]), .IN3(n2958), .IN4(n3537), 
        .IN5(N3462), .IN6(n3337), .Q(n2435) );
  AO222X1 U4692 ( .IN1(n3525), .IN2(Datao[29]), .IN3(n2957), .IN4(n3537), 
        .IN5(N3463), .IN6(n3337), .Q(n2434) );
  AO222X1 U4693 ( .IN1(n3525), .IN2(Datao[30]), .IN3(n2846), .IN4(n3538), 
        .IN5(test_so20), .IN6(n3337), .Q(n2433) );
  INVX0 U4694 ( .IN(n4013), .QN(n4111) );
  NOR2X0 U4695 ( .IN1(n4091), .IN2(n3525), .QN(n5204) );
  AND2X1 U4696 ( .IN1(n4013), .IN2(n5205), .Q(n5203) );
  NAND4X0 U4697 ( .IN1(n4651), .IN2(n4017), .IN3(n5206), .IN4(n4019), .QN(
        n5205) );
  NOR2X0 U4698 ( .IN1(n4097), .IN2(n1492), .QN(n4116) );
  NAND3X0 U4699 ( .IN1(n2865), .IN2(n2844), .IN3(n5200), .QN(n4013) );
  NOR2X0 U4700 ( .IN1(n4097), .IN2(n2842), .QN(n5200) );
  OAI221X1 U4701 ( .IN1(n2864), .IN2(rEIP_1_), .IN3(n5207), .IN4(n3693), .IN5(
        n5208), .QN(n2432) );
  MUX21X1 U4702 ( .IN1(n5209), .IN2(BE_n[3]), .S(n3205), .Q(n2431) );
  AO222X1 U4703 ( .IN1(n5210), .IN2(rEIP_0_), .IN3(n5211), .IN4(n1415), .IN5(
        n5212), .IN6(n5213), .Q(n2430) );
  OA21X1 U4704 ( .IN1(n1416), .IN2(n2845), .IN3(n2888), .Q(n5211) );
  INVX0 U4705 ( .IN(n5214), .QN(n5210) );
  MUX21X1 U4706 ( .IN1(n5213), .IN2(BE_n[2]), .S(n3205), .Q(n2429) );
  NAND3X0 U4707 ( .IN1(n5214), .IN2(n5208), .IN3(n5215), .QN(n2428) );
  NAND2X0 U4708 ( .IN1(n5212), .IN2(n5216), .QN(n5215) );
  NAND3X0 U4709 ( .IN1(n1415), .IN2(n2845), .IN3(n1416), .QN(n5208) );
  MUX21X1 U4710 ( .IN1(n5216), .IN2(BE_n[1]), .S(n3205), .Q(n2427) );
  NAND2X0 U4711 ( .IN1(n5217), .IN2(n5214), .QN(n2426) );
  NAND2X0 U4712 ( .IN1(rEIP_1_), .IN2(n5207), .QN(n5214) );
  MUX21X1 U4713 ( .IN1(n2845), .IN2(n3692), .S(n5212), .Q(n5217) );
  INVX0 U4714 ( .IN(n5207), .QN(n5212) );
  NAND2X0 U4715 ( .IN1(n2864), .IN2(test_so2), .QN(n5207) );
  MUX21X1 U4716 ( .IN1(n5218), .IN2(BE_n[0]), .S(n3206), .Q(n2425) );
  AND2X1 U4717 ( .IN1(n4814), .IN2(n4030), .Q(n4024) );
  NAND3X0 U4718 ( .IN1(n2867), .IN2(n2847), .IN3(n1436), .QN(n4030) );
  NAND2X0 U4719 ( .IN1(n3874), .IN2(n5219), .QN(N811) );
  OAI21X1 U4720 ( .IN1(n5220), .IN2(n5221), .IN3(Datai[31]), .QN(n5219) );
  OR4X1 U4721 ( .IN1(Datai[16]), .IN2(Datai[17]), .IN3(Datai[18]), .IN4(
        Datai[19]), .Q(n5221) );
  OR4X1 U4722 ( .IN1(Datai[20]), .IN2(Datai[21]), .IN3(Datai[22]), .IN4(
        Datai[23]), .Q(n5220) );
  NAND2X0 U4723 ( .IN1(Datai[31]), .IN2(n5222), .QN(n3874) );
  OR4X1 U4724 ( .IN1(n5223), .IN2(n5224), .IN3(n5225), .IN4(n5226), .Q(n5222)
         );
  OR4X1 U4725 ( .IN1(n3084), .IN2(n3086), .IN3(n3088), .IN4(n3090), .Q(n5226)
         );
  OR4X1 U4726 ( .IN1(n3092), .IN2(n3094), .IN3(n2941), .IN4(n2945), .Q(n5225)
         );
  OR4X1 U4727 ( .IN1(n3080), .IN2(n2937), .IN3(n2943), .IN4(n2947), .Q(n5224)
         );
  OR4X1 U4728 ( .IN1(n2935), .IN2(n2939), .IN3(Datai[15]), .IN4(n3082), .Q(
        n5223) );
  NOR2X0 U4729 ( .IN1(n3871), .IN2(n2870), .QN(N3493) );
  AO21X1 U4730 ( .IN1(rEIP_1_), .IN2(rEIP_31_), .IN3(N498), .Q(N425) );
  NOR2X0 U4731 ( .IN1(n2845), .IN2(n2866), .QN(N498) );
  MUX21X1 U4732 ( .IN1(N2737), .IN2(n1557), .S(n2870), .Q(N3486) );
  MUX21X1 U4733 ( .IN1(n4137), .IN2(InstQueueRd_Addr[1]), .S(n1590), .Q(N3485)
         );
  NOR2X0 U4734 ( .IN1(n1557), .IN2(n4143), .QN(n4137) );
  INVX0 U4735 ( .IN(n5227), .QN(n4143) );
  MUX21X1 U4736 ( .IN1(n5228), .IN2(n4140), .S(n1590), .Q(N3484) );
  NOR2X0 U4737 ( .IN1(n1557), .IN2(n5227), .QN(n5228) );
  XOR2X1 U4738 ( .IN1(n3867), .IN2(N3467), .Q(n5227) );
  MUX21X1 U4739 ( .IN1(N2737), .IN2(n4134), .S(n5066), .Q(N3420) );
  AO21X1 U4740 ( .IN1(N2737), .IN2(n5229), .IN3(n5230), .Q(n4134) );
  MUX21X1 U4741 ( .IN1(n5231), .IN2(n4658), .S(n1552), .Q(n5230) );
  MUX21X1 U4742 ( .IN1(n4138), .IN2(InstQueueRd_Addr[1]), .S(n5232), .Q(N3419)
         );
  AO222X1 U4743 ( .IN1(n1550), .IN2(n5231), .IN3(n4136), .IN4(n4658), .IN5(
        n1550), .IN6(n5229), .Q(n4138) );
  NAND2X0 U4744 ( .IN1(n5063), .IN2(n5062), .QN(n4658) );
  NAND2X0 U4745 ( .IN1(n3996), .IN2(n3887), .QN(n4136) );
  MUX21X1 U4746 ( .IN1(n4144), .IN2(n4140), .S(n5232), .Q(N3418) );
  AO221X1 U4747 ( .IN1(n5233), .IN2(n5231), .IN3(N2739), .IN4(n5229), .IN5(
        n5234), .Q(n4144) );
  MUX21X1 U4748 ( .IN1(n5235), .IN2(n5236), .S(n4141), .Q(n5234) );
  XOR2X1 U4749 ( .IN1(n3839), .IN2(n3889), .Q(n4141) );
  XOR2X1 U4750 ( .IN1(n3839), .IN2(n1550), .Q(n5233) );
  MUX21X1 U4751 ( .IN1(n4080), .IN2(n4078), .S(n5232), .Q(N3417) );
  AO221X1 U4752 ( .IN1(n5237), .IN2(n5231), .IN3(n5238), .IN4(n5235), .IN5(
        n5239), .Q(n4080) );
  AO22X1 U4753 ( .IN1(N2740), .IN2(n5229), .IN3(n5236), .IN4(n4082), .Q(n5239)
         );
  NAND2X0 U4754 ( .IN1(n5240), .IN2(n3111), .QN(n4082) );
  MUX21X1 U4755 ( .IN1(n3124), .IN2(n1548), .S(n3889), .Q(n5240) );
  INVX0 U4756 ( .IN(n5062), .QN(n5236) );
  NAND2X0 U4757 ( .IN1(n5241), .IN2(n3124), .QN(n5238) );
  MUX21X1 U4758 ( .IN1(n4078), .IN2(n3110), .S(n3889), .Q(n5241) );
  NAND2X0 U4759 ( .IN1(n5242), .IN2(n3111), .QN(n5237) );
  MUX21X1 U4760 ( .IN1(n3124), .IN2(n1548), .S(n1550), .Q(n5242) );
  MUX21X1 U4761 ( .IN1(n5243), .IN2(InstQueueRd_Addr[4]), .S(n5232), .Q(N3427)
         );
  INVX0 U4762 ( .IN(n5066), .QN(n5232) );
  NAND4X0 U4763 ( .IN1(n5244), .IN2(n5245), .IN3(n5062), .IN4(n5246), .QN(
        n5066) );
  NAND3X0 U4764 ( .IN1(n5247), .IN2(n5199), .IN3(n5061), .QN(n5062) );
  NOR2X0 U4765 ( .IN1(n5231), .IN2(n5229), .QN(n5061) );
  INVX0 U4766 ( .IN(n4148), .QN(n5229) );
  NAND3X0 U4767 ( .IN1(n5246), .IN2(n4812), .IN3(n4020), .QN(n5231) );
  INVX0 U4768 ( .IN(n5206), .QN(n4020) );
  INVX0 U4769 ( .IN(n4656), .QN(n5246) );
  NOR4X0 U4770 ( .IN1(n4129), .IN2(n4124), .IN3(n4628), .IN4(n4126), .QN(n4656) );
  NAND4X0 U4771 ( .IN1(n4644), .IN2(n5248), .IN3(n5249), .IN4(n5250), .QN(
        n4129) );
  NAND2X0 U4772 ( .IN1(n5251), .IN2(n5252), .QN(n5199) );
  INVX0 U4773 ( .IN(n4662), .QN(n5247) );
  NAND2X0 U4774 ( .IN1(n5063), .IN2(n5064), .QN(n4662) );
  NAND3X0 U4775 ( .IN1(n4126), .IN2(n5253), .IN3(n5251), .QN(n5064) );
  INVX0 U4776 ( .IN(n5235), .QN(n5063) );
  NAND3X0 U4777 ( .IN1(n4659), .IN2(n2948), .IN3(n4651), .QN(n5245) );
  INVX0 U4778 ( .IN(n4661), .QN(n4651) );
  AO21X1 U4779 ( .IN1(n5201), .IN2(n5254), .IN3(n2955), .Q(n4661) );
  INVX0 U4780 ( .IN(r680_B_1_), .QN(n5254) );
  NOR3X0 U4781 ( .IN1(r680_B_3_), .IN2(r680_B_4_), .IN3(r680_B_2_), .QN(n5201)
         );
  AO21X1 U4782 ( .IN1(n5206), .IN2(n4019), .IN3(n4869), .Q(n4659) );
  NAND2X0 U4783 ( .IN1(n4148), .IN2(n4812), .QN(n4869) );
  NAND3X0 U4784 ( .IN1(n4125), .IN2(n5250), .IN3(n5255), .QN(n4812) );
  NAND2X0 U4785 ( .IN1(n4040), .IN2(n4814), .QN(n4019) );
  NAND3X0 U4786 ( .IN1(n1434), .IN2(n2847), .IN3(n1436), .QN(n4814) );
  NAND3X0 U4787 ( .IN1(n1436), .IN2(n2867), .IN3(n1435), .QN(n4040) );
  NAND2X0 U4788 ( .IN1(n4822), .IN2(n4021), .QN(n5206) );
  NAND4X0 U4789 ( .IN1(n4126), .IN2(n5256), .IN3(n4125), .IN4(n5250), .QN(
        n4021) );
  INVX0 U4790 ( .IN(n4638), .QN(n4125) );
  NAND2X0 U4791 ( .IN1(n5257), .IN2(n4628), .QN(n4822) );
  NAND2X0 U4792 ( .IN1(n4868), .IN2(n5235), .QN(n5244) );
  NAND2X0 U4793 ( .IN1(n4120), .IN2(n4863), .QN(n5235) );
  NAND4X0 U4794 ( .IN1(n4638), .IN2(n4641), .IN3(n5256), .IN4(n4870), .QN(
        n4863) );
  AND3X1 U4795 ( .IN1(n5253), .IN2(n5258), .IN3(n4647), .Q(n5256) );
  AND3X1 U4796 ( .IN1(n4128), .IN2(n5248), .IN3(n4635), .Q(n5253) );
  INVX0 U4797 ( .IN(n4631), .QN(n5248) );
  NAND3X0 U4798 ( .IN1(n4641), .IN2(n5255), .IN3(n4638), .QN(n4120) );
  AND3X1 U4799 ( .IN1(n4647), .IN2(n5258), .IN3(n5252), .Q(n5255) );
  NOR4X0 U4800 ( .IN1(n4128), .IN2(n4870), .IN3(n5249), .IN4(n4631), .QN(n5252) );
  ISOLANDX1 U4801 ( .D(n5259), .ISO(n2955), .Q(n4868) );
  OR3X1 U4802 ( .IN1(r680_B_3_), .IN2(r680_B_4_), .IN3(n5260), .Q(n5259) );
  OA21X1 U4803 ( .IN1(r680_B_1_), .IN2(gte_355_B_0_), .IN3(r680_B_2_), .Q(
        n5260) );
  NOR2X0 U4804 ( .IN1(n4148), .IN2(n2883), .QN(n5243) );
  NAND2X0 U4805 ( .IN1(n5257), .IN2(n4128), .QN(n4148) );
  INVX0 U4806 ( .IN(n4628), .QN(n4128) );
  OA222X1 U4807 ( .IN1(n3903), .IN2(n3996), .IN3(n5261), .IN4(n3998), .IN5(
        n1552), .IN6(n3907), .Q(n4628) );
  MUX21X1 U4808 ( .IN1(n3900), .IN2(n5262), .S(n1550), .Q(n3907) );
  OA221X1 U4809 ( .IN1(n3107), .IN2(n4461), .IN3(n3121), .IN4(n4349), .IN5(
        n5263), .Q(n5262) );
  OA22X1 U4810 ( .IN1(n3141), .IN2(n4574), .IN3(n3165), .IN4(n4234), .Q(n5263)
         );
  AOI221X1 U4811 ( .IN1(n3751), .IN2(n3128), .IN3(n3783), .IN4(n3116), .IN5(
        n5264), .QN(n3900) );
  AO22X1 U4812 ( .IN1(n3719), .IN2(n3162), .IN3(n3815), .IN4(n3150), .Q(n5264)
         );
  OA221X1 U4813 ( .IN1(n3107), .IN2(n4430), .IN3(n3122), .IN4(n4317), .IN5(
        n5265), .Q(n5261) );
  OA22X1 U4814 ( .IN1(n3142), .IN2(n4541), .IN3(n3165), .IN4(N2549), .Q(n5265)
         );
  AOI221X1 U4815 ( .IN1(n3743), .IN2(n3128), .IN3(n3775), .IN4(n3116), .IN5(
        n5266), .QN(n3903) );
  AO22X1 U4816 ( .IN1(n3711), .IN2(n3163), .IN3(n3807), .IN4(n3139), .Q(n5266)
         );
  AND4X1 U4817 ( .IN1(n5251), .IN2(n4631), .IN3(n5249), .IN4(n4870), .Q(n5257)
         );
  INVX0 U4818 ( .IN(n4126), .QN(n4870) );
  OA222X1 U4819 ( .IN1(n3880), .IN2(n3996), .IN3(n5267), .IN4(n3998), .IN5(
        n1552), .IN6(n3886), .Q(n4126) );
  MUX21X1 U4820 ( .IN1(n3876), .IN2(n5268), .S(n1550), .Q(n3886) );
  OA221X1 U4821 ( .IN1(test_so9), .IN2(n3164), .IN3(n3140), .IN4(n4570), .IN5(
        n5269), .Q(n5268) );
  OA22X1 U4822 ( .IN1(n4345), .IN2(n3124), .IN3(n4457), .IN4(n3111), .Q(n5269)
         );
  AOI221X1 U4823 ( .IN1(n3750), .IN2(n3128), .IN3(n3782), .IN4(n3116), .IN5(
        n5270), .QN(n3876) );
  AO22X1 U4824 ( .IN1(n3718), .IN2(n3162), .IN3(n3814), .IN4(n3137), .Q(n5270)
         );
  OA221X1 U4825 ( .IN1(n3108), .IN2(n4426), .IN3(n3122), .IN4(n4313), .IN5(
        n5271), .Q(n5267) );
  OA22X1 U4826 ( .IN1(n3142), .IN2(n4537), .IN3(n3165), .IN4(N2548), .Q(n5271)
         );
  AOI221X1 U4827 ( .IN1(n3742), .IN2(n3129), .IN3(n3774), .IN4(n3116), .IN5(
        n5272), .QN(n3880) );
  AO22X1 U4828 ( .IN1(n3710), .IN2(n3163), .IN3(n3806), .IN4(n3137), .Q(n5272)
         );
  INVX0 U4829 ( .IN(n4635), .QN(n5249) );
  OA222X1 U4830 ( .IN1(n3933), .IN2(n3996), .IN3(n5273), .IN4(n3998), .IN5(
        n1552), .IN6(n3937), .Q(n4635) );
  MUX21X1 U4831 ( .IN1(n5274), .IN2(n3930), .S(InstQueueRd_Addr[1]), .Q(n3937)
         );
  AOI221X1 U4832 ( .IN1(n3753), .IN2(n3129), .IN3(n3785), .IN4(n3116), .IN5(
        n5275), .QN(n3930) );
  AO22X1 U4833 ( .IN1(n3721), .IN2(n3175), .IN3(n3817), .IN4(n3154), .Q(n5275)
         );
  OA221X1 U4834 ( .IN1(n3108), .IN2(n4467), .IN3(n3122), .IN4(n4355), .IN5(
        n5276), .Q(n5274) );
  OA22X1 U4835 ( .IN1(n3142), .IN2(n4580), .IN3(n3166), .IN4(n4241), .Q(n5276)
         );
  OA221X1 U4836 ( .IN1(n3108), .IN2(n4436), .IN3(n3121), .IN4(n4323), .IN5(
        n5277), .Q(n5273) );
  OA22X1 U4837 ( .IN1(n3142), .IN2(n4547), .IN3(n3166), .IN4(N2551), .Q(n5277)
         );
  AOI221X1 U4838 ( .IN1(n3745), .IN2(n3126), .IN3(n3777), .IN4(n3112), .IN5(
        n5278), .QN(n3933) );
  AO22X1 U4839 ( .IN1(n3713), .IN2(n3175), .IN3(n3809), .IN4(n3154), .Q(n5278)
         );
  OA222X1 U4840 ( .IN1(n3918), .IN2(n3996), .IN3(n5279), .IN4(n3998), .IN5(
        n1552), .IN6(n3922), .Q(n4631) );
  MUX21X1 U4841 ( .IN1(n3915), .IN2(n5280), .S(n1550), .Q(n3922) );
  OA221X1 U4842 ( .IN1(n3108), .IN2(n4464), .IN3(n3121), .IN4(n4352), .IN5(
        n5281), .Q(n5280) );
  OA22X1 U4843 ( .IN1(n3143), .IN2(n4577), .IN3(n3166), .IN4(n4238), .Q(n5281)
         );
  AOI221X1 U4844 ( .IN1(n3752), .IN2(n3129), .IN3(n3784), .IN4(n3116), .IN5(
        n5282), .QN(n3915) );
  AO22X1 U4845 ( .IN1(n3720), .IN2(n3162), .IN3(n3816), .IN4(n3139), .Q(n5282)
         );
  OA221X1 U4846 ( .IN1(n3109), .IN2(n4433), .IN3(n3123), .IN4(n4320), .IN5(
        n5283), .Q(n5279) );
  OA22X1 U4847 ( .IN1(n3143), .IN2(n4544), .IN3(n3167), .IN4(N2550), .Q(n5283)
         );
  AOI221X1 U4848 ( .IN1(n3744), .IN2(n3129), .IN3(n3776), .IN4(n3112), .IN5(
        n5284), .QN(n3918) );
  AO22X1 U4849 ( .IN1(n3712), .IN2(n3163), .IN3(n3808), .IN4(n3149), .Q(n5284)
         );
  NOR4X0 U4850 ( .IN1(n5250), .IN2(n5258), .IN3(n4124), .IN4(n4638), .QN(n5251) );
  OA222X1 U4851 ( .IN1(n3948), .IN2(n3996), .IN3(n5285), .IN4(n3998), .IN5(
        n1552), .IN6(n3952), .Q(n4638) );
  MUX21X1 U4852 ( .IN1(n5286), .IN2(n3945), .S(InstQueueRd_Addr[1]), .Q(n3952)
         );
  AOI221X1 U4853 ( .IN1(n3754), .IN2(n3129), .IN3(n3786), .IN4(n3118), .IN5(
        n5287), .QN(n3945) );
  AO22X1 U4854 ( .IN1(n3722), .IN2(n3174), .IN3(n3818), .IN4(n3149), .Q(n5287)
         );
  OA221X1 U4855 ( .IN1(n3109), .IN2(n4471), .IN3(n3122), .IN4(n4359), .IN5(
        n5288), .Q(n5286) );
  OA22X1 U4856 ( .IN1(n3143), .IN2(n4584), .IN3(n3167), .IN4(n4244), .Q(n5288)
         );
  OA221X1 U4857 ( .IN1(n3109), .IN2(n4439), .IN3(n3123), .IN4(n4326), .IN5(
        n5289), .Q(n5285) );
  OA22X1 U4858 ( .IN1(n3143), .IN2(n4551), .IN3(n3167), .IN4(N2552), .Q(n5289)
         );
  AOI221X1 U4859 ( .IN1(n3746), .IN2(n3129), .IN3(n3778), .IN4(n3118), .IN5(
        n5290), .QN(n3948) );
  AO22X1 U4860 ( .IN1(n3714), .IN2(n3174), .IN3(n3810), .IN4(n3147), .Q(n5290)
         );
  INVX0 U4861 ( .IN(n4647), .QN(n4124) );
  OA222X1 U4862 ( .IN1(n3993), .IN2(n3996), .IN3(n5291), .IN4(n3998), .IN5(
        n1552), .IN6(n3999), .Q(n4647) );
  MUX21X1 U4863 ( .IN1(n5292), .IN2(n3990), .S(InstQueueRd_Addr[1]), .Q(n3999)
         );
  AOI221X1 U4864 ( .IN1(n3757), .IN2(n3130), .IN3(n3789), .IN4(n3117), .IN5(
        n5293), .QN(n3990) );
  AO22X1 U4865 ( .IN1(n3725), .IN2(n3173), .IN3(n3821), .IN4(n3148), .Q(n5293)
         );
  OA221X1 U4866 ( .IN1(n3109), .IN2(n4480), .IN3(n3123), .IN4(n4368), .IN5(
        n5294), .Q(n5292) );
  OA22X1 U4867 ( .IN1(n3144), .IN2(n4593), .IN3(n3168), .IN4(n4253), .Q(n5294)
         );
  OA221X1 U4868 ( .IN1(n3110), .IN2(test_so12), .IN3(n3122), .IN4(n4336), 
        .IN5(n5295), .Q(n5291) );
  OA22X1 U4869 ( .IN1(n3143), .IN2(n4560), .IN3(n3167), .IN4(N2555), .Q(n5295)
         );
  AOI221X1 U4870 ( .IN1(n3749), .IN2(n3130), .IN3(n3781), .IN4(n3117), .IN5(
        n5296), .QN(n3993) );
  AO22X1 U4871 ( .IN1(n3717), .IN2(n3173), .IN3(n3813), .IN4(n3148), .Q(n5296)
         );
  INVX0 U4872 ( .IN(n4644), .QN(n5258) );
  OA222X1 U4873 ( .IN1(n3978), .IN2(n3996), .IN3(n5297), .IN4(n3998), .IN5(
        n1552), .IN6(n3982), .Q(n4644) );
  MUX21X1 U4874 ( .IN1(n5298), .IN2(n3975), .S(InstQueueRd_Addr[1]), .Q(n3982)
         );
  AOI221X1 U4875 ( .IN1(n3756), .IN2(n3130), .IN3(n3788), .IN4(n3117), .IN5(
        n5299), .QN(n3975) );
  AO22X1 U4876 ( .IN1(n3724), .IN2(n3172), .IN3(n3820), .IN4(n3148), .Q(n5299)
         );
  OA221X1 U4877 ( .IN1(n3109), .IN2(n4477), .IN3(n3123), .IN4(n4365), .IN5(
        n5300), .Q(n5298) );
  OA22X1 U4878 ( .IN1(n3144), .IN2(n4590), .IN3(n3168), .IN4(n4250), .Q(n5300)
         );
  OA221X1 U4879 ( .IN1(n3110), .IN2(n4446), .IN3(n3124), .IN4(n4333), .IN5(
        n5301), .Q(n5297) );
  OA22X1 U4880 ( .IN1(n3144), .IN2(n4557), .IN3(n3168), .IN4(N2554), .Q(n5301)
         );
  AOI221X1 U4881 ( .IN1(n3748), .IN2(n3131), .IN3(n3780), .IN4(n3118), .IN5(
        n5302), .QN(n3978) );
  AO22X1 U4882 ( .IN1(n3716), .IN2(n3172), .IN3(n3812), .IN4(n3147), .Q(n5302)
         );
  INVX0 U4883 ( .IN(n4641), .QN(n5250) );
  OA222X1 U4884 ( .IN1(n3963), .IN2(n3996), .IN3(n5303), .IN4(n3998), .IN5(
        n1552), .IN6(n3967), .Q(n4641) );
  MUX21X1 U4885 ( .IN1(n5304), .IN2(n3960), .S(InstQueueRd_Addr[1]), .Q(n3967)
         );
  AOI221X1 U4886 ( .IN1(n3755), .IN2(n3131), .IN3(n3787), .IN4(n3118), .IN5(
        n5305), .QN(n3960) );
  AO22X1 U4887 ( .IN1(n3723), .IN2(n3171), .IN3(n3819), .IN4(n3147), .Q(n5305)
         );
  OA221X1 U4888 ( .IN1(n3110), .IN2(n4474), .IN3(n3123), .IN4(n4362), .IN5(
        n5306), .Q(n5304) );
  OA22X1 U4889 ( .IN1(n3144), .IN2(n4587), .IN3(n3168), .IN4(n4247), .Q(n5306)
         );
  OA221X1 U4890 ( .IN1(n3106), .IN2(n4443), .IN3(n3123), .IN4(n4330), .IN5(
        n5307), .Q(n5303) );
  OA22X1 U4891 ( .IN1(n3140), .IN2(n4554), .IN3(n3164), .IN4(N2553), .Q(n5307)
         );
  AOI221X1 U4892 ( .IN1(n3747), .IN2(n3131), .IN3(n3779), .IN4(n3118), .IN5(
        n5308), .QN(n3963) );
  AO22X1 U4893 ( .IN1(n3715), .IN2(n3171), .IN3(n3811), .IN4(n3148), .Q(n5308)
         );
  NAND2X0 U4894 ( .IN1(n4078), .IN2(n4140), .QN(n3896) );
  NAND2X0 U4895 ( .IN1(n3839), .IN2(n1548), .QN(n3897) );
  NAND2X0 U4896 ( .IN1(n3839), .IN2(n4078), .QN(n3893) );
  INVX0 U4897 ( .IN(n1548), .QN(n4078) );
  NAND2X0 U4898 ( .IN1(n1548), .IN2(n4140), .QN(n3894) );
  INVX0 U4899 ( .IN(n3839), .QN(n4140) );
  MUX21X1 U4900 ( .IN1(Datai[0]), .IN2(N3434), .S(n5309), .Q(N2103) );
  MUX21X1 U4901 ( .IN1(Datai[1]), .IN2(N3435), .S(n5309), .Q(N2104) );
  MUX21X1 U4902 ( .IN1(Datai[2]), .IN2(test_so17), .S(n5309), .Q(N2105) );
  MUX21X1 U4903 ( .IN1(Datai[3]), .IN2(N3437), .S(n5309), .Q(N2106) );
  MUX21X1 U4904 ( .IN1(Datai[4]), .IN2(N3438), .S(n5309), .Q(N2107) );
  MUX21X1 U4905 ( .IN1(Datai[5]), .IN2(N3439), .S(n5309), .Q(N2108) );
  MUX21X1 U4906 ( .IN1(Datai[6]), .IN2(N3440), .S(n5309), .Q(N2109) );
  MUX21X1 U4907 ( .IN1(Datai[7]), .IN2(N3441), .S(n5309), .Q(N2110) );
  MUX21X1 U4908 ( .IN1(n2941), .IN2(N3442), .S(n5309), .Q(N2111) );
  MUX21X1 U4909 ( .IN1(n2945), .IN2(N3443), .S(n5309), .Q(N2112) );
  MUX21X1 U4910 ( .IN1(n2937), .IN2(N3444), .S(n5309), .Q(N2113) );
  MUX21X1 U4911 ( .IN1(n2943), .IN2(N3445), .S(n5309), .Q(N2114) );
  MUX21X1 U4912 ( .IN1(n2947), .IN2(N3446), .S(n5309), .Q(N2115) );
  MUX21X1 U4913 ( .IN1(n2935), .IN2(N3447), .S(n5309), .Q(N2116) );
  MUX21X1 U4914 ( .IN1(n2939), .IN2(N3448), .S(n5309), .Q(N2117) );
  MUX21X1 U4915 ( .IN1(Datai[15]), .IN2(N3449), .S(n5309), .Q(N2118) );
  NOR2X0 U4916 ( .IN1(n3822), .IN2(n5310), .QN(N1749) );
  NOR4X0 U4917 ( .IN1(n5311), .IN2(n5312), .IN3(n5313), .IN4(n5314), .QN(n5310) );
  NAND4X0 U4918 ( .IN1(n3838), .IN2(n3837), .IN3(n3836), .IN4(n3835), .QN(
        n5314) );
  NAND4X0 U4919 ( .IN1(n3834), .IN2(n3833), .IN3(n3832), .IN4(n3831), .QN(
        n5313) );
  NAND4X0 U4920 ( .IN1(n3830), .IN2(n3829), .IN3(n3828), .IN4(n3827), .QN(
        n5312) );
  NAND4X0 U4921 ( .IN1(n3826), .IN2(n3825), .IN3(n3824), .IN4(n3823), .QN(
        n5311) );
endmodule

