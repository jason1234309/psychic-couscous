module top(
  input LIOB33_SING_X0Y100_IOB_X0Y100_IPAD,
  input LIOB33_X0Y101_IOB_X0Y101_IPAD,
  input LIOB33_X0Y101_IOB_X0Y102_IPAD,
  input LIOB33_X0Y103_IOB_X0Y103_IPAD,
  input LIOB33_X0Y103_IOB_X0Y104_IPAD,
  input LIOB33_X0Y105_IOB_X0Y105_IPAD,
  input LIOB33_X0Y105_IOB_X0Y106_IPAD,
  input LIOB33_X0Y107_IOB_X0Y107_IPAD,
  input LIOB33_X0Y107_IOB_X0Y108_IPAD,
  input LIOB33_X0Y109_IOB_X0Y109_IPAD,
  input LIOB33_X0Y109_IOB_X0Y110_IPAD,
  input LIOB33_X0Y111_IOB_X0Y111_IPAD,
  input LIOB33_X0Y111_IOB_X0Y112_IPAD,
  input LIOB33_X0Y113_IOB_X0Y113_IPAD,
  input LIOB33_X0Y113_IOB_X0Y114_IPAD,
  input LIOB33_X0Y115_IOB_X0Y115_IPAD,
  input LIOB33_X0Y115_IOB_X0Y116_IPAD,
  input LIOB33_X0Y117_IOB_X0Y117_IPAD,
  input LIOB33_X0Y117_IOB_X0Y118_IPAD,
  input LIOB33_X0Y119_IOB_X0Y119_IPAD,
  input LIOB33_X0Y119_IOB_X0Y120_IPAD,
  input LIOB33_X0Y121_IOB_X0Y121_IPAD,
  input LIOB33_X0Y121_IOB_X0Y122_IPAD,
  input LIOB33_X0Y123_IOB_X0Y123_IPAD,
  input RIOB33_SING_X105Y100_IOB_X1Y100_IPAD,
  input RIOB33_X105Y101_IOB_X1Y101_IPAD,
  input RIOB33_X105Y101_IOB_X1Y102_IPAD,
  input RIOB33_X105Y103_IOB_X1Y103_IPAD,
  input RIOB33_X105Y103_IOB_X1Y104_IPAD,
  input RIOB33_X105Y105_IOB_X1Y105_IPAD,
  input RIOB33_X105Y105_IOB_X1Y106_IPAD,
  input RIOB33_X105Y127_IOB_X1Y128_IPAD,
  output LIOB33_SING_X0Y149_IOB_X0Y149_OPAD,
  output LIOB33_X0Y123_IOB_X0Y124_OPAD,
  output LIOB33_X0Y125_IOB_X0Y125_OPAD,
  output LIOB33_X0Y125_IOB_X0Y126_OPAD,
  output LIOB33_X0Y127_IOB_X0Y127_OPAD,
  output LIOB33_X0Y127_IOB_X0Y128_OPAD,
  output LIOB33_X0Y129_IOB_X0Y129_OPAD,
  output LIOB33_X0Y129_IOB_X0Y130_OPAD,
  output LIOB33_X0Y131_IOB_X0Y131_OPAD,
  output LIOB33_X0Y131_IOB_X0Y132_OPAD,
  output LIOB33_X0Y133_IOB_X0Y133_OPAD,
  output LIOB33_X0Y133_IOB_X0Y134_OPAD,
  output LIOB33_X0Y135_IOB_X0Y135_OPAD,
  output LIOB33_X0Y135_IOB_X0Y136_OPAD,
  output LIOB33_X0Y137_IOB_X0Y137_OPAD,
  output LIOB33_X0Y137_IOB_X0Y138_OPAD,
  output LIOB33_X0Y139_IOB_X0Y139_OPAD,
  output LIOB33_X0Y139_IOB_X0Y140_OPAD,
  output LIOB33_X0Y141_IOB_X0Y141_OPAD,
  output LIOB33_X0Y141_IOB_X0Y142_OPAD,
  output LIOB33_X0Y143_IOB_X0Y143_OPAD,
  output LIOB33_X0Y145_IOB_X0Y145_OPAD,
  output LIOB33_X0Y145_IOB_X0Y146_OPAD,
  output LIOB33_X0Y147_IOB_X0Y147_OPAD,
  output LIOB33_X0Y147_IOB_X0Y148_OPAD,
  output RIOB33_X105Y107_IOB_X1Y107_OPAD,
  output RIOB33_X105Y107_IOB_X1Y108_OPAD,
  output RIOB33_X105Y109_IOB_X1Y109_OPAD,
  output RIOB33_X105Y109_IOB_X1Y110_OPAD,
  output RIOB33_X105Y111_IOB_X1Y111_OPAD,
  output RIOB33_X105Y111_IOB_X1Y112_OPAD,
  output RIOB33_X105Y113_IOB_X1Y113_OPAD,
  output RIOB33_X105Y113_IOB_X1Y114_OPAD,
  output RIOB33_X105Y115_IOB_X1Y115_OPAD,
  output RIOB33_X105Y115_IOB_X1Y116_OPAD,
  output RIOB33_X105Y117_IOB_X1Y117_OPAD,
  output RIOB33_X105Y117_IOB_X1Y118_OPAD,
  output RIOB33_X105Y119_IOB_X1Y119_OPAD,
  output RIOB33_X105Y119_IOB_X1Y120_OPAD,
  output RIOB33_X105Y121_IOB_X1Y121_OPAD,
  output RIOB33_X105Y121_IOB_X1Y122_OPAD,
  output RIOB33_X105Y123_IOB_X1Y123_OPAD,
  output RIOB33_X105Y123_IOB_X1Y124_OPAD,
  output RIOB33_X105Y125_IOB_X1Y125_OPAD,
  output RIOB33_X105Y125_IOB_X1Y126_OPAD,
  output RIOB33_X105Y127_IOB_X1Y127_OPAD,
  output RIOB33_X105Y129_IOB_X1Y129_OPAD,
  output RIOB33_X105Y129_IOB_X1Y130_OPAD,
  output RIOB33_X105Y131_IOB_X1Y131_OPAD,
  output RIOB33_X105Y131_IOB_X1Y132_OPAD,
  output RIOB33_X105Y133_IOB_X1Y133_OPAD,
  output RIOB33_X105Y133_IOB_X1Y134_OPAD,
  output RIOB33_X105Y135_IOB_X1Y135_OPAD,
  output RIOB33_X105Y135_IOB_X1Y136_OPAD,
  output RIOB33_X105Y137_IOB_X1Y137_OPAD,
  output RIOB33_X105Y137_IOB_X1Y138_OPAD,
  output RIOB33_X105Y139_IOB_X1Y139_OPAD,
  output RIOB33_X105Y139_IOB_X1Y140_OPAD,
  output RIOB33_X105Y141_IOB_X1Y141_OPAD,
  output RIOB33_X105Y141_IOB_X1Y142_OPAD,
  output RIOB33_X105Y143_IOB_X1Y143_OPAD,
  output RIOB33_X105Y143_IOB_X1Y144_OPAD,
  output RIOB33_X105Y145_IOB_X1Y145_OPAD
  );
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_A;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_A1;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_A2;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_A3;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_A4;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_A5;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_A6;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_AO5;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_AO6;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_A_CY;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_A_XOR;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_B;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_B1;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_B2;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_B3;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_B4;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_B5;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_B6;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_BO5;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_BO6;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_B_CY;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_B_XOR;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_C;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_C1;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_C2;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_C3;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_C4;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_C5;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_C6;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_CO5;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_CO6;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_C_CY;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_C_XOR;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_D;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_D1;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_D2;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_D3;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_D4;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_D5;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_D6;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_DO5;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_DO6;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_D_CY;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X78Y101_D_XOR;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_A;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_A1;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_A2;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_A3;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_A4;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_A5;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_A6;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_AO5;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_AO6;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_A_CY;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_A_XOR;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_B;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_B1;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_B2;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_B3;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_B4;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_B5;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_B6;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_BO5;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_BO6;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_B_CY;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_B_XOR;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_C;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_C1;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_C2;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_C3;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_C4;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_C5;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_C6;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_CO5;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_CO6;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_C_CY;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_C_XOR;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_D;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_D1;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_D2;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_D3;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_D4;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_D5;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_D6;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_DO5;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_DO6;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_D_CY;
  wire [0:0] CLBLL_L_X52Y101_SLICE_X79Y101_D_XOR;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_A;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_A1;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_A2;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_A3;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_A4;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_A5;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_A6;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_AMUX;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_AO5;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_AO6;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_A_CY;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_A_XOR;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_B;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_B1;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_B2;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_B3;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_B4;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_B5;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_B6;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_BMUX;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_BO5;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_BO6;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_B_CY;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_B_XOR;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_C;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_C1;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_C2;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_C3;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_C4;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_C5;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_C6;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_CO5;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_CO6;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_C_CY;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_C_XOR;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_D;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_D1;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_D2;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_D3;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_D4;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_D5;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_D6;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_DO5;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_DO6;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_D_CY;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X78Y105_D_XOR;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_A;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_A1;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_A2;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_A3;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_A4;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_A5;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_A6;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_AO5;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_AO6;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_A_CY;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_A_XOR;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_B;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_B1;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_B2;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_B3;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_B4;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_B5;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_B6;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_BO5;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_BO6;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_B_CY;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_B_XOR;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_C;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_C1;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_C2;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_C3;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_C4;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_C5;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_C6;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_CO5;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_CO6;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_C_CY;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_C_XOR;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_D;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_D1;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_D2;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_D3;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_D4;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_D5;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_D6;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_DO5;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_DO6;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_D_CY;
  wire [0:0] CLBLL_L_X52Y105_SLICE_X79Y105_D_XOR;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_A;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_A1;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_A2;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_A3;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_A4;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_A5;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_A6;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_AMUX;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_AO5;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_AO6;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_A_CY;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_A_XOR;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_B;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_B1;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_B2;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_B3;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_B4;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_B5;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_B6;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_BO5;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_BO6;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_B_CY;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_B_XOR;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_C;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_C1;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_C2;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_C3;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_C4;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_C5;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_C6;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_CO5;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_CO6;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_C_CY;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_C_XOR;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_D;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_D1;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_D2;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_D3;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_D4;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_D5;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_D6;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_DO5;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_DO6;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_D_CY;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X78Y106_D_XOR;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_A;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_A1;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_A2;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_A3;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_A4;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_A5;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_A6;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_AMUX;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_AO5;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_AO6;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_A_CY;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_A_XOR;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_B;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_B1;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_B2;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_B3;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_B4;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_B5;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_B6;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_BO5;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_BO6;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_B_CY;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_B_XOR;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_C;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_C1;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_C2;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_C3;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_C4;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_C5;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_C6;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_CO5;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_CO6;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_C_CY;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_C_XOR;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_D;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_D1;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_D2;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_D3;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_D4;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_D5;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_D6;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_DO5;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_DO6;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_D_CY;
  wire [0:0] CLBLL_L_X52Y106_SLICE_X79Y106_D_XOR;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_A;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_A1;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_A2;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_A3;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_A4;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_A5;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_A6;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_AMUX;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_AO5;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_AO6;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_A_CY;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_A_XOR;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_B;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_B1;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_B2;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_B3;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_B4;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_B5;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_B6;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_BMUX;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_BO5;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_BO6;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_B_CY;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_B_XOR;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_C;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_C1;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_C2;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_C3;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_C4;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_C5;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_C6;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_CO5;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_CO6;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_C_CY;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_C_XOR;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_D;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_D1;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_D2;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_D3;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_D4;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_D5;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_D6;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_DO5;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_DO6;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_D_CY;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X78Y107_D_XOR;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_A;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_A1;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_A2;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_A3;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_A4;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_A5;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_A6;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_AO5;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_AO6;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_A_CY;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_A_XOR;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_B;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_B1;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_B2;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_B3;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_B4;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_B5;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_B6;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_BO5;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_BO6;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_B_CY;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_B_XOR;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_C;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_C1;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_C2;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_C3;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_C4;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_C5;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_C6;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_CO5;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_CO6;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_C_CY;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_C_XOR;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_D;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_D1;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_D2;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_D3;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_D4;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_D5;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_D6;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_DO5;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_DO6;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_D_CY;
  wire [0:0] CLBLL_L_X52Y107_SLICE_X79Y107_D_XOR;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_A;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_A1;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_A2;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_A3;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_A4;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_A5;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_A6;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_AO5;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_AO6;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_A_CY;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_A_XOR;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_B;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_B1;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_B2;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_B3;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_B4;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_B5;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_B6;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_BO5;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_BO6;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_B_CY;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_B_XOR;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_C;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_C1;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_C2;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_C3;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_C4;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_C5;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_C6;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_CO5;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_CO6;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_C_CY;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_C_XOR;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_D;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_D1;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_D2;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_D3;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_D4;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_D5;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_D6;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_DO5;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_DO6;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_D_CY;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X78Y99_D_XOR;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_A;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_A1;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_A2;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_A3;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_A4;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_A5;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_A6;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_AMUX;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_AO5;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_AO6;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_A_CY;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_A_XOR;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_B;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_B1;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_B2;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_B3;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_B4;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_B5;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_B6;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_BO5;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_BO6;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_B_CY;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_B_XOR;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_C;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_C1;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_C2;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_C3;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_C4;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_C5;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_C6;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_CO5;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_CO6;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_C_CY;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_C_XOR;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_D;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_D1;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_D2;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_D3;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_D4;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_D5;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_D6;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_DO5;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_DO6;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_D_CY;
  wire [0:0] CLBLL_L_X52Y99_SLICE_X79Y99_D_XOR;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_A;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_A1;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_A2;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_A3;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_A4;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_A5;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_A6;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_AMUX;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_AO5;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_AO6;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_A_CY;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_A_XOR;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_B;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_B1;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_B2;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_B3;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_B4;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_B5;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_B6;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_BO5;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_BO6;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_BQ;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_B_CY;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_B_XOR;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_C;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_C1;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_C2;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_C3;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_C4;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_C5;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_C6;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_CE;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_CLK;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_CO5;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_CO6;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_C_CY;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_C_XOR;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_D;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_D1;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_D2;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_D3;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_D4;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_D5;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_D6;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_DO5;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_DO6;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_D_CY;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_D_XOR;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X82Y100_SR;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_A;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_A1;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_A2;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_A3;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_A4;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_A5;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_A6;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_AMUX;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_AO5;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_AO6;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_A_CY;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_A_XOR;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_B;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_B1;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_B2;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_B3;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_B4;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_B5;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_B6;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_BO5;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_BO6;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_B_CY;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_B_XOR;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_C;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_C1;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_C2;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_C3;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_C4;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_C5;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_C6;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_CO5;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_CO6;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_C_CY;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_C_XOR;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_D;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_D1;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_D2;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_D3;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_D4;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_D5;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_D6;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_DO5;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_DO6;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_D_CY;
  wire [0:0] CLBLL_L_X54Y100_SLICE_X83Y100_D_XOR;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_A;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_A1;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_A2;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_A3;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_A4;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_A5;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_A6;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_AMUX;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_AO5;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_AO6;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_AQ;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_A_CY;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_A_XOR;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_B;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_B1;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_B2;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_B3;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_B4;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_B5;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_B6;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_BO5;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_BO6;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_BQ;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_BX;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_B_CY;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_B_XOR;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_C;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_C1;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_C2;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_C3;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_C4;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_C5;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_C6;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_CE;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_CLK;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_CO5;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_CO6;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_C_CY;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_C_XOR;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_D;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_D1;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_D2;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_D3;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_D4;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_D5;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_D6;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_DO5;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_DO6;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_D_CY;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_D_XOR;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X82Y101_SR;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_A;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_A1;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_A2;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_A3;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_A4;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_A5;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_A6;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_AO5;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_AO6;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_A_CY;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_A_XOR;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_B;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_B1;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_B2;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_B3;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_B4;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_B5;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_B6;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_BO5;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_BO6;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_B_CY;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_B_XOR;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_C;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_C1;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_C2;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_C3;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_C4;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_C5;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_C6;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_CO5;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_CO6;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_C_CY;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_C_XOR;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_D;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_D1;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_D2;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_D3;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_D4;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_D5;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_D6;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_DO5;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_DO6;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_D_CY;
  wire [0:0] CLBLL_L_X54Y101_SLICE_X83Y101_D_XOR;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_A;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_A1;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_A2;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_A3;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_A4;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_A5;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_A6;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_AMUX;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_AO5;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_AO6;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_A_CY;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_A_XOR;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_B;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_B1;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_B2;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_B3;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_B4;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_B5;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_B6;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_BO5;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_BO6;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_B_CY;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_B_XOR;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_C;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_C1;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_C2;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_C3;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_C4;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_C5;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_C6;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_CO5;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_CO6;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_C_CY;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_C_XOR;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_D;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_D1;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_D2;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_D3;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_D4;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_D5;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_D6;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_DO5;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_DO6;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_D_CY;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X82Y102_D_XOR;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_A;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_A1;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_A2;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_A3;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_A4;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_A5;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_A6;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_AO5;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_AO6;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_A_CY;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_A_XOR;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_B;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_B1;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_B2;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_B3;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_B4;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_B5;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_B6;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_BO5;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_BO6;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_B_CY;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_B_XOR;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_C;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_C1;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_C2;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_C3;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_C4;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_C5;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_C6;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_CO5;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_CO6;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_C_CY;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_C_XOR;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_D;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_D1;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_D2;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_D3;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_D4;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_D5;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_D6;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_DO5;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_DO6;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_D_CY;
  wire [0:0] CLBLL_L_X54Y102_SLICE_X83Y102_D_XOR;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_A;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_A1;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_A2;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_A3;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_A4;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_A5;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_A6;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_AO5;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_AO6;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_AQ;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_A_CY;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_A_XOR;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_B;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_B1;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_B2;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_B3;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_B4;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_B5;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_B6;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_BO5;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_BO6;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_B_CY;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_B_XOR;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_C;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_C1;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_C2;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_C3;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_C4;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_C5;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_C6;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_CLK;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_CO5;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_CO6;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_C_CY;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_C_XOR;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_D;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_D1;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_D2;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_D3;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_D4;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_D5;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_D6;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_DO5;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_DO6;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_D_CY;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_D_XOR;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X82Y103_SR;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_A;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_A1;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_A2;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_A3;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_A4;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_A5;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_A6;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_AO5;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_AO6;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_A_CY;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_A_XOR;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_B;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_B1;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_B2;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_B3;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_B4;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_B5;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_B6;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_BO5;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_BO6;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_B_CY;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_B_XOR;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_C;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_C1;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_C2;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_C3;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_C4;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_C5;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_C6;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_CO5;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_CO6;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_C_CY;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_C_XOR;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_D;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_D1;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_D2;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_D3;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_D4;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_D5;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_D6;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_DO5;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_DO6;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_D_CY;
  wire [0:0] CLBLL_L_X54Y103_SLICE_X83Y103_D_XOR;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_A;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_A1;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_A2;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_A3;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_A4;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_A5;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_A6;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_AO5;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_AO6;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_A_CY;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_A_XOR;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_B;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_B1;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_B2;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_B3;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_B4;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_B5;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_B6;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_BO5;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_BO6;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_B_CY;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_B_XOR;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_C;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_C1;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_C2;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_C3;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_C4;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_C5;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_C6;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_CO5;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_CO6;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_C_CY;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_C_XOR;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_D;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_D1;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_D2;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_D3;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_D4;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_D5;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_D6;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_DO5;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_DO6;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_D_CY;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X82Y104_D_XOR;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_A;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_A1;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_A2;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_A3;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_A4;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_A5;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_A6;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_AO5;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_AO6;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_A_CY;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_A_XOR;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_B;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_B1;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_B2;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_B3;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_B4;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_B5;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_B6;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_BO5;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_BO6;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_B_CY;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_B_XOR;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_C;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_C1;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_C2;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_C3;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_C4;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_C5;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_C6;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_CO5;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_CO6;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_C_CY;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_C_XOR;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_D;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_D1;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_D2;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_D3;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_D4;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_D5;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_D6;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_DO5;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_DO6;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_D_CY;
  wire [0:0] CLBLL_L_X54Y104_SLICE_X83Y104_D_XOR;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_A;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_A1;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_A2;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_A3;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_A4;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_A5;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_A6;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_AO5;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_AO6;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_AX;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_A_CY;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_A_XOR;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_B;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_B1;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_B2;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_B3;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_B4;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_B5;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_B6;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_BMUX;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_BO5;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_BO6;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_BX;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_B_CY;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_B_XOR;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_C;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_C1;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_C2;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_C3;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_C4;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_C5;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_C6;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_CMUX;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_CO5;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_CO6;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_COUT;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_CX;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_C_CY;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_C_XOR;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_D;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_D1;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_D2;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_D3;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_D4;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_D5;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_D6;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_DMUX;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_DO5;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_DO6;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_D_CY;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X82Y105_D_XOR;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_A;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_A1;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_A2;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_A3;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_A4;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_A5;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_A6;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_AO5;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_AO6;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_A_CY;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_A_XOR;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_B;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_B1;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_B2;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_B3;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_B4;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_B5;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_B6;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_BO5;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_BO6;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_B_CY;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_B_XOR;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_C;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_C1;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_C2;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_C3;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_C4;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_C5;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_C6;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_CO5;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_CO6;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_C_CY;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_C_XOR;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_D;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_D1;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_D2;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_D3;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_D4;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_D5;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_D6;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_DO5;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_DO6;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_D_CY;
  wire [0:0] CLBLL_L_X54Y105_SLICE_X83Y105_D_XOR;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_A;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_A1;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_A2;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_A3;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_A4;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_A5;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_A6;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_AMUX;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_AO5;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_AO6;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_AX;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_A_CY;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_A_XOR;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_B;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_B1;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_B2;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_B3;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_B4;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_B5;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_B6;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_BMUX;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_BO5;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_BO6;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_BX;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_B_CY;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_B_XOR;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_C;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_C1;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_C2;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_C3;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_C4;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_C5;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_C6;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_CIN;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_CMUX;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_CO5;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_CO6;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_COUT;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_CX;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_C_CY;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_C_XOR;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_D;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_D1;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_D2;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_D3;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_D4;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_D5;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_D6;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_DMUX;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_DO5;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_DO6;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_DX;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_D_CY;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X82Y106_D_XOR;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_A;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_A1;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_A2;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_A3;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_A4;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_A5;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_A6;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_AMUX;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_AO5;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_AO6;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_A_CY;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_A_XOR;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_B;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_B1;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_B2;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_B3;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_B4;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_B5;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_B6;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_BMUX;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_BO5;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_BO6;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_B_CY;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_B_XOR;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_C;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_C1;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_C2;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_C3;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_C4;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_C5;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_C6;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_CMUX;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_CO5;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_CO6;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_C_CY;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_C_XOR;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_D;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_D1;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_D2;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_D3;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_D4;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_D5;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_D6;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_DO5;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_DO6;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_D_CY;
  wire [0:0] CLBLL_L_X54Y106_SLICE_X83Y106_D_XOR;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_A;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_A1;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_A2;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_A3;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_A4;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_A5;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_A6;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_AMUX;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_AO5;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_AO6;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_AX;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_A_CY;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_A_XOR;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_B;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_B1;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_B2;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_B3;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_B4;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_B5;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_B6;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_BMUX;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_BO5;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_BO6;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_BX;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_B_CY;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_B_XOR;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_C;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_C1;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_C2;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_C3;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_C4;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_C5;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_C6;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_CIN;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_CMUX;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_CO5;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_CO6;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_COUT;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_CX;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_C_CY;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_C_XOR;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_D;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_D1;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_D2;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_D3;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_D4;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_D5;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_D6;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_DMUX;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_DO5;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_DO6;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_DX;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_D_CY;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X82Y107_D_XOR;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_A;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_A1;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_A2;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_A3;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_A4;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_A5;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_A6;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_AMUX;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_AO5;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_AO6;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_A_CY;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_A_XOR;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_B;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_B1;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_B2;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_B3;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_B4;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_B5;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_B6;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_BMUX;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_BO5;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_BO6;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_B_CY;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_B_XOR;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_C;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_C1;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_C2;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_C3;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_C4;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_C5;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_C6;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_CO5;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_CO6;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_C_CY;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_C_XOR;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_D;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_D1;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_D2;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_D3;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_D4;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_D5;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_D6;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_DMUX;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_DO5;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_DO6;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_D_CY;
  wire [0:0] CLBLL_L_X54Y107_SLICE_X83Y107_D_XOR;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_A;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_A1;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_A2;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_A3;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_A4;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_A5;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_A6;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_AMUX;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_AO5;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_AO6;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_AX;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_A_CY;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_A_XOR;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_B;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_B1;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_B2;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_B3;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_B4;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_B5;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_B6;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_BO5;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_BO6;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_BX;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_B_CY;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_B_XOR;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_C;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_C1;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_C2;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_C3;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_C4;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_C5;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_C6;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_CIN;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_CO5;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_CO6;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_COUT;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_CX;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_C_CY;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_C_XOR;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_D;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_D1;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_D2;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_D3;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_D4;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_D5;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_D6;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_DO5;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_DO6;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_DX;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_D_CY;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X82Y108_D_XOR;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_A;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_A1;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_A2;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_A3;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_A4;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_A5;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_A6;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_AMUX;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_AO5;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_AO6;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_A_CY;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_A_XOR;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_B;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_B1;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_B2;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_B3;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_B4;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_B5;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_B6;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_BO5;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_BO6;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_B_CY;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_B_XOR;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_C;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_C1;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_C2;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_C3;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_C4;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_C5;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_C6;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_CO5;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_CO6;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_C_CY;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_C_XOR;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_D;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_D1;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_D2;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_D3;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_D4;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_D5;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_D6;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_DO5;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_DO6;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_D_CY;
  wire [0:0] CLBLL_L_X54Y108_SLICE_X83Y108_D_XOR;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_A;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_A1;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_A2;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_A3;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_A4;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_A5;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_A6;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_AO5;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_AQ;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_AX;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_A_CY;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_A_XOR;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_B;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_B1;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_B2;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_B3;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_B4;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_B5;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_B6;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_BO5;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_BO6;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_B_CY;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_B_XOR;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_C;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_C1;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_C2;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_C3;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_C4;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_C5;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_C6;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_CLK;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_CO5;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_CO6;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_C_CY;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_C_XOR;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_D;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_D1;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_D2;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_D3;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_D4;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_D5;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_D6;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_DO5;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_DO6;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_D_CY;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_D_XOR;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X82Y109_SR;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_A;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_A1;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_A2;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_A3;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_A4;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_A5;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_A6;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_AO5;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_AO6;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_A_CY;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_A_XOR;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_B;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_B1;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_B2;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_B3;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_B4;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_B5;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_B6;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_BO5;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_BO6;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_B_CY;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_B_XOR;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_C;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_C1;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_C2;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_C3;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_C4;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_C5;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_C6;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_CO5;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_CO6;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_C_CY;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_C_XOR;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_D;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_D1;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_D2;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_D3;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_D4;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_D5;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_D6;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_DO5;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_DO6;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_D_CY;
  wire [0:0] CLBLL_L_X54Y109_SLICE_X83Y109_D_XOR;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_A;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_A1;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_A2;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_A3;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_A4;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_A5;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_A6;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_AO5;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_AO6;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_A_CY;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_A_XOR;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_B;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_B1;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_B2;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_B3;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_B4;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_B5;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_B6;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_BO5;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_BO6;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_B_CY;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_B_XOR;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_C;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_C1;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_C2;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_C3;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_C4;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_C5;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_C6;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_CO5;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_CO6;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_C_CY;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_C_XOR;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_D;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_D1;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_D2;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_D3;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_D4;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_D5;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_D6;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_DO5;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_DO6;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_D_CY;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X82Y97_D_XOR;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_A;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_A1;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_A2;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_A3;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_A4;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_A5;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_A6;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_AO5;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_AO6;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_A_CY;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_A_XOR;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_B;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_B1;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_B2;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_B3;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_B4;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_B5;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_B6;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_BO5;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_BO6;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_B_CY;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_B_XOR;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_C;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_C1;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_C2;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_C3;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_C4;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_C5;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_C6;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_CO5;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_CO6;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_C_CY;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_C_XOR;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_D;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_D1;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_D2;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_D3;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_D4;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_D5;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_D6;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_DO5;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_DO6;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_D_CY;
  wire [0:0] CLBLL_L_X54Y97_SLICE_X83Y97_D_XOR;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_A;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_A1;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_A2;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_A3;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_A4;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_A5;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_A6;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_AO5;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_AO6;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_A_CY;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_A_XOR;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_B;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_B1;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_B2;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_B3;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_B4;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_B5;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_B6;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_BMUX;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_BO5;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_BO6;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_B_CY;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_B_XOR;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_C;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_C1;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_C2;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_C3;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_C4;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_C5;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_C6;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_CO5;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_CO6;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_C_CY;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_C_XOR;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_D;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_D1;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_D2;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_D3;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_D4;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_D5;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_D6;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_DO5;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_DO6;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_D_CY;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X82Y98_D_XOR;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_A;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_A1;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_A2;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_A3;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_A4;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_A5;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_A6;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_AO5;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_AO6;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_AQ;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_A_CY;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_A_XOR;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_B;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_B1;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_B2;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_B3;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_B4;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_B5;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_B6;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_BO5;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_BO6;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_BQ;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_B_CY;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_B_XOR;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_C;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_C1;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_C2;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_C3;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_C4;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_C5;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_C6;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_CE;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_CLK;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_CMUX;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_CO5;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_CO6;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_C_CY;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_C_XOR;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_D;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_D1;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_D2;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_D3;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_D4;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_D5;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_D6;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_DO5;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_DO6;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_D_CY;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_D_XOR;
  wire [0:0] CLBLL_L_X54Y98_SLICE_X83Y98_SR;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_A;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_A1;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_A2;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_A3;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_A4;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_A5;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_A6;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_AMUX;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_AO5;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_AO6;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_AQ;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_AX;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_A_CY;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_A_XOR;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_B;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_B1;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_B2;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_B3;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_B4;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_B5;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_B6;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_BMUX;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_BO5;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_BO6;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_B_CY;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_B_XOR;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_C;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_C1;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_C2;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_C3;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_C4;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_C5;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_C6;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_CE;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_CLK;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_CO5;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_CO6;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_CQ;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_C_CY;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_C_XOR;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_D;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_D1;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_D2;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_D3;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_D4;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_D5;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_D6;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_DO5;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_DO6;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_D_CY;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_D_XOR;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X82Y99_SR;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_A;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_A1;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_A2;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_A3;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_A4;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_A5;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_A5Q;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_A6;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_AMUX;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_AO5;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_AO6;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_AQ;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_AX;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_A_CY;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_A_XOR;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_B;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_B1;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_B2;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_B3;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_B4;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_B5;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_B6;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_BMUX;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_BO5;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_BO6;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_B_CY;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_B_XOR;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_C;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_C1;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_C2;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_C3;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_C4;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_C5;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_C6;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_CE;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_CLK;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_CO5;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_CO6;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_C_CY;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_C_XOR;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_D;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_D1;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_D2;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_D3;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_D4;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_D5;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_D6;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_DO5;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_DO6;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_D_CY;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_D_XOR;
  wire [0:0] CLBLL_L_X54Y99_SLICE_X83Y99_SR;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_A;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_A1;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_A2;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_A3;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_A4;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_A5;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_A6;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_AMUX;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_AO5;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_AO6;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_AQ;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_A_CY;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_A_XOR;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_B;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_B1;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_B2;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_B3;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_B4;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_B5;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_B6;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_BO5;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_BO6;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_BQ;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_B_CY;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_B_XOR;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_C;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_C1;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_C2;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_C3;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_C4;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_C5;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_C6;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_CE;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_CLK;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_CO5;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_CO6;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_CQ;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_C_CY;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_C_XOR;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_D;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_D1;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_D2;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_D3;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_D4;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_D5;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_D6;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_DO5;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_DO6;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_DQ;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_D_CY;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_D_XOR;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X86Y100_SR;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_A;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_A1;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_A2;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_A3;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_A4;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_A5;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_A6;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_AO5;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_AO6;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_AQ;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_A_CY;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_A_XOR;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_B;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_B1;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_B2;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_B3;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_B4;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_B5;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_B6;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_BO5;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_BO6;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_BQ;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_B_CY;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_B_XOR;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_C;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_C1;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_C2;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_C3;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_C4;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_C5;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_C6;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_CE;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_CLK;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_CO5;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_CO6;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_CQ;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_C_CY;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_C_XOR;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_D;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_D1;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_D2;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_D3;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_D4;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_D5;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_D6;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_DO5;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_DO6;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_D_CY;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_D_XOR;
  wire [0:0] CLBLL_R_X57Y100_SLICE_X87Y100_SR;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_A;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_A1;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_A2;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_A3;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_A4;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_A5;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_A6;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_AMUX;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_AO5;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_AO6;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_AQ;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_A_CY;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_A_XOR;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_B;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_B1;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_B2;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_B3;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_B4;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_B5;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_B6;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_BO5;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_BO6;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_B_CY;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_B_XOR;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_C;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_C1;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_C2;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_C3;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_C4;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_C5;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_C6;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_CE;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_CLK;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_CO5;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_CO6;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_C_CY;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_C_XOR;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_D;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_D1;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_D2;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_D3;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_D4;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_D5;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_D6;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_DO5;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_DO6;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_D_CY;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_D_XOR;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X86Y101_SR;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_A;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_A1;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_A2;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_A3;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_A4;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_A5;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_A6;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_AO5;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_AO6;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_AQ;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_A_CY;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_A_XOR;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_B;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_B1;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_B2;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_B3;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_B4;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_B5;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_B6;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_BMUX;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_BO5;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_BO6;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_B_CY;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_B_XOR;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_C;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_C1;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_C2;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_C3;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_C4;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_C5;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_C6;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_CE;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_CLK;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_CO5;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_CO6;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_CQ;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_C_CY;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_C_XOR;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_D;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_D1;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_D2;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_D3;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_D4;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_D5;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_D6;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_DO5;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_DO6;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_DQ;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_D_CY;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_D_XOR;
  wire [0:0] CLBLL_R_X57Y101_SLICE_X87Y101_SR;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_A;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_A1;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_A2;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_A3;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_A4;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_A5;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_A6;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_AMUX;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_AO5;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_AO6;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_AQ;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_AX;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_A_CY;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_A_XOR;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_B;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_B1;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_B2;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_B3;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_B4;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_B5;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_B6;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_BO5;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_BO6;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_BQ;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_B_CY;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_B_XOR;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_C;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_C1;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_C2;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_C3;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_C4;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_C5;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_C6;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_CE;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_CLK;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_CMUX;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_CO5;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_CO6;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_C_CY;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_C_XOR;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_D;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_D1;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_D2;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_D3;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_D4;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_D5;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_D6;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_DO5;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_DO6;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_D_CY;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_D_XOR;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X86Y102_SR;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_A;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_A1;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_A2;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_A3;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_A4;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_A5;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_A6;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_AO5;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_AO6;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_A_CY;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_A_XOR;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_B;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_B1;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_B2;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_B3;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_B4;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_B5;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_B6;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_BO5;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_BO6;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_B_CY;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_B_XOR;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_C;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_C1;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_C2;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_C3;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_C4;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_C5;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_C6;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_CO5;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_CO6;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_C_CY;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_C_XOR;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_D;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_D1;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_D2;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_D3;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_D4;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_D5;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_D6;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_DO5;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_DO6;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_D_CY;
  wire [0:0] CLBLL_R_X57Y102_SLICE_X87Y102_D_XOR;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_A;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_A1;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_A2;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_A3;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_A4;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_A5;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_A5Q;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_A6;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_AMUX;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_AO5;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_AO6;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_AQ;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_A_CY;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_A_XOR;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_B;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_B1;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_B2;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_B3;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_B4;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_B5;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_B6;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_BO5;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_BO6;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_B_CY;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_B_XOR;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_C;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_C1;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_C2;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_C3;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_C4;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_C5;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_C6;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_CLK;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_CO5;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_CO6;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_C_CY;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_C_XOR;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_D;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_D1;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_D2;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_D3;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_D4;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_D5;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_D6;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_DO5;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_DO6;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_D_CY;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_D_XOR;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X86Y103_SR;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_A;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_A1;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_A2;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_A3;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_A4;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_A5;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_A6;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_AO5;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_AO6;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_AQ;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_A_CY;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_A_XOR;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_B;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_B1;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_B2;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_B3;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_B4;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_B5;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_B6;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_BO5;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_BO6;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_B_CY;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_B_XOR;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_C;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_C1;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_C2;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_C3;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_C4;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_C5;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_C6;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_CE;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_CLK;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_CO5;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_CO6;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_C_CY;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_C_XOR;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_D;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_D1;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_D2;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_D3;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_D4;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_D5;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_D6;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_DO5;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_DO6;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_D_CY;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_D_XOR;
  wire [0:0] CLBLL_R_X57Y103_SLICE_X87Y103_SR;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_A;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_A1;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_A2;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_A3;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_A4;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_A5;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_A6;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_AO5;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_AO6;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_AQ;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_A_CY;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_A_XOR;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_B;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_B1;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_B2;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_B3;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_B4;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_B5;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_B6;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_BO5;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_BO6;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_BQ;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_B_CY;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_B_XOR;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_C;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_C1;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_C2;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_C3;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_C4;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_C5;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_C6;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_CE;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_CLK;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_CO5;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_CO6;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_CQ;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_C_CY;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_C_XOR;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_D;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_D1;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_D2;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_D3;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_D4;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_D5;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_D6;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_DO5;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_DO6;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_D_CY;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_D_XOR;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X86Y104_SR;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_A;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_A1;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_A2;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_A3;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_A4;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_A5;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_A6;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_AO5;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_AO6;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_AQ;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_A_CY;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_A_XOR;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_B;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_B1;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_B2;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_B3;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_B4;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_B5;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_B6;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_BO5;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_BO6;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_BQ;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_B_CY;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_B_XOR;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_C;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_C1;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_C2;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_C3;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_C4;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_C5;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_C6;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_CE;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_CLK;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_CO5;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_CO6;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_CQ;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_C_CY;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_C_XOR;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_D;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_D1;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_D2;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_D3;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_D4;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_D5;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_D6;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_DO5;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_DO6;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_D_CY;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_D_XOR;
  wire [0:0] CLBLL_R_X57Y104_SLICE_X87Y104_SR;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_A;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_A1;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_A2;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_A3;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_A4;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_A5;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_A6;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_AO5;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_AO6;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_AQ;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_A_CY;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_A_XOR;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_B;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_B1;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_B2;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_B3;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_B4;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_B5;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_B6;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_BO5;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_BO6;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_BQ;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_B_CY;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_B_XOR;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_C;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_C1;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_C2;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_C3;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_C4;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_C5;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_C6;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_CE;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_CLK;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_CO5;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_CO6;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_C_CY;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_C_XOR;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_D;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_D1;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_D2;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_D3;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_D4;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_D5;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_D6;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_DO5;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_DO6;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_D_CY;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_D_XOR;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X86Y105_SR;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_A;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_A1;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_A2;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_A3;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_A4;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_A5;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_A6;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_AMUX;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_AO5;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_AO6;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_AX;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_A_CY;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_A_XOR;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_B;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_B1;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_B2;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_B3;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_B4;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_B5;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_B6;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_BMUX;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_BO5;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_BO6;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_BX;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_B_CY;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_B_XOR;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_C;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_C1;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_C2;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_C3;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_C4;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_C5;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_C6;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_CMUX;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_CO5;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_CO6;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_COUT;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_CX;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_C_CY;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_C_XOR;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_D;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_D1;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_D2;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_D3;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_D4;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_D5;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_D6;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_DMUX;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_DO5;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_DO6;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_DX;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_D_CY;
  wire [0:0] CLBLL_R_X57Y105_SLICE_X87Y105_D_XOR;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_A;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_A1;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_A2;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_A3;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_A4;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_A5;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_A6;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_AMUX;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_AO5;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_AO6;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_AX;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_A_CY;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_A_XOR;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_B;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_B1;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_B2;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_B3;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_B4;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_B5;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_B6;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_BMUX;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_BO5;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_BO6;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_BX;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_B_CY;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_B_XOR;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_C;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_C1;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_C2;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_C3;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_C4;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_C5;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_C6;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_CMUX;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_CO5;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_CO6;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_COUT;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_CX;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_C_CY;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_C_XOR;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_D;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_D1;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_D2;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_D3;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_D4;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_D5;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_D6;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_DMUX;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_DO5;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_DO6;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_DX;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_D_CY;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X86Y106_D_XOR;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_A;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_A1;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_A2;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_A3;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_A4;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_A5;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_A6;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_AMUX;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_AO5;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_AO6;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_AQ;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_AX;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_A_CY;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_A_XOR;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_B;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_B1;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_B2;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_B3;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_B4;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_B5;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_B6;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_BMUX;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_BO5;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_BO6;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_BX;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_B_CY;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_B_XOR;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_C;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_C1;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_C2;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_C3;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_C4;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_C5;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_C6;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_CE;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_CIN;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_CLK;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_CMUX;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_CO5;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_CO6;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_COUT;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_CX;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_C_CY;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_C_XOR;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_D;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_D1;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_D2;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_D3;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_D4;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_D5;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_D6;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_DMUX;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_DO5;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_DO6;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_DX;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_D_CY;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_D_XOR;
  wire [0:0] CLBLL_R_X57Y106_SLICE_X87Y106_SR;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_A;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_A1;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_A2;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_A3;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_A4;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_A5;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_A6;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_AMUX;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_AO5;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_AO6;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_AX;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_A_CY;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_A_XOR;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_B;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_B1;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_B2;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_B3;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_B4;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_B5;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_B6;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_BMUX;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_BO5;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_BO6;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_BX;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_B_CY;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_B_XOR;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_C;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_C1;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_C2;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_C3;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_C4;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_C5;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_C6;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_CIN;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_CMUX;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_CO5;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_CO6;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_COUT;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_CX;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_C_CY;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_C_XOR;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_D;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_D1;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_D2;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_D3;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_D4;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_D5;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_D6;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_DMUX;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_DO5;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_DO6;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_DX;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_D_CY;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X86Y107_D_XOR;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_A;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_A1;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_A2;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_A3;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_A4;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_A5;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_A6;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_AMUX;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_AO5;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_AO6;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_AX;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_A_CY;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_A_XOR;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_B;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_B1;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_B2;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_B3;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_B4;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_B5;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_B6;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_BMUX;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_BO5;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_BO6;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_BX;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_B_CY;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_B_XOR;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_C;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_C1;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_C2;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_C3;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_C4;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_C5;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_C6;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_CIN;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_CMUX;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_CO5;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_CO6;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_COUT;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_CX;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_C_CY;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_C_XOR;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_D;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_D1;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_D2;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_D3;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_D4;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_D5;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_D6;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_DO5;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_DO6;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_DX;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_D_CY;
  wire [0:0] CLBLL_R_X57Y107_SLICE_X87Y107_D_XOR;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_A;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_A1;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_A2;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_A3;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_A4;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_A5;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_A6;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_AMUX;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_AO5;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_AO6;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_AX;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_A_CY;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_A_XOR;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_B;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_B1;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_B2;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_B3;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_B4;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_B5;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_B6;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_BMUX;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_BO5;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_BO6;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_BX;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_B_CY;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_B_XOR;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_C;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_C1;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_C2;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_C3;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_C4;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_C5;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_C6;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_CIN;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_CMUX;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_CO5;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_CO6;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_COUT;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_CX;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_C_CY;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_C_XOR;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_D;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_D1;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_D2;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_D3;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_D4;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_D5;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_D6;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_DO5;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_DO6;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_DX;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_D_CY;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X86Y108_D_XOR;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_A;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_A1;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_A2;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_A3;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_A4;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_A5;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_A6;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_AO5;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_AO6;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_AQ;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_A_CY;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_A_XOR;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_B;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_B1;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_B2;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_B3;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_B4;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_B5;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_B6;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_BO5;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_BO6;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_BQ;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_B_CY;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_B_XOR;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_C;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_C1;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_C2;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_C3;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_C4;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_C5;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_C6;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_CE;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_CLK;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_CO5;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_CO6;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_C_CY;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_C_XOR;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_D;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_D1;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_D2;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_D3;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_D4;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_D5;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_D6;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_DO5;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_DO6;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_D_CY;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_D_XOR;
  wire [0:0] CLBLL_R_X57Y108_SLICE_X87Y108_SR;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_A;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_A1;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_A2;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_A3;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_A4;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_A5;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_A6;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_AO5;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_AO6;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_AQ;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_A_CY;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_A_XOR;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_B;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_B1;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_B2;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_B3;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_B4;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_B5;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_B6;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_BO5;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_BO6;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_BQ;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_B_CY;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_B_XOR;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_C;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_C1;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_C2;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_C3;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_C4;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_C5;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_C6;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_CE;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_CLK;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_CO5;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_CO6;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_CQ;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_C_CY;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_C_XOR;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_D;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_D1;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_D2;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_D3;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_D4;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_D5;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_D6;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_DO5;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_DO6;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_D_CY;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_D_XOR;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X86Y109_SR;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_A;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_A1;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_A2;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_A3;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_A4;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_A5;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_A6;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_AMUX;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_AO5;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_AO6;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_AX;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_A_CY;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_A_XOR;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_B;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_B1;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_B2;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_B3;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_B4;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_B5;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_B6;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_BMUX;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_BO5;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_BO6;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_BX;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_B_CY;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_B_XOR;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_C;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_C1;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_C2;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_C3;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_C4;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_C5;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_C6;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_CMUX;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_CO5;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_CO6;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_COUT;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_CX;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_C_CY;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_C_XOR;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_D;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_D1;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_D2;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_D3;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_D4;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_D5;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_D6;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_DMUX;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_DO5;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_DO6;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_DX;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_D_CY;
  wire [0:0] CLBLL_R_X57Y109_SLICE_X87Y109_D_XOR;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_A;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_A1;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_A2;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_A3;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_A4;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_A5;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_A6;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_AO5;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_AO6;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_A_CY;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_A_XOR;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_B;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_B1;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_B2;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_B3;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_B4;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_B5;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_B6;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_BO5;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_BO6;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_B_CY;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_B_XOR;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_C;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_C1;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_C2;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_C3;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_C4;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_C5;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_C6;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_CO5;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_CO6;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_C_CY;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_C_XOR;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_D;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_D1;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_D2;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_D3;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_D4;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_D5;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_D6;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_DO5;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_DO6;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_D_CY;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X86Y110_D_XOR;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_A;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_A1;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_A2;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_A3;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_A4;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_A5;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_A6;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_AMUX;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_AO5;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_AO6;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_AX;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_A_CY;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_A_XOR;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_B;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_B1;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_B2;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_B3;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_B4;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_B5;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_B6;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_BMUX;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_BO5;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_BO6;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_BX;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_B_CY;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_B_XOR;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_C;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_C1;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_C2;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_C3;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_C4;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_C5;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_C6;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_CIN;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_CMUX;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_CO5;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_CO6;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_COUT;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_CX;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_C_CY;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_C_XOR;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_D;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_D1;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_D2;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_D3;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_D4;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_D5;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_D6;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_DMUX;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_DO5;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_DO6;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_DX;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_D_CY;
  wire [0:0] CLBLL_R_X57Y110_SLICE_X87Y110_D_XOR;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_A;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_A1;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_A2;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_A3;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_A4;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_A5;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_A6;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_AO5;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_AO6;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_A_CY;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_A_XOR;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_B;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_B1;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_B2;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_B3;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_B4;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_B5;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_B6;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_BO5;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_BO6;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_B_CY;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_B_XOR;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_C;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_C1;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_C2;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_C3;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_C4;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_C5;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_C6;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_CO5;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_CO6;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_C_CY;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_C_XOR;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_D;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_D1;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_D2;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_D3;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_D4;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_D5;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_D6;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_DO5;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_DO6;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_D_CY;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X86Y111_D_XOR;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_A;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_A1;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_A2;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_A3;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_A4;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_A5;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_A6;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_AMUX;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_AO5;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_AO6;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_AX;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_A_CY;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_A_XOR;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_B;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_B1;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_B2;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_B3;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_B4;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_B5;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_B6;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_BMUX;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_BO5;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_BO6;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_BX;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_B_CY;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_B_XOR;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_C;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_C1;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_C2;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_C3;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_C4;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_C5;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_C6;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_CIN;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_CMUX;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_CO5;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_CO6;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_COUT;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_CX;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_C_CY;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_C_XOR;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_D;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_D1;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_D2;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_D3;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_D4;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_D5;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_D6;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_DMUX;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_DO5;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_DO6;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_DX;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_D_CY;
  wire [0:0] CLBLL_R_X57Y111_SLICE_X87Y111_D_XOR;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_A;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_A1;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_A2;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_A3;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_A4;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_A5;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_A6;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_AO5;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_AO6;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_AQ;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_A_CY;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_A_XOR;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_B;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_B1;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_B2;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_B3;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_B4;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_B5;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_B6;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_BMUX;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_BO5;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_BO6;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_B_CY;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_B_XOR;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_C;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_C1;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_C2;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_C3;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_C4;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_C5;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_C6;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_CLK;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_CO5;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_CO6;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_C_CY;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_C_XOR;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_D;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_D1;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_D2;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_D3;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_D4;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_D5;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_D6;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_DO5;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_DO6;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_D_CY;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_D_XOR;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X86Y97_SR;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_A;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_A1;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_A2;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_A3;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_A4;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_A5;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_A6;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_AO5;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_AO6;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_AQ;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_AX;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_A_CY;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_A_XOR;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_B;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_B1;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_B2;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_B3;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_B4;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_B5;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_B6;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_BO5;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_BO6;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_B_CY;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_B_XOR;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_C;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_C1;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_C2;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_C3;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_C4;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_C5;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_C6;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_CE;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_CLK;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_CO5;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_CO6;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_C_CY;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_C_XOR;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_D;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_D1;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_D2;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_D3;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_D4;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_D5;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_D6;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_DO5;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_DO6;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_D_CY;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_D_XOR;
  wire [0:0] CLBLL_R_X57Y97_SLICE_X87Y97_SR;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_A;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_A1;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_A2;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_A3;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_A4;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_A5;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_A6;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_AO5;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_AO6;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_A_CY;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_A_XOR;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_B;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_B1;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_B2;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_B3;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_B4;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_B5;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_B6;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_BO5;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_BO6;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_B_CY;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_B_XOR;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_C;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_C1;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_C2;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_C3;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_C4;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_C5;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_C6;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_CO5;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_CO6;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_C_CY;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_C_XOR;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_D;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_D1;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_D2;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_D3;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_D4;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_D5;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_D6;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_DO5;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_DO6;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_D_CY;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X86Y98_D_XOR;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_A;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_A1;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_A2;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_A3;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_A4;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_A5;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_A6;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_AO5;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_AO6;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_AQ;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_AX;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_A_CY;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_A_XOR;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_B;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_B1;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_B2;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_B3;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_B4;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_B5;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_B6;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_BO5;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_BO6;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_BQ;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_BX;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_B_CY;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_B_XOR;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_C;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_C1;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_C2;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_C3;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_C4;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_C5;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_C6;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_CE;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_CLK;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_CO5;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_CO6;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_CQ;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_CX;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_C_CY;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_C_XOR;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_D;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_D1;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_D2;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_D3;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_D4;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_D5;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_D6;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_DO5;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_DO6;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_DQ;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_DX;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_D_CY;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_D_XOR;
  wire [0:0] CLBLL_R_X57Y98_SLICE_X87Y98_SR;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_A;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_A1;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_A2;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_A3;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_A4;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_A5;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_A6;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_AO5;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_AO6;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_AQ;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_A_CY;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_A_XOR;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_B;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_B1;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_B2;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_B3;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_B4;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_B5;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_B6;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_BO5;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_BO6;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_BQ;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_B_CY;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_B_XOR;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_C;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_C1;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_C2;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_C3;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_C4;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_C5;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_C6;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_CE;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_CLK;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_CO5;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_CO6;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_C_CY;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_C_XOR;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_D;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_D1;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_D2;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_D3;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_D4;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_D5;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_D6;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_DO5;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_DO6;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_D_CY;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_D_XOR;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X86Y99_SR;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_A;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_A1;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_A2;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_A3;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_A4;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_A5;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_A6;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_AO5;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_AO6;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_AQ;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_A_CY;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_A_XOR;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_B;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_B1;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_B2;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_B3;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_B4;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_B5;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_B6;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_BO5;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_BO6;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_B_CY;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_B_XOR;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_C;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_C1;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_C2;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_C3;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_C4;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_C5;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_C6;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_CLK;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_CO5;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_CO6;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_C_CY;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_C_XOR;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_D;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_D1;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_D2;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_D3;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_D4;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_D5;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_D6;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_DO5;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_DO6;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_D_CY;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_D_XOR;
  wire [0:0] CLBLL_R_X57Y99_SLICE_X87Y99_SR;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_A;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_A1;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_A2;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_A3;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_A4;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_A5;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_A6;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_AO5;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_AO6;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_AQ;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_AX;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_A_CY;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_A_XOR;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_B;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_B1;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_B2;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_B3;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_B4;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_B5;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_B6;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_BO5;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_BO6;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_BQ;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_BX;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_B_CY;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_B_XOR;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_C;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_C1;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_C2;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_C3;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_C4;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_C5;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_C6;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_CLK;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_CO5;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_CO6;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_C_CY;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_C_XOR;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_D;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_D1;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_D2;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_D3;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_D4;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_D5;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_D6;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_DO5;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_DO6;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_D_CY;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_D_XOR;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X46Y119_SR;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_A;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_A1;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_A2;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_A3;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_A4;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_A5;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_A6;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_AO5;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_AO6;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_A_CY;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_A_XOR;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_B;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_B1;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_B2;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_B3;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_B4;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_B5;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_B6;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_BO5;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_BO6;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_B_CY;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_B_XOR;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_C;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_C1;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_C2;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_C3;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_C4;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_C5;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_C6;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_CO5;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_CO6;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_C_CY;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_C_XOR;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_D;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_D1;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_D2;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_D3;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_D4;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_D5;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_D6;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_DO5;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_DO6;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_D_CY;
  wire [0:0] CLBLM_L_X32Y119_SLICE_X47Y119_D_XOR;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_A;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_A1;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_A2;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_A3;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_A4;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_A5;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_A6;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_AO5;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_AO6;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_AQ;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_A_CY;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_A_XOR;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_B;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_B1;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_B2;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_B3;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_B4;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_B5;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_B6;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_BO5;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_BO6;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_B_CY;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_B_XOR;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_C;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_C1;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_C2;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_C3;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_C4;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_C5;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_C6;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_CE;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_CLK;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_CO5;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_CO6;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_C_CY;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_C_XOR;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_D;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_D1;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_D2;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_D3;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_D4;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_D5;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_D6;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_DO5;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_DO6;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_D_CY;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_D_XOR;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X76Y104_SR;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_A;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_A1;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_A2;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_A3;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_A4;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_A5;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_A6;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_AO5;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_AO6;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_A_CY;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_A_XOR;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_B;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_B1;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_B2;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_B3;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_B4;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_B5;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_B6;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_BO5;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_BO6;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_B_CY;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_B_XOR;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_C;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_C1;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_C2;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_C3;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_C4;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_C5;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_C6;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_CO5;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_CO6;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_C_CY;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_C_XOR;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_D;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_D1;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_D2;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_D3;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_D4;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_D5;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_D6;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_DO5;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_DO6;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_D_CY;
  wire [0:0] CLBLM_L_X50Y104_SLICE_X77Y104_D_XOR;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_A;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_A1;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_A2;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_A3;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_A4;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_A5;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_A6;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_AO5;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_AO6;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_AQ;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_A_CY;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_A_XOR;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_B;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_B1;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_B2;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_B3;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_B4;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_B5;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_B6;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_BMUX;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_BO5;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_BO6;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_B_CY;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_B_XOR;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_C;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_C1;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_C2;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_C3;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_C4;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_C5;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_C6;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_CE;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_CLK;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_CMUX;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_CO5;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_CO6;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_C_CY;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_C_XOR;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_D;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_D1;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_D2;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_D3;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_D4;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_D5;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_D6;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_DO5;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_DO6;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_D_CY;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_D_XOR;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X76Y105_SR;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_A;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_A1;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_A2;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_A3;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_A4;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_A5;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_A6;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_AO5;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_AO6;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_AQ;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_AX;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_A_CY;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_A_XOR;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_B;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_B1;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_B2;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_B3;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_B4;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_B5;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_B6;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_BO5;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_BO6;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_B_CY;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_B_XOR;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_C;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_C1;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_C2;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_C3;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_C4;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_C5;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_C6;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_CE;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_CLK;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_CO5;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_CO6;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_C_CY;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_C_XOR;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_D;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_D1;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_D2;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_D3;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_D4;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_D5;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_D6;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_DO5;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_DO6;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_D_CY;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_D_XOR;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_F7AMUX_O;
  wire [0:0] CLBLM_L_X50Y105_SLICE_X77Y105_SR;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_A;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_A1;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_A2;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_A3;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_A4;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_A5;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_A6;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_AO5;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_AO6;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_AQ;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_A_CY;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_A_XOR;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_B;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_B1;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_B2;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_B3;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_B4;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_B5;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_B6;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_BMUX;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_BO5;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_BO6;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_B_CY;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_B_XOR;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_C;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_C1;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_C2;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_C3;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_C4;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_C5;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_C6;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_CE;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_CLK;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_CO5;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_CO6;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_CQ;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_C_CY;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_C_XOR;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_D;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_D1;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_D2;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_D3;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_D4;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_D5;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_D6;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_DO5;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_DO6;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_D_CY;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_D_XOR;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X76Y106_SR;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_A;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_A1;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_A2;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_A3;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_A4;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_A5;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_A6;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_AMUX;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_AO5;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_AO6;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_A_CY;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_A_XOR;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_B;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_B1;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_B2;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_B3;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_B4;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_B5;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_B6;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_BMUX;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_BO5;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_BO6;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_B_CY;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_B_XOR;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_C;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_C1;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_C2;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_C3;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_C4;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_C5;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_C6;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_CO5;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_CO6;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_C_CY;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_C_XOR;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_D;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_D1;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_D2;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_D3;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_D4;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_D5;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_D6;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_DO5;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_DO6;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_D_CY;
  wire [0:0] CLBLM_L_X50Y106_SLICE_X77Y106_D_XOR;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_A;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_A1;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_A2;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_A3;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_A4;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_A5;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_A6;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_AMUX;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_AO5;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_AO6;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_A_CY;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_A_XOR;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_B;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_B1;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_B2;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_B3;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_B4;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_B5;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_B6;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_BO5;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_BO6;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_BQ;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_B_CY;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_B_XOR;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_C;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_C1;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_C2;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_C3;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_C4;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_C5;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_C6;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_CE;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_CLK;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_CO5;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_CO6;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_C_CY;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_C_XOR;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_D;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_D1;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_D2;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_D3;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_D4;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_D5;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_D6;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_DO5;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_DO6;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_D_CY;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_D_XOR;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X76Y107_SR;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_A;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_A1;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_A2;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_A3;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_A4;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_A5;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_A6;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_AO5;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_AO6;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_AQ;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_A_CY;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_A_XOR;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_B;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_B1;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_B2;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_B3;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_B4;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_B5;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_B6;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_BO5;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_BO6;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_B_CY;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_B_XOR;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_C;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_C1;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_C2;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_C3;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_C4;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_C5;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_C6;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_CE;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_CLK;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_CO5;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_CO6;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_C_CY;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_C_XOR;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_D;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_D1;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_D2;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_D3;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_D4;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_D5;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_D6;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_DO5;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_DO6;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_D_CY;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_D_XOR;
  wire [0:0] CLBLM_L_X50Y107_SLICE_X77Y107_SR;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_A;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_A1;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_A2;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_A3;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_A4;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_A5;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_A6;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_AMUX;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_AO5;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_AO6;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_AX;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_A_CY;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_A_XOR;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_B;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_B1;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_B2;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_B3;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_B4;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_B5;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_B6;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_BMUX;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_BO5;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_BO6;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_BX;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_B_CY;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_B_XOR;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_C;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_C1;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_C2;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_C3;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_C4;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_C5;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_C6;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_CMUX;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_CO5;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_CO6;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_COUT;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_CX;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_C_CY;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_C_XOR;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_D;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_D1;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_D2;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_D3;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_D4;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_D5;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_D6;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_DMUX;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_DO5;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_DO6;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_DX;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_D_CY;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X76Y108_D_XOR;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_A;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_A1;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_A2;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_A3;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_A4;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_A5;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_A6;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_AMUX;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_AO5;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_AO6;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_AX;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_A_CY;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_A_XOR;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_B;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_B1;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_B2;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_B3;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_B4;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_B5;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_B6;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_BMUX;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_BO5;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_BO6;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_B_CY;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_B_XOR;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_C;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_C1;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_C2;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_C3;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_C4;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_C5;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_C6;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_CMUX;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_CO5;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_CO6;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_COUT;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_C_CY;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_C_XOR;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_D;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_D1;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_D2;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_D3;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_D4;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_D5;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_D6;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_DMUX;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_DO5;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_DO6;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_D_CY;
  wire [0:0] CLBLM_L_X50Y108_SLICE_X77Y108_D_XOR;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_A;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_A1;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_A2;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_A3;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_A4;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_A5;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_A6;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_AMUX;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_AO5;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_AO6;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_AX;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_A_CY;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_A_XOR;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_B;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_B1;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_B2;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_B3;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_B4;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_B5;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_B6;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_BMUX;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_BO5;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_BO6;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_BX;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_B_CY;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_B_XOR;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_C;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_C1;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_C2;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_C3;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_C4;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_C5;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_C6;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_CIN;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_CMUX;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_CO5;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_CO6;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_COUT;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_CX;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_C_CY;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_C_XOR;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_D;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_D1;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_D2;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_D3;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_D4;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_D5;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_D6;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_DMUX;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_DO5;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_DO6;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_DX;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_D_CY;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X76Y109_D_XOR;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_A;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_A1;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_A2;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_A3;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_A4;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_A5;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_A6;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_AMUX;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_AO5;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_AO6;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_A_CY;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_A_XOR;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_B;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_B1;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_B2;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_B3;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_B4;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_B5;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_B6;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_BMUX;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_BO5;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_BO6;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_B_CY;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_B_XOR;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_C;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_C1;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_C2;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_C3;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_C4;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_C5;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_C6;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_CIN;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_CMUX;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_CO5;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_CO6;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_COUT;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_C_CY;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_C_XOR;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_D;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_D1;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_D2;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_D3;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_D4;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_D5;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_D6;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_DMUX;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_DO5;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_DO6;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_D_CY;
  wire [0:0] CLBLM_L_X50Y109_SLICE_X77Y109_D_XOR;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_A;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_A1;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_A2;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_A3;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_A4;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_A5;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_A6;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_AMUX;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_AO5;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_AO6;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_AX;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_A_CY;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_A_XOR;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_B;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_B1;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_B2;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_B3;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_B4;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_B5;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_B6;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_BO5;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_BO6;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_BX;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_B_CY;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_B_XOR;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_C;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_C1;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_C2;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_C3;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_C4;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_C5;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_C6;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_CIN;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_CO5;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_CO6;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_COUT;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_CX;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_C_CY;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_C_XOR;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_D;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_D1;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_D2;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_D3;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_D4;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_D5;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_D6;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_DO5;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_DO6;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_DX;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_D_CY;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X76Y110_D_XOR;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_A;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_A1;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_A2;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_A3;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_A4;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_A5;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_A6;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_AMUX;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_AO5;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_AO6;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_AX;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_A_CY;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_A_XOR;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_B;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_B1;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_B2;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_B3;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_B4;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_B5;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_B6;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_BO5;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_BO6;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_BX;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_B_CY;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_B_XOR;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_C;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_C1;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_C2;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_C3;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_C4;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_C5;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_C6;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_CIN;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_CO5;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_CO6;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_COUT;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_CX;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_C_CY;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_C_XOR;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_D;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_D1;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_D2;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_D3;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_D4;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_D5;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_D6;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_DO5;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_DO6;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_DX;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_D_CY;
  wire [0:0] CLBLM_L_X50Y110_SLICE_X77Y110_D_XOR;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_A;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_A1;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_A2;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_A3;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_A4;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_A5;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_A6;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_AO5;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_AO6;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_A_CY;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_A_XOR;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_B;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_B1;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_B2;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_B3;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_B4;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_B5;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_B6;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_BO5;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_BO6;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_B_CY;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_B_XOR;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_C;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_C1;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_C2;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_C3;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_C4;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_C5;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_C6;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_CMUX;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_CO5;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_CO6;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_C_CY;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_C_XOR;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_D;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_D1;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_D2;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_D3;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_D4;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_D5;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_D6;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_DO5;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_DO6;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_D_CY;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X76Y111_D_XOR;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_A;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_A1;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_A2;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_A3;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_A4;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_A5;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_A6;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_AO5;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_AO6;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_A_CY;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_A_XOR;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_B;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_B1;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_B2;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_B3;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_B4;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_B5;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_B6;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_BO5;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_BO6;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_B_CY;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_B_XOR;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_C;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_C1;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_C2;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_C3;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_C4;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_C5;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_C6;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_CO5;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_CO6;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_C_CY;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_C_XOR;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_D;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_D1;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_D2;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_D3;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_D4;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_D5;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_D6;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_DO5;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_DO6;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_D_CY;
  wire [0:0] CLBLM_L_X50Y111_SLICE_X77Y111_D_XOR;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_A;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_A1;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_A2;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_A3;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_A4;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_A5;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_A6;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_AO5;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_AO6;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_AQ;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_A_CY;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_A_XOR;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_B;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_B1;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_B2;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_B3;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_B4;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_B5;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_B6;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_BO5;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_BO6;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_BQ;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_BX;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_B_CY;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_B_XOR;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_C;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_C1;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_C2;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_C3;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_C4;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_C5;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_C6;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_CE;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_CLK;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_CO5;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_CO6;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_COUT;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_CQ;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_CX;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_C_CY;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_C_XOR;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_D;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_D1;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_D2;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_D3;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_D4;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_D5;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_D6;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_DO5;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_DO6;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_DQ;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_DX;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_D_CY;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_D_XOR;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X84Y100_SR;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_A;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_A1;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_A2;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_A3;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_A4;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_A5;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_A6;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_AMUX;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_AO5;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_AO6;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_AQ;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_AX;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_A_CY;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_A_XOR;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_B;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_B1;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_B2;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_B3;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_B4;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_B5;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_B6;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_BMUX;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_BO5;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_BO6;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_BQ;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_BX;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_B_CY;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_B_XOR;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_C;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_C1;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_C2;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_C3;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_C4;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_C5;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_C6;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_CE;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_CLK;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_CO5;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_CO6;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_CQ;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_CX;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_C_CY;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_C_XOR;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_D;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_D1;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_D2;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_D3;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_D4;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_D5;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_D6;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_DO5;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_DO6;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_DQ;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_DX;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_D_CY;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_D_XOR;
  wire [0:0] CLBLM_L_X56Y100_SLICE_X85Y100_SR;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_A;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_A1;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_A2;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_A3;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_A4;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_A5;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_A6;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_AO5;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_AO6;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_AQ;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_AX;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_A_CY;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_A_XOR;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_B;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_B1;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_B2;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_B3;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_B4;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_B5;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_B6;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_BO5;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_BO6;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_BQ;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_BX;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_B_CY;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_B_XOR;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_C;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_C1;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_C2;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_C3;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_C4;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_C5;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_C6;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_CE;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_CIN;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_CLK;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_CO5;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_CO6;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_COUT;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_CQ;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_CX;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_C_CY;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_C_XOR;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_D;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_D1;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_D2;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_D3;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_D4;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_D5;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_D6;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_DO5;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_DO6;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_DQ;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_DX;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_D_CY;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_D_XOR;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X84Y101_SR;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_A;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_A1;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_A2;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_A3;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_A4;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_A5;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_A6;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_AO5;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_AO6;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_AQ;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_A_CY;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_A_XOR;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_B;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_B1;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_B2;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_B3;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_B4;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_B5;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_B6;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_BO5;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_BO6;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_BQ;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_B_CY;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_B_XOR;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_C;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_C1;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_C2;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_C3;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_C4;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_C5;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_C6;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_CE;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_CLK;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_CO5;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_CO6;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_CQ;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_C_CY;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_C_XOR;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_D;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_D1;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_D2;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_D3;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_D4;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_D5;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_D6;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_DO5;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_DO6;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_DQ;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_D_CY;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_D_XOR;
  wire [0:0] CLBLM_L_X56Y101_SLICE_X85Y101_SR;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_A;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_A1;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_A2;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_A3;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_A4;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_A5;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_A6;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_AO5;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_AO6;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_AQ;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_AX;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_A_CY;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_A_XOR;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_B;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_B1;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_B2;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_B3;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_B4;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_B5;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_B6;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_BO5;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_BO6;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_BQ;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_BX;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_B_CY;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_B_XOR;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_C;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_C1;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_C2;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_C3;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_C4;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_C5;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_C6;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_CE;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_CIN;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_CLK;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_CO5;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_CO6;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_COUT;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_CQ;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_CX;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_C_CY;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_C_XOR;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_D;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_D1;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_D2;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_D3;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_D4;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_D5;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_D6;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_DO5;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_DO6;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_DQ;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_DX;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_D_CY;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_D_XOR;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X84Y102_SR;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_A;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_A1;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_A2;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_A3;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_A4;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_A5;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_A5Q;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_A6;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_AMUX;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_AO5;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_AO6;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_AQ;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_A_CY;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_A_XOR;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_B;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_B1;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_B2;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_B3;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_B4;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_B5;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_B6;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_BO5;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_BO6;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_B_CY;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_B_XOR;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_C;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_C1;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_C2;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_C3;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_C4;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_C5;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_C6;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_CLK;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_CO5;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_CO6;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_C_CY;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_C_XOR;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_D;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_D1;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_D2;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_D3;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_D4;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_D5;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_D6;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_DO5;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_DO6;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_D_CY;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_D_XOR;
  wire [0:0] CLBLM_L_X56Y102_SLICE_X85Y102_SR;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_A;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_A1;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_A2;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_A3;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_A4;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_A5;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_A6;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_AO5;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_AO6;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_AQ;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_AX;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_A_CY;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_A_XOR;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_B;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_B1;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_B2;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_B3;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_B4;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_B5;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_B6;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_BO5;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_BO6;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_BQ;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_BX;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_B_CY;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_B_XOR;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_C;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_C1;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_C2;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_C3;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_C4;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_C5;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_C6;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_CE;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_CIN;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_CLK;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_CO5;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_CO6;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_COUT;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_CQ;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_CX;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_C_CY;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_C_XOR;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_D;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_D1;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_D2;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_D3;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_D4;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_D5;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_D6;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_DO5;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_DO6;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_DQ;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_DX;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_D_CY;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_D_XOR;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X84Y103_SR;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_A;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_A1;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_A2;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_A3;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_A4;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_A5;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_A6;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_AO5;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_AO6;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_AQ;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_A_CY;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_A_XOR;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_B;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_B1;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_B2;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_B3;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_B4;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_B5;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_B6;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_BO5;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_BO6;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_BQ;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_B_CY;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_B_XOR;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_C;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_C1;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_C2;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_C3;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_C4;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_C5;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_C6;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_CE;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_CLK;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_CO5;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_CO6;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_C_CY;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_C_XOR;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_D;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_D1;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_D2;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_D3;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_D4;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_D5;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_D6;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_DO5;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_DO6;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_D_CY;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_D_XOR;
  wire [0:0] CLBLM_L_X56Y103_SLICE_X85Y103_SR;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_A;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_A1;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_A2;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_A3;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_A4;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_A5;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_A6;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_AO5;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_AO6;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_AQ;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_AX;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_A_CY;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_A_XOR;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_B;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_B1;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_B2;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_B3;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_B4;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_B5;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_B6;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_BO5;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_BO6;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_BX;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_B_CY;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_B_XOR;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_C;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_C1;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_C2;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_C3;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_C4;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_C5;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_C6;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_CE;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_CIN;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_CLK;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_CO5;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_CO6;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_COUT;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_CX;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_C_CY;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_C_XOR;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_D;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_D1;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_D2;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_D3;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_D4;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_D5;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_D6;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_DO5;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_DO6;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_DX;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_D_CY;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_D_XOR;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X84Y104_SR;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_A;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_A1;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_A2;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_A3;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_A4;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_A5;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_A6;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_AO5;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_AO6;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_AQ;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_A_CY;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_A_XOR;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_B;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_B1;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_B2;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_B3;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_B4;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_B5;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_B6;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_BO5;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_BO6;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_B_CY;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_B_XOR;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_C;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_C1;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_C2;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_C3;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_C4;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_C5;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_C6;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_CE;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_CLK;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_CO5;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_CO6;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_C_CY;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_C_XOR;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_D;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_D1;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_D2;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_D3;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_D4;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_D5;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_D6;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_DO5;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_DO6;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_D_CY;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_D_XOR;
  wire [0:0] CLBLM_L_X56Y104_SLICE_X85Y104_SR;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_A;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_A1;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_A2;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_A3;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_A4;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_A5;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_A6;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_AO5;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_AO6;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_AQ;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_A_CY;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_A_XOR;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_B;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_B1;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_B2;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_B3;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_B4;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_B5;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_B6;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_BO5;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_BO6;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_BQ;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_B_CY;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_B_XOR;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_C;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_C1;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_C2;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_C3;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_C4;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_C5;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_C6;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_CE;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_CLK;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_CO5;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_CO6;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_CQ;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_C_CY;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_C_XOR;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_D;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_D1;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_D2;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_D3;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_D4;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_D5;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_D6;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_DO5;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_DO6;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_D_CY;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_D_XOR;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X84Y105_SR;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_A;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_A1;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_A2;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_A3;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_A4;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_A5;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_A6;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_AO5;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_AO6;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_AQ;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_A_CY;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_A_XOR;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_B;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_B1;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_B2;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_B3;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_B4;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_B5;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_B6;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_BO5;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_BO6;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_BQ;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_B_CY;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_B_XOR;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_C;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_C1;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_C2;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_C3;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_C4;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_C5;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_C6;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_CE;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_CLK;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_CO5;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_CO6;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_CQ;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_C_CY;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_C_XOR;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_D;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_D1;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_D2;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_D3;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_D4;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_D5;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_D6;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_DO5;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_DO6;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_DQ;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_D_CY;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_D_XOR;
  wire [0:0] CLBLM_L_X56Y105_SLICE_X85Y105_SR;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_A;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_A1;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_A2;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_A3;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_A4;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_A5;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_A6;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_AO5;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_AO6;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_AQ;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_A_CY;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_A_XOR;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_B;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_B1;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_B2;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_B3;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_B4;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_B5;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_B6;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_BO5;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_BO6;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_B_CY;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_B_XOR;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_C;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_C1;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_C2;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_C3;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_C4;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_C5;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_C6;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_CE;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_CLK;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_CO5;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_CO6;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_C_CY;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_C_XOR;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_D;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_D1;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_D2;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_D3;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_D4;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_D5;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_D6;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_DO5;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_DO6;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_D_CY;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_D_XOR;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X84Y111_SR;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_A;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_A1;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_A2;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_A3;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_A4;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_A5;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_A6;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_AO5;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_AO6;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_A_CY;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_A_XOR;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_B;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_B1;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_B2;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_B3;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_B4;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_B5;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_B6;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_BO5;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_BO6;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_B_CY;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_B_XOR;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_C;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_C1;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_C2;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_C3;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_C4;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_C5;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_C6;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_CO5;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_CO6;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_C_CY;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_C_XOR;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_D;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_D1;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_D2;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_D3;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_D4;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_D5;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_D6;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_DO5;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_DO6;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_D_CY;
  wire [0:0] CLBLM_L_X56Y111_SLICE_X85Y111_D_XOR;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_A;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_A1;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_A2;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_A3;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_A4;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_A5;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_A6;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_AMUX;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_AO5;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_AO6;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_A_CY;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_A_XOR;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_B;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_B1;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_B2;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_B3;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_B4;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_B5;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_B6;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_BO5;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_BO6;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_B_CY;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_B_XOR;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_C;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_C1;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_C2;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_C3;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_C4;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_C5;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_C6;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_CE;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_CLK;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_CMUX;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_CO5;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_CO6;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_C_CY;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_C_XOR;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_D;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_D1;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_D2;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_D3;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_D4;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_D5;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_D6;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_DO5;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_DO6;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_DQ;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_D_CY;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_D_XOR;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X84Y97_SR;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_A;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_A1;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_A2;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_A3;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_A4;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_A5;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_A6;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_AO5;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_AO6;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_AQ;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_A_CY;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_A_XOR;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_B;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_B1;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_B2;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_B3;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_B4;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_B5;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_B6;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_BMUX;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_BO5;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_BO6;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_B_CY;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_B_XOR;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_C;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_C1;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_C2;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_C3;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_C4;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_C5;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_C6;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_CE;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_CLK;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_CO5;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_CO6;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_CQ;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_C_CY;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_C_XOR;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_D;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_D1;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_D2;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_D3;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_D4;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_D5;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_D6;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_DO5;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_DO6;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_D_CY;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_D_XOR;
  wire [0:0] CLBLM_L_X56Y97_SLICE_X85Y97_SR;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_A;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_A1;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_A2;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_A3;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_A4;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_A5;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_A6;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_AMUX;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_AO5;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_AO6;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_AQ;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_A_CY;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_A_XOR;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_B;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_B1;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_B2;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_B3;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_B4;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_B5;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_B6;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_BMUX;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_BO5;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_BO6;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_BQ;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_BX;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_B_CY;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_B_XOR;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_C;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_C1;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_C2;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_C3;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_C4;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_C5;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_C6;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_CE;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_CLK;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_CMUX;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_CO5;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_CO6;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_C_CY;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_C_XOR;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_D;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_D1;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_D2;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_D3;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_D4;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_D5;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_D6;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_DMUX;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_DO5;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_DO6;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_D_CY;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_D_XOR;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X84Y98_SR;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_A;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_A1;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_A2;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_A3;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_A4;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_A5;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_A5Q;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_A6;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_AMUX;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_AO5;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_AO6;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_AQ;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_A_CY;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_A_XOR;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_B;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_B1;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_B2;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_B3;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_B4;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_B5;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_B6;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_BMUX;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_BO5;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_BO6;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_BQ;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_B_CY;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_B_XOR;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_C;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_C1;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_C2;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_C3;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_C4;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_C5;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_C6;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_CE;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_CLK;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_CO5;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_CO6;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_CQ;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_C_CY;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_C_XOR;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_D;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_D1;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_D2;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_D3;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_D4;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_D5;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_D6;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_DO5;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_DO6;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_DQ;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_D_CY;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_D_XOR;
  wire [0:0] CLBLM_L_X56Y98_SLICE_X85Y98_SR;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_A;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_A1;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_A2;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_A3;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_A4;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_A5;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_A6;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_AO5;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_AO6;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_AQ;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_A_CY;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_A_XOR;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_B;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_B1;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_B2;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_B3;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_B4;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_B5;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_B6;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_BO5;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_BO6;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_BQ;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_B_CY;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_B_XOR;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_C;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_C1;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_C2;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_C3;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_C4;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_C5;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_C6;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_CE;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_CLK;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_CO5;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_CO6;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_C_CY;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_C_XOR;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_D;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_D1;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_D2;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_D3;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_D4;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_D5;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_D6;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_DO5;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_DO6;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_D_CY;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_D_XOR;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X84Y99_SR;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_A;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_A1;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_A2;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_A3;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_A4;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_A5;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_A5Q;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_A6;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_AMUX;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_AO5;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_AO6;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_AQ;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_AX;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_A_CY;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_A_XOR;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_B;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_B1;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_B2;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_B3;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_B4;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_B5;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_B6;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_BO5;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_BO6;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_BQ;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_B_CY;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_B_XOR;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_C;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_C1;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_C2;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_C3;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_C4;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_C5;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_C6;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_CE;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_CLK;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_CO5;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_CO6;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_CQ;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_C_CY;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_C_XOR;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_D;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_D1;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_D2;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_D3;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_D4;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_D5;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_D6;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_DO5;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_DO6;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_D_CY;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_D_XOR;
  wire [0:0] CLBLM_L_X56Y99_SLICE_X85Y99_SR;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_A;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_A1;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_A2;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_A3;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_A4;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_A5;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_A6;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_AMUX;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_AO5;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_AO6;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_AQ;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_AX;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_A_CY;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_A_XOR;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_B;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_B1;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_B2;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_B3;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_B4;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_B5;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_B6;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_BO5;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_BO6;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_B_CY;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_B_XOR;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_C;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_C1;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_C2;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_C3;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_C4;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_C5;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_C6;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_CE;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_CLK;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_CO5;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_CO6;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_C_CY;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_C_XOR;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_D;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_D1;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_D2;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_D3;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_D4;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_D5;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_D6;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_DO5;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_DO6;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_D_CY;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_D_XOR;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X90Y100_SR;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_A;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_A1;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_A2;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_A3;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_A4;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_A5;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_A6;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_AMUX;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_AO5;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_AO6;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_A_CY;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_A_XOR;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_B;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_B1;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_B2;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_B3;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_B4;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_B5;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_B6;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_BO5;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_BO6;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_BQ;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_B_CY;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_B_XOR;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_C;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_C1;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_C2;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_C3;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_C4;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_C5;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_C6;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_CE;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_CLK;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_CMUX;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_CO5;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_CO6;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_C_CY;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_C_XOR;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_D;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_D1;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_D2;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_D3;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_D4;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_D5;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_D6;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_DO5;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_DO6;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_D_CY;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_D_XOR;
  wire [0:0] CLBLM_L_X60Y100_SLICE_X91Y100_SR;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_A;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_A1;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_A2;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_A3;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_A4;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_A5;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_A6;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_AO5;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_AO6;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_AQ;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_A_CY;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_A_XOR;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_B;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_B1;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_B2;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_B3;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_B4;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_B5;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_B6;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_BO5;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_BO6;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_B_CY;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_B_XOR;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_C;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_C1;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_C2;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_C3;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_C4;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_C5;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_C6;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_CE;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_CLK;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_CO5;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_CO6;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_C_CY;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_C_XOR;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_D;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_D1;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_D2;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_D3;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_D4;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_D5;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_D6;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_DO5;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_DO6;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_D_CY;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_D_XOR;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X90Y101_SR;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_A;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_A1;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_A2;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_A3;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_A4;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_A5;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_A6;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_AO5;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_AO6;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_AQ;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_A_CY;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_A_XOR;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_B;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_B1;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_B2;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_B3;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_B4;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_B5;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_B6;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_BO5;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_BO6;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_BQ;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_B_CY;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_B_XOR;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_C;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_C1;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_C2;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_C3;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_C4;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_C5;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_C6;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_CE;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_CLK;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_CMUX;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_CO5;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_CO6;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_C_CY;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_C_XOR;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_D;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_D1;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_D2;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_D3;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_D4;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_D5;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_D6;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_DO5;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_DO6;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_D_CY;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_D_XOR;
  wire [0:0] CLBLM_L_X60Y101_SLICE_X91Y101_SR;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_A;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_A1;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_A2;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_A3;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_A4;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_A5;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_A6;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_AO5;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_AO6;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_AQ;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_A_CY;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_A_XOR;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_B;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_B1;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_B2;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_B3;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_B4;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_B5;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_B6;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_BO5;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_BO6;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_BQ;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_B_CY;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_B_XOR;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_C;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_C1;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_C2;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_C3;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_C4;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_C5;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_C6;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_CE;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_CLK;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_CO5;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_CO6;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_CQ;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_C_CY;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_C_XOR;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_D;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_D1;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_D2;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_D3;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_D4;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_D5;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_D6;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_DO5;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_DO6;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_D_CY;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_D_XOR;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X90Y102_SR;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_A;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_A1;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_A2;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_A3;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_A4;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_A5;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_A6;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_AMUX;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_AO5;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_AO6;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_AX;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_A_CY;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_A_XOR;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_B;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_B1;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_B2;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_B3;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_B4;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_B5;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_B6;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_BMUX;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_BO5;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_BO6;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_BQ;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_BX;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_B_CY;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_B_XOR;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_C;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_C1;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_C2;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_C3;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_C4;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_C5;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_C6;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_CE;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_CLK;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_CMUX;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_CO5;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_CO6;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_COUT;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_CX;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_C_CY;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_C_XOR;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_D;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_D1;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_D2;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_D3;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_D4;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_D5;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_D6;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_DMUX;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_DO5;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_DO6;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_DX;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_D_CY;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_D_XOR;
  wire [0:0] CLBLM_L_X60Y102_SLICE_X91Y102_SR;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_A;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_A1;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_A2;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_A3;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_A4;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_A5;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_A6;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_AO5;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_AO6;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_AX;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_A_CY;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_A_XOR;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_B;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_B1;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_B2;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_B3;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_B4;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_B5;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_B6;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_BMUX;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_BO5;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_BO6;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_BX;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_B_CY;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_B_XOR;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_C;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_C1;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_C2;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_C3;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_C4;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_C5;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_C6;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_CO5;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_CO6;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_CX;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_C_CY;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_C_XOR;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_D;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_D1;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_D2;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_D3;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_D4;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_D5;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_D6;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_DO5;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_DO6;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_D_CY;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_D_XOR;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_F7AMUX_O;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_F7BMUX_O;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X90Y103_F8MUX_O;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_A;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_A1;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_A2;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_A3;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_A4;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_A5;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_A6;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_AMUX;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_AO5;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_AO6;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_AQ;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_AX;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_A_CY;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_A_XOR;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_B;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_B1;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_B2;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_B3;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_B4;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_B5;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_B6;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_BMUX;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_BO5;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_BO6;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_BX;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_B_CY;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_B_XOR;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_C;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_C1;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_C2;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_C3;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_C4;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_C5;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_C6;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_CE;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_CIN;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_CLK;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_CMUX;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_CO5;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_CO6;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_COUT;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_CX;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_C_CY;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_C_XOR;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_D;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_D1;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_D2;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_D3;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_D4;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_D5;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_D6;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_DMUX;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_DO5;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_DO6;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_DX;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_D_CY;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_D_XOR;
  wire [0:0] CLBLM_L_X60Y103_SLICE_X91Y103_SR;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_A;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_A1;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_A2;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_A3;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_A4;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_A5;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_A6;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_AO5;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_AO6;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_AQ;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_A_CY;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_A_XOR;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_B;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_B1;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_B2;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_B3;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_B4;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_B5;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_B6;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_BO5;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_BO6;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_B_CY;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_B_XOR;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_C;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_C1;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_C2;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_C3;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_C4;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_C5;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_C6;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_CE;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_CLK;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_CO5;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_CO6;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_C_CY;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_C_XOR;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_D;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_D1;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_D2;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_D3;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_D4;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_D5;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_D6;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_DO5;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_DO6;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_D_CY;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_D_XOR;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X90Y104_SR;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_A;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_A1;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_A2;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_A3;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_A4;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_A5;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_A6;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_AMUX;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_AO5;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_AO6;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_AQ;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_AX;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_A_CY;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_A_XOR;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_B;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_B1;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_B2;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_B3;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_B4;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_B5;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_B6;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_BMUX;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_BO5;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_BO6;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_BX;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_B_CY;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_B_XOR;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_C;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_C1;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_C2;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_C3;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_C4;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_C5;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_C6;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_CE;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_CIN;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_CLK;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_CMUX;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_CO5;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_CO6;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_COUT;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_CX;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_C_CY;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_C_XOR;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_D;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_D1;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_D2;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_D3;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_D4;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_D5;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_D6;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_DO5;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_DO6;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_DX;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_D_CY;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_D_XOR;
  wire [0:0] CLBLM_L_X60Y104_SLICE_X91Y104_SR;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_A;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_A1;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_A2;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_A3;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_A4;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_A5;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_A6;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_AMUX;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_AO5;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_AO6;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_AX;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_A_CY;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_A_XOR;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_B;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_B1;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_B2;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_B3;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_B4;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_B5;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_B6;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_BMUX;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_BO5;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_BO6;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_BX;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_B_CY;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_B_XOR;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_C;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_C1;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_C2;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_C3;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_C4;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_C5;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_C6;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_CMUX;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_CO5;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_CO6;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_COUT;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_CX;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_C_CY;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_C_XOR;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_D;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_D1;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_D2;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_D3;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_D4;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_D5;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_D6;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_DMUX;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_DO5;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_DO6;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_DX;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_D_CY;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X90Y105_D_XOR;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_A;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_A1;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_A2;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_A3;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_A4;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_A5;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_A6;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_AMUX;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_AO5;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_AO6;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_AX;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_A_CY;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_A_XOR;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_B;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_B1;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_B2;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_B3;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_B4;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_B5;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_B6;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_BMUX;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_BO5;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_BO6;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_BX;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_B_CY;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_B_XOR;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_C;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_C1;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_C2;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_C3;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_C4;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_C5;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_C6;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_CMUX;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_CO5;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_CO6;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_COUT;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_CX;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_C_CY;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_C_XOR;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_D;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_D1;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_D2;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_D3;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_D4;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_D5;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_D6;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_DMUX;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_DO5;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_DO6;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_DX;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_D_CY;
  wire [0:0] CLBLM_L_X60Y105_SLICE_X91Y105_D_XOR;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_A;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_A1;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_A2;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_A3;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_A4;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_A5;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_A6;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_AMUX;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_AO5;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_AO6;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_AQ;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_AX;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_A_CY;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_A_XOR;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_B;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_B1;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_B2;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_B3;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_B4;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_B5;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_B6;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_BMUX;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_BO5;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_BO6;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_BX;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_B_CY;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_B_XOR;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_C;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_C1;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_C2;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_C3;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_C4;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_C5;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_C6;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_CE;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_CIN;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_CLK;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_CMUX;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_CO5;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_CO6;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_COUT;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_CX;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_C_CY;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_C_XOR;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_D;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_D1;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_D2;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_D3;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_D4;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_D5;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_D6;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_DMUX;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_DO5;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_DO6;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_DX;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_D_CY;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_D_XOR;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X90Y106_SR;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_A;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_A1;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_A2;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_A3;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_A4;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_A5;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_A6;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_AMUX;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_AO5;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_AO6;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_AX;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_A_CY;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_A_XOR;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_B;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_B1;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_B2;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_B3;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_B4;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_B5;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_B6;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_BMUX;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_BO5;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_BO6;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_BX;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_B_CY;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_B_XOR;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_C;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_C1;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_C2;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_C3;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_C4;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_C5;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_C6;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_CIN;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_CMUX;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_CO5;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_CO6;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_COUT;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_CX;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_C_CY;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_C_XOR;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_D;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_D1;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_D2;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_D3;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_D4;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_D5;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_D6;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_DMUX;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_DO5;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_DO6;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_DX;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_D_CY;
  wire [0:0] CLBLM_L_X60Y106_SLICE_X91Y106_D_XOR;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_A;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_A1;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_A2;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_A3;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_A4;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_A5;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_A6;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_AMUX;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_AO5;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_AO6;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_AQ;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_AX;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_A_CY;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_A_XOR;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_B;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_B1;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_B2;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_B3;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_B4;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_B5;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_B6;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_BMUX;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_BO5;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_BO6;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_BX;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_B_CY;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_B_XOR;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_C;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_C1;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_C2;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_C3;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_C4;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_C5;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_C6;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_CE;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_CIN;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_CLK;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_CMUX;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_CO5;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_CO6;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_COUT;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_CX;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_C_CY;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_C_XOR;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_D;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_D1;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_D2;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_D3;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_D4;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_D5;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_D6;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_DMUX;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_DO5;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_DO6;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_DX;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_D_CY;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_D_XOR;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X90Y107_SR;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_A;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_A1;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_A2;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_A3;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_A4;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_A5;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_A6;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_AMUX;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_AO5;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_AO6;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_AQ;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_AX;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_A_CY;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_A_XOR;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_B;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_B1;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_B2;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_B3;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_B4;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_B5;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_B6;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_BMUX;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_BO5;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_BO6;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_BX;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_B_CY;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_B_XOR;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_C;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_C1;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_C2;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_C3;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_C4;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_C5;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_C6;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_CE;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_CIN;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_CLK;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_CMUX;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_CO5;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_CO6;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_COUT;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_CX;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_C_CY;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_C_XOR;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_D;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_D1;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_D2;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_D3;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_D4;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_D5;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_D6;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_DO5;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_DO6;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_DX;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_D_CY;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_D_XOR;
  wire [0:0] CLBLM_L_X60Y107_SLICE_X91Y107_SR;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_A;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_A1;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_A2;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_A3;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_A4;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_A5;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_A6;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_AMUX;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_AO5;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_AO6;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_AX;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_A_CY;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_A_XOR;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_B;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_B1;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_B2;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_B3;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_B4;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_B5;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_B6;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_BMUX;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_BO5;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_BO6;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_BQ;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_BX;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_B_CY;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_B_XOR;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_C;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_C1;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_C2;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_C3;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_C4;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_C5;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_C6;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_CE;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_CLK;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_CMUX;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_CO5;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_CO6;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_COUT;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_CX;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_C_CY;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_C_XOR;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_D;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_D1;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_D2;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_D3;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_D4;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_D5;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_D6;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_DMUX;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_DO5;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_DO6;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_DX;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_D_CY;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_D_XOR;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X90Y108_SR;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_A;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_A1;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_A2;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_A3;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_A4;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_A5;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_A6;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_AO5;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_AO6;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_AQ;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_A_CY;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_A_XOR;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_B;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_B1;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_B2;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_B3;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_B4;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_B5;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_B6;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_BO5;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_BO6;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_B_CY;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_B_XOR;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_C;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_C1;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_C2;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_C3;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_C4;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_C5;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_C6;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_CE;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_CLK;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_CO5;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_CO6;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_C_CY;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_C_XOR;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_D;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_D1;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_D2;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_D3;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_D4;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_D5;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_D6;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_DO5;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_DO6;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_D_CY;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_D_XOR;
  wire [0:0] CLBLM_L_X60Y108_SLICE_X91Y108_SR;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_A;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_A1;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_A2;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_A3;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_A4;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_A5;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_A6;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_AMUX;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_AO5;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_AO6;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_AX;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_A_CY;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_A_XOR;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_B;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_B1;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_B2;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_B3;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_B4;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_B5;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_B6;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_BMUX;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_BO5;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_BO6;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_BX;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_B_CY;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_B_XOR;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_C;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_C1;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_C2;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_C3;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_C4;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_C5;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_C6;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_CIN;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_CMUX;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_CO5;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_CO6;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_COUT;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_CX;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_C_CY;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_C_XOR;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_D;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_D1;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_D2;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_D3;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_D4;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_D5;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_D6;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_DMUX;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_DO5;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_DO6;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_DX;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_D_CY;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X90Y109_D_XOR;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_A;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_A1;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_A2;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_A3;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_A4;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_A5;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_A6;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_AO5;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_AO6;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_AQ;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_A_CY;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_A_XOR;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_B;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_B1;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_B2;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_B3;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_B4;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_B5;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_B6;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_BO5;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_BO6;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_BQ;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_B_CY;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_B_XOR;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_C;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_C1;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_C2;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_C3;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_C4;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_C5;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_C6;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_CE;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_CLK;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_CO5;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_CO6;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_C_CY;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_C_XOR;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_D;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_D1;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_D2;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_D3;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_D4;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_D5;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_D6;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_DO5;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_DO6;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_D_CY;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_D_XOR;
  wire [0:0] CLBLM_L_X60Y109_SLICE_X91Y109_SR;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_A;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_A1;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_A2;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_A3;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_A4;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_A5;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_A6;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_AMUX;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_AO5;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_AO6;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_AX;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_A_CY;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_A_XOR;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_B;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_B1;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_B2;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_B3;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_B4;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_B5;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_B6;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_BMUX;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_BO5;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_BO6;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_BX;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_B_CY;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_B_XOR;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_C;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_C1;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_C2;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_C3;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_C4;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_C5;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_C6;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_CIN;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_CMUX;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_CO5;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_CO6;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_COUT;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_CX;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_C_CY;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_C_XOR;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_D;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_D1;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_D2;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_D3;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_D4;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_D5;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_D6;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_DO5;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_DO6;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_DX;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_D_CY;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X90Y110_D_XOR;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_A;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_A1;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_A2;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_A3;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_A4;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_A5;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_A6;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_AO5;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_AO6;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_AQ;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_A_CY;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_A_XOR;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_B;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_B1;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_B2;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_B3;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_B4;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_B5;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_B6;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_BO5;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_BO6;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_B_CY;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_B_XOR;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_C;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_C1;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_C2;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_C3;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_C4;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_C5;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_C6;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_CE;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_CLK;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_CO5;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_CO6;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_C_CY;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_C_XOR;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_D;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_D1;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_D2;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_D3;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_D4;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_D5;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_D6;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_DO5;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_DO6;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_D_CY;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_D_XOR;
  wire [0:0] CLBLM_L_X60Y110_SLICE_X91Y110_SR;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_A;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_A1;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_A2;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_A3;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_A4;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_A5;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_A6;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_AO5;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_AO6;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_AQ;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_A_CY;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_A_XOR;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_B;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_B1;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_B2;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_B3;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_B4;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_B5;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_B6;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_BO5;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_BO6;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_B_CY;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_B_XOR;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_C;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_C1;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_C2;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_C3;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_C4;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_C5;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_C6;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_CE;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_CLK;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_CO5;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_CO6;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_C_CY;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_C_XOR;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_D;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_D1;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_D2;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_D3;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_D4;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_D5;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_D6;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_DO5;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_DO6;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_D_CY;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_D_XOR;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X90Y111_SR;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_A;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_A1;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_A2;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_A3;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_A4;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_A5;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_A6;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_AO5;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_AO6;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_AQ;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_A_CY;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_A_XOR;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_B;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_B1;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_B2;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_B3;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_B4;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_B5;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_B6;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_BO5;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_BO6;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_BQ;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_B_CY;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_B_XOR;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_C;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_C1;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_C2;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_C3;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_C4;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_C5;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_C6;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_CE;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_CLK;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_CO5;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_CO6;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_C_CY;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_C_XOR;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_D;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_D1;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_D2;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_D3;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_D4;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_D5;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_D6;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_DO5;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_DO6;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_D_CY;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_D_XOR;
  wire [0:0] CLBLM_L_X60Y111_SLICE_X91Y111_SR;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_A;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_A1;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_A2;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_A3;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_A4;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_A5;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_A6;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_AO5;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_AO6;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_A_CY;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_A_XOR;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_B;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_B1;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_B2;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_B3;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_B4;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_B5;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_B6;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_BO5;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_BO6;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_B_CY;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_B_XOR;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_C;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_C1;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_C2;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_C3;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_C4;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_C5;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_C6;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_CO5;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_CO6;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_C_CY;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_C_XOR;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_D;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_D1;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_D2;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_D3;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_D4;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_D5;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_D6;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_DO5;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_DO6;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_D_CY;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X90Y112_D_XOR;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_A;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_A1;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_A2;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_A3;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_A4;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_A5;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_A6;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_AO5;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_AO6;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_A_CY;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_A_XOR;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_B;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_B1;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_B2;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_B3;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_B4;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_B5;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_B6;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_BO5;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_BO6;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_B_CY;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_B_XOR;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_C;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_C1;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_C2;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_C3;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_C4;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_C5;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_C6;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_CO5;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_CO6;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_C_CY;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_C_XOR;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_D;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_D1;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_D2;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_D3;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_D4;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_D5;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_D6;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_DO5;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_DO6;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_D_CY;
  wire [0:0] CLBLM_L_X60Y112_SLICE_X91Y112_D_XOR;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_A;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_A1;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_A2;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_A3;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_A4;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_A5;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_A6;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_AO5;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_AO6;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_AQ;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_AX;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_A_CY;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_A_XOR;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_B;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_B1;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_B2;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_B3;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_B4;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_B5;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_B6;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_BO5;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_BO6;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_BQ;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_BX;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_B_CY;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_B_XOR;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_C;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_C1;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_C2;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_C3;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_C4;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_C5;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_C6;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_CE;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_CLK;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_CO5;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_CO6;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_C_CY;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_C_XOR;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_D;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_D1;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_D2;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_D3;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_D4;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_D5;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_D6;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_DO5;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_DO6;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_D_CY;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_D_XOR;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X90Y96_SR;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_A;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_A1;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_A2;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_A3;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_A4;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_A5;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_A6;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_AO5;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_AO6;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_A_CY;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_A_XOR;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_B;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_B1;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_B2;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_B3;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_B4;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_B5;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_B6;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_BO5;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_BO6;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_B_CY;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_B_XOR;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_C;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_C1;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_C2;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_C3;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_C4;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_C5;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_C6;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_CO5;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_CO6;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_C_CY;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_C_XOR;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_D;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_D1;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_D2;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_D3;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_D4;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_D5;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_D6;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_DO5;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_DO6;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_D_CY;
  wire [0:0] CLBLM_L_X60Y96_SLICE_X91Y96_D_XOR;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_A;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_A1;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_A2;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_A3;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_A4;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_A5;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_A5Q;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_A6;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_AMUX;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_AO5;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_AO6;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_AX;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_A_CY;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_A_XOR;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_B;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_B1;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_B2;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_B3;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_B4;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_B5;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_B6;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_BO5;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_BO6;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_BQ;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_BX;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_B_CY;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_B_XOR;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_C;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_C1;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_C2;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_C3;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_C4;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_C5;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_C6;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_CE;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_CLK;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_CO5;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_CO6;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_CX;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_C_CY;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_C_XOR;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_D;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_D1;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_D2;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_D3;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_D4;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_D5;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_D6;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_DO5;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_DO6;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_D_CY;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_D_XOR;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X90Y97_SR;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_A;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_A1;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_A2;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_A3;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_A4;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_A5;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_A6;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_AMUX;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_AO5;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_AO6;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_AQ;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_AX;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_A_CY;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_A_XOR;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_B;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_B1;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_B2;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_B3;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_B4;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_B5;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_B6;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_BO5;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_BO6;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_BQ;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_B_CY;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_B_XOR;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_C;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_C1;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_C2;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_C3;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_C4;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_C5;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_C6;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_CE;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_CLK;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_CO5;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_CO6;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_C_CY;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_C_XOR;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_D;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_D1;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_D2;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_D3;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_D4;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_D5;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_D6;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_DO5;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_DO6;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_D_CY;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_D_XOR;
  wire [0:0] CLBLM_L_X60Y97_SLICE_X91Y97_SR;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_A;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_A1;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_A2;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_A3;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_A4;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_A5;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_A6;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_AO5;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_AO6;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_AQ;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_A_CY;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_A_XOR;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_B;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_B1;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_B2;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_B3;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_B4;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_B5;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_B6;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_BO5;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_BO6;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_BQ;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_B_CY;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_B_XOR;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_C;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_C1;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_C2;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_C3;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_C4;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_C5;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_C6;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_CLK;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_CMUX;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_CO5;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_CO6;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_C_CY;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_C_XOR;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_D;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_D1;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_D2;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_D3;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_D4;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_D5;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_D6;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_DO5;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_DO6;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_D_CY;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_D_XOR;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X90Y98_SR;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_A;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_A1;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_A2;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_A3;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_A4;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_A5;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_A6;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_AMUX;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_AO5;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_AO6;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_AQ;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_AX;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_A_CY;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_A_XOR;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_B;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_B1;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_B2;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_B3;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_B4;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_B5;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_B6;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_BO5;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_BO6;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_BQ;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_BX;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_B_CY;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_B_XOR;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_C;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_C1;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_C2;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_C3;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_C4;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_C5;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_C6;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_CE;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_CLK;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_CO5;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_CO6;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_CQ;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_CX;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_C_CY;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_C_XOR;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_D;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_D1;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_D2;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_D3;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_D4;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_D5;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_D6;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_DO5;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_DO6;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_DQ;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_DX;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_D_CY;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_D_XOR;
  wire [0:0] CLBLM_L_X60Y98_SLICE_X91Y98_SR;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_A;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_A1;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_A2;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_A3;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_A4;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_A5;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_A6;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_AMUX;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_AO5;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_AO6;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_AQ;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_AX;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_A_CY;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_A_XOR;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_B;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_B1;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_B2;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_B3;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_B4;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_B5;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_B6;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_BMUX;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_BO5;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_BO6;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_B_CY;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_B_XOR;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_C;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_C1;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_C2;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_C3;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_C4;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_C5;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_C6;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_CE;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_CLK;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_CO5;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_CO6;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_CQ;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_C_CY;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_C_XOR;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_D;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_D1;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_D2;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_D3;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_D4;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_D5;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_D6;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_DO5;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_DO6;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_D_CY;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_D_XOR;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X90Y99_SR;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_A;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_A1;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_A2;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_A3;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_A4;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_A5;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_A6;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_AMUX;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_AO5;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_AO6;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_A_CY;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_A_XOR;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_B;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_B1;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_B2;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_B3;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_B4;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_B5;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_B6;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_BMUX;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_BO5;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_BO6;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_B_CY;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_B_XOR;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_C;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_C1;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_C2;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_C3;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_C4;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_C5;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_C6;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_CMUX;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_CO5;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_CO6;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_C_CY;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_C_XOR;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_D;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_D1;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_D2;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_D3;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_D4;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_D5;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_D6;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_DO5;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_DO6;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_D_CY;
  wire [0:0] CLBLM_L_X60Y99_SLICE_X91Y99_D_XOR;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_A;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_A1;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_A2;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_A3;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_A4;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_A5;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_A6;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_AMUX;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_AO5;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_AO6;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_AQ;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_AX;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_A_CY;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_A_XOR;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_B;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_B1;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_B2;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_B3;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_B4;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_B5;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_B6;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_BO5;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_BO6;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_BQ;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_BX;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_B_CY;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_B_XOR;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_C;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_C1;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_C2;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_C3;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_C4;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_C5;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_C6;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_CE;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_CLK;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_CO5;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_CO6;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_CQ;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_CX;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_C_CY;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_C_XOR;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_D;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_D1;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_D2;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_D3;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_D4;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_D5;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_D6;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_DO5;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_DO6;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_D_CY;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_D_XOR;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X92Y100_SR;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_A;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_A1;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_A2;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_A3;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_A4;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_A5;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_A6;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_AO5;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_AO6;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_AQ;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_A_CY;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_A_XOR;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_B;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_B1;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_B2;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_B3;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_B4;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_B5;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_B6;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_BO5;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_BO6;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_BQ;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_B_CY;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_B_XOR;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_C;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_C1;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_C2;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_C3;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_C4;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_C5;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_C6;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_CE;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_CLK;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_CO5;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_CO6;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_C_CY;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_C_XOR;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_D;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_D1;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_D2;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_D3;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_D4;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_D5;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_D6;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_DO5;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_DO6;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_D_CY;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_D_XOR;
  wire [0:0] CLBLM_L_X62Y100_SLICE_X93Y100_SR;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_A;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_A1;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_A2;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_A3;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_A4;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_A5;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_A6;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_AO5;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_AO6;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_AQ;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_A_CY;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_A_XOR;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_B;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_B1;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_B2;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_B3;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_B4;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_B5;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_B6;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_BO5;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_BO6;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_BQ;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_B_CY;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_B_XOR;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_C;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_C1;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_C2;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_C3;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_C4;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_C5;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_C6;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_CE;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_CLK;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_CO5;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_CO6;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_CQ;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_C_CY;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_C_XOR;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_D;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_D1;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_D2;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_D3;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_D4;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_D5;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_D6;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_DMUX;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_DO5;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_DO6;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_D_CY;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_D_XOR;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X92Y101_SR;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_A;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_A1;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_A2;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_A3;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_A4;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_A5;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_A6;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_AO5;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_AO6;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_AQ;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_AX;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_A_CY;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_A_XOR;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_B;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_B1;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_B2;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_B3;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_B4;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_B5;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_B6;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_BO5;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_BO6;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_BQ;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_BX;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_B_CY;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_B_XOR;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_C;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_C1;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_C2;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_C3;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_C4;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_C5;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_C6;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_CE;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_CLK;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_CO5;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_CO6;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_CQ;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_CX;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_C_CY;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_C_XOR;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_D;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_D1;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_D2;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_D3;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_D4;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_D5;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_D6;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_DO5;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_DO6;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_D_CY;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_D_XOR;
  wire [0:0] CLBLM_L_X62Y101_SLICE_X93Y101_SR;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_A;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_A1;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_A2;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_A3;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_A4;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_A5;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_A6;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_AMUX;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_AO5;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_AO6;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_A_CY;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_A_XOR;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_B;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_B1;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_B2;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_B3;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_B4;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_B5;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_B6;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_BO5;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_BO6;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_BQ;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_B_CY;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_B_XOR;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_C;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_C1;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_C2;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_C3;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_C4;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_C5;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_C6;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_CE;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_CLK;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_CO5;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_CO6;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_C_CY;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_C_XOR;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_D;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_D1;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_D2;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_D3;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_D4;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_D5;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_D6;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_DMUX;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_DO5;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_DO6;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_D_CY;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_D_XOR;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X92Y102_SR;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_A;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_A1;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_A2;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_A3;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_A4;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_A5;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_A6;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_AMUX;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_AO5;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_AO6;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_A_CY;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_A_XOR;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_B;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_B1;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_B2;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_B3;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_B4;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_B5;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_B6;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_BO5;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_BO6;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_B_CY;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_B_XOR;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_C;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_C1;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_C2;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_C3;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_C4;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_C5;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_C6;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_CO5;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_CO6;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_C_CY;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_C_XOR;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_D;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_D1;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_D2;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_D3;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_D4;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_D5;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_D6;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_DO5;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_DO6;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_D_CY;
  wire [0:0] CLBLM_L_X62Y102_SLICE_X93Y102_D_XOR;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_A;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_A1;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_A2;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_A3;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_A4;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_A5;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_A6;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_AO5;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_AO6;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_AQ;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_A_CY;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_A_XOR;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_B;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_B1;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_B2;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_B3;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_B4;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_B5;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_B6;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_BO5;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_BO6;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_B_CY;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_B_XOR;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_C;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_C1;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_C2;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_C3;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_C4;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_C5;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_C6;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_CE;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_CLK;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_CMUX;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_CO5;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_CO6;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_C_CY;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_C_XOR;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_D;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_D1;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_D2;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_D3;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_D4;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_D5;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_D6;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_DO5;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_DO6;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_D_CY;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_D_XOR;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X92Y103_SR;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_A;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_A1;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_A2;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_A3;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_A4;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_A5;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_A6;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_AO5;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_AO6;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_AQ;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_A_CY;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_A_XOR;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_B;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_B1;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_B2;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_B3;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_B4;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_B5;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_B6;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_BO5;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_BO6;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_B_CY;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_B_XOR;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_C;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_C1;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_C2;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_C3;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_C4;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_C5;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_C6;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_CE;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_CLK;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_CO5;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_CO6;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_C_CY;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_C_XOR;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_D;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_D1;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_D2;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_D3;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_D4;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_D5;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_D6;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_DO5;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_DO6;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_D_CY;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_D_XOR;
  wire [0:0] CLBLM_L_X62Y103_SLICE_X93Y103_SR;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_A;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_A1;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_A2;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_A3;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_A4;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_A5;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_A6;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_AO5;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_AO6;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_AQ;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_A_CY;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_A_XOR;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_B;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_B1;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_B2;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_B3;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_B4;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_B5;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_B6;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_BO5;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_BO6;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_BQ;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_B_CY;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_B_XOR;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_C;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_C1;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_C2;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_C3;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_C4;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_C5;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_C6;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_CE;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_CLK;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_CMUX;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_CO5;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_CO6;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_C_CY;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_C_XOR;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_D;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_D1;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_D2;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_D3;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_D4;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_D5;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_D6;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_DO5;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_DO6;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_D_CY;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_D_XOR;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X92Y104_SR;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_A;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_A1;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_A2;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_A3;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_A4;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_A5;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_A6;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_AO5;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_AO6;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_AQ;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_A_CY;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_A_XOR;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_B;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_B1;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_B2;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_B3;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_B4;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_B5;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_B6;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_BO5;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_BO6;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_B_CY;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_B_XOR;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_C;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_C1;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_C2;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_C3;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_C4;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_C5;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_C6;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_CE;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_CLK;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_CO5;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_CO6;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_C_CY;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_C_XOR;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_D;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_D1;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_D2;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_D3;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_D4;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_D5;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_D6;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_DO5;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_DO6;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_D_CY;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_D_XOR;
  wire [0:0] CLBLM_L_X62Y104_SLICE_X93Y104_SR;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_A;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_A1;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_A2;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_A3;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_A4;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_A5;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_A6;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_AMUX;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_AO5;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_AO6;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_A_CY;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_A_XOR;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_B;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_B1;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_B2;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_B3;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_B4;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_B5;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_B6;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_BMUX;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_BO5;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_BO6;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_B_CY;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_B_XOR;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_C;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_C1;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_C2;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_C3;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_C4;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_C5;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_C6;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_CE;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_CLK;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_CO5;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_CO6;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_CQ;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_C_CY;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_C_XOR;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_D;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_D1;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_D2;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_D3;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_D4;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_D5;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_D6;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_DO5;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_DO6;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_D_CY;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_D_XOR;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X92Y105_SR;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_A;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_A1;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_A2;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_A3;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_A4;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_A5;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_A6;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_AMUX;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_AO5;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_AO6;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_A_CY;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_A_XOR;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_B;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_B1;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_B2;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_B3;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_B4;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_B5;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_B6;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_BO5;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_BO6;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_BQ;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_B_CY;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_B_XOR;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_C;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_C1;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_C2;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_C3;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_C4;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_C5;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_C6;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_CE;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_CLK;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_CO5;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_CO6;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_C_CY;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_C_XOR;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_D;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_D1;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_D2;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_D3;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_D4;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_D5;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_D6;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_DO5;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_DO6;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_D_CY;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_D_XOR;
  wire [0:0] CLBLM_L_X62Y105_SLICE_X93Y105_SR;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_A;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_A1;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_A2;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_A3;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_A4;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_A5;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_A6;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_AMUX;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_AO5;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_AO6;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_A_CY;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_A_XOR;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_B;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_B1;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_B2;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_B3;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_B4;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_B5;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_B6;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_BO5;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_BO6;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_BQ;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_B_CY;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_B_XOR;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_C;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_C1;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_C2;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_C3;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_C4;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_C5;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_C6;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_CE;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_CLK;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_CO5;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_CO6;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_CQ;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_C_CY;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_C_XOR;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_D;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_D1;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_D2;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_D3;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_D4;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_D5;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_D6;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_DO5;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_DO6;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_D_CY;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_D_XOR;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X92Y106_SR;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_A;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_A1;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_A2;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_A3;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_A4;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_A5;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_A6;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_AO5;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_AO6;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_AQ;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_A_CY;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_A_XOR;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_B;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_B1;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_B2;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_B3;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_B4;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_B5;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_B6;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_BMUX;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_BO5;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_BO6;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_B_CY;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_B_XOR;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_C;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_C1;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_C2;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_C3;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_C4;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_C5;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_C6;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_CE;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_CLK;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_CMUX;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_CO5;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_CO6;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_C_CY;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_C_XOR;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_D;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_D1;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_D2;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_D3;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_D4;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_D5;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_D6;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_DO5;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_DO6;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_D_CY;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_D_XOR;
  wire [0:0] CLBLM_L_X62Y106_SLICE_X93Y106_SR;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_A;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_A1;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_A2;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_A3;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_A4;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_A5;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_A5Q;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_A6;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_AMUX;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_AO5;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_AO6;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_AQ;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_AX;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_A_CY;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_A_XOR;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_B;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_B1;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_B2;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_B3;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_B4;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_B5;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_B6;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_BMUX;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_BO5;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_BO6;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_BQ;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_B_CY;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_B_XOR;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_C;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_C1;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_C2;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_C3;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_C4;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_C5;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_C6;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_CE;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_CLK;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_CO5;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_CO6;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_C_CY;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_C_XOR;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_D;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_D1;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_D2;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_D3;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_D4;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_D5;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_D6;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_DO5;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_DO6;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_D_CY;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_D_XOR;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X92Y107_SR;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_A;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_A1;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_A2;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_A3;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_A4;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_A5;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_A6;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_AO5;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_A_CY;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_A_XOR;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_B;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_B1;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_B2;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_B3;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_B4;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_B5;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_B6;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_BMUX;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_BO5;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_B_CY;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_B_XOR;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_C;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_C1;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_C2;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_C3;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_C4;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_C5;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_C6;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_CO5;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_CO6;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_C_CY;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_C_XOR;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_D;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_D1;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_D2;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_D3;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_D4;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_D5;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_D6;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_DO5;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_DO6;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_D_CY;
  wire [0:0] CLBLM_L_X62Y107_SLICE_X93Y107_D_XOR;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_A;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_A1;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_A2;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_A3;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_A4;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_A5;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_A5Q;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_A6;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_AMUX;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_AO5;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_AO6;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_AQ;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_A_CY;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_A_XOR;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_B;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_B1;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_B2;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_B3;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_B4;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_B5;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_B6;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_BMUX;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_BO5;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_BO6;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_B_CY;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_B_XOR;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_C;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_C1;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_C2;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_C3;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_C4;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_C5;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_C6;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_CE;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_CLK;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_CO5;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_CO6;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_C_CY;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_C_XOR;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_D;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_D1;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_D2;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_D3;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_D4;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_D5;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_D6;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_DO5;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_DO6;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_D_CY;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_D_XOR;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X92Y108_SR;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_A;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_A1;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_A2;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_A3;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_A4;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_A5;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_A6;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_AO5;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_AO6;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_AQ;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_A_CY;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_A_XOR;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_B;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_B1;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_B2;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_B3;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_B4;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_B5;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_B6;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_BO5;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_BO6;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_B_CY;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_B_XOR;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_C;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_C1;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_C2;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_C3;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_C4;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_C5;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_C6;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_CE;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_CLK;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_CO5;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_CO6;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_C_CY;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_C_XOR;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_D;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_D1;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_D2;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_D3;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_D4;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_D5;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_D6;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_DO5;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_DO6;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_D_CY;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_D_XOR;
  wire [0:0] CLBLM_L_X62Y108_SLICE_X93Y108_SR;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_A;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_A1;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_A2;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_A3;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_A4;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_A5;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_A6;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_AO5;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_AO6;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_A_CY;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_A_XOR;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_B;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_B1;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_B2;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_B3;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_B4;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_B5;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_B6;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_BO5;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_BO6;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_B_CY;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_B_XOR;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_C;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_C1;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_C2;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_C3;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_C4;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_C5;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_C6;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_CO5;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_CO6;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_C_CY;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_C_XOR;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_D;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_D1;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_D2;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_D3;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_D4;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_D5;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_D6;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_DO5;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_DO6;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_D_CY;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X92Y109_D_XOR;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_A;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_A1;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_A2;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_A3;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_A4;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_A5;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_A6;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_AO5;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_AO6;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_A_CY;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_A_XOR;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_B;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_B1;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_B2;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_B3;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_B4;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_B5;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_B6;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_BO5;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_BO6;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_B_CY;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_B_XOR;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_C;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_C1;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_C2;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_C3;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_C4;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_C5;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_C6;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_CO5;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_CO6;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_C_CY;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_C_XOR;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_D;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_D1;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_D2;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_D3;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_D4;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_D5;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_D6;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_DO5;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_DO6;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_D_CY;
  wire [0:0] CLBLM_L_X62Y109_SLICE_X93Y109_D_XOR;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_A;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_A1;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_A2;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_A3;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_A4;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_A5;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_A6;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_AO5;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_AO6;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_AQ;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_A_CY;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_A_XOR;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_B;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_B1;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_B2;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_B3;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_B4;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_B5;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_B6;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_BO5;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_BO6;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_BQ;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_B_CY;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_B_XOR;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_C;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_C1;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_C2;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_C3;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_C4;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_C5;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_C6;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_CE;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_CLK;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_CO5;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_CO6;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_C_CY;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_C_XOR;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_D;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_D1;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_D2;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_D3;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_D4;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_D5;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_D6;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_DO5;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_DO6;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_D_CY;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_D_XOR;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X92Y110_SR;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_A;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_A1;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_A2;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_A3;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_A4;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_A5;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_A6;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_AO5;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_AO6;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_AQ;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_A_CY;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_A_XOR;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_B;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_B1;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_B2;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_B3;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_B4;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_B5;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_B6;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_BO5;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_BO6;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_B_CY;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_B_XOR;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_C;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_C1;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_C2;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_C3;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_C4;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_C5;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_C6;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_CLK;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_CMUX;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_CO5;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_CO6;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_C_CY;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_C_XOR;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_D;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_D1;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_D2;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_D3;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_D4;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_D5;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_D6;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_DO5;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_DO6;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_D_CY;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_D_XOR;
  wire [0:0] CLBLM_L_X62Y110_SLICE_X93Y110_SR;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_A;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_A1;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_A2;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_A3;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_A4;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_A5;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_A5Q;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_A6;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_AMUX;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_AO5;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_AO6;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_AQ;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_A_CY;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_A_XOR;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_B;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_B1;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_B2;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_B3;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_B4;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_B5;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_B6;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_BO5;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_BO6;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_B_CY;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_B_XOR;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_C;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_C1;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_C2;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_C3;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_C4;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_C5;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_C6;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_CE;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_CLK;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_CO5;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_CO6;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_C_CY;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_C_XOR;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_D;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_D1;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_D2;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_D3;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_D4;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_D5;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_D6;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_DO5;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_DO6;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_D_CY;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_D_XOR;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X92Y111_SR;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_A;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_A1;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_A2;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_A3;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_A4;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_A5;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_A6;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_AO5;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_AO6;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_A_CY;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_A_XOR;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_B;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_B1;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_B2;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_B3;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_B4;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_B5;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_B6;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_BO5;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_BO6;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_B_CY;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_B_XOR;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_C;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_C1;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_C2;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_C3;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_C4;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_C5;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_C6;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_CO5;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_CO6;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_C_CY;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_C_XOR;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_D;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_D1;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_D2;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_D3;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_D4;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_D5;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_D6;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_DO5;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_DO6;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_D_CY;
  wire [0:0] CLBLM_L_X62Y111_SLICE_X93Y111_D_XOR;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_A;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_A1;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_A2;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_A3;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_A4;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_A5;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_A6;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_AO5;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_AO6;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_A_CY;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_A_XOR;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_B;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_B1;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_B2;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_B3;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_B4;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_B5;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_B6;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_BO5;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_BO6;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_B_CY;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_B_XOR;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_C;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_C1;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_C2;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_C3;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_C4;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_C5;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_C6;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_CE;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_CLK;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_CO5;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_CO6;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_C_CY;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_C_XOR;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_D;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_D1;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_D2;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_D3;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_D4;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_D5;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_D6;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_DO5;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_DO6;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_D_CY;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_D_XOR;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X92Y112_SR;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_A;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_A1;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_A2;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_A3;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_A4;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_A5;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_A6;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_AO5;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_AO6;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_A_CY;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_A_XOR;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_B;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_B1;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_B2;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_B3;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_B4;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_B5;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_B6;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_BO5;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_BO6;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_B_CY;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_B_XOR;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_C;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_C1;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_C2;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_C3;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_C4;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_C5;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_C6;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_CO5;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_CO6;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_C_CY;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_C_XOR;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_D;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_D1;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_D2;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_D3;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_D4;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_D5;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_D6;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_DO5;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_DO6;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_D_CY;
  wire [0:0] CLBLM_L_X62Y112_SLICE_X93Y112_D_XOR;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_A;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_A1;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_A2;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_A3;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_A4;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_A5;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_A5Q;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_A6;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_AMUX;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_AO5;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_AO6;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_AQ;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_A_CY;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_A_XOR;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_B;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_B1;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_B2;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_B3;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_B4;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_B5;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_B6;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_BO5;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_BO6;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_B_CY;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_B_XOR;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_C;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_C1;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_C2;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_C3;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_C4;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_C5;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_C6;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_CE;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_CLK;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_CO5;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_CO6;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_C_CY;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_C_XOR;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_D;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_D1;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_D2;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_D3;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_D4;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_D5;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_D6;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_DO5;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_DO6;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_D_CY;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_D_XOR;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X92Y95_SR;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_A;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_A1;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_A2;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_A3;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_A4;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_A5;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_A6;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_AMUX;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_AO5;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_AO6;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_AQ;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_AX;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_A_CY;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_A_XOR;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_B;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_B1;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_B2;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_B3;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_B4;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_B5;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_B6;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_BMUX;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_BO5;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_BO6;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_BQ;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_BX;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_B_CY;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_B_XOR;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_C;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_C1;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_C2;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_C3;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_C4;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_C5;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_C6;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_CE;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_CLK;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_CO5;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_CO6;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_CQ;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_C_CY;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_C_XOR;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_D;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_D1;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_D2;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_D3;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_D4;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_D5;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_D5Q;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_D6;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_DMUX;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_DO5;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_DO6;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_DQ;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_D_CY;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_D_XOR;
  wire [0:0] CLBLM_L_X62Y95_SLICE_X93Y95_SR;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_A;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_A1;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_A2;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_A3;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_A4;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_A5;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_A6;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_AMUX;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_AO5;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_AO6;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_AX;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_A_CY;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_A_XOR;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_B;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_B1;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_B2;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_B3;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_B4;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_B5;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_B6;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_BO5;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_BO6;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_B_CY;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_B_XOR;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_C;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_C1;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_C2;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_C3;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_C4;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_C5;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_C6;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_CE;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_CLK;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_CO5;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_CO6;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_CQ;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_C_CY;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_C_XOR;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_D;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_D1;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_D2;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_D3;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_D4;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_D5;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_D6;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_DO5;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_DO6;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_D_CY;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_D_XOR;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_F7AMUX_O;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X92Y96_SR;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_A;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_A1;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_A2;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_A3;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_A4;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_A5;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_A6;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_AMUX;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_AO5;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_AO6;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_AX;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_A_CY;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_A_XOR;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_B;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_B1;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_B2;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_B3;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_B4;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_B5;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_B6;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_BO5;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_BO6;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_BQ;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_BX;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_B_CY;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_B_XOR;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_C;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_C1;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_C2;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_C3;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_C4;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_C5;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_C6;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_CE;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_CLK;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_CO5;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_CO6;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_CQ;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_C_CY;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_C_XOR;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_D;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_D1;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_D2;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_D3;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_D4;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_D5;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_D6;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_DO5;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_DO6;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_DQ;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_D_CY;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_D_XOR;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_F7AMUX_O;
  wire [0:0] CLBLM_L_X62Y96_SLICE_X93Y96_SR;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_A;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_A1;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_A2;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_A3;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_A4;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_A5;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_A6;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_AO5;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_AO6;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_AQ;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_A_CY;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_A_XOR;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_B;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_B1;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_B2;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_B3;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_B4;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_B5;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_B6;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_BO5;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_BO6;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_BQ;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_B_CY;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_B_XOR;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_C;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_C1;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_C2;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_C3;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_C4;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_C5;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_C5Q;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_C6;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_CE;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_CLK;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_CMUX;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_CO5;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_CO6;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_CQ;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_C_CY;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_C_XOR;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_D;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_D1;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_D2;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_D3;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_D4;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_D5;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_D5Q;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_D6;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_DMUX;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_DO5;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_DO6;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_DQ;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_DX;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_D_CY;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_D_XOR;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X92Y97_SR;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_A;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_A1;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_A2;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_A3;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_A4;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_A5;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_A6;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_AMUX;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_AO5;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_AO6;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_AX;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_A_CY;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_A_XOR;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_B;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_B1;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_B2;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_B3;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_B4;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_B5;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_B6;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_BO5;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_BO6;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_BQ;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_BX;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_B_CY;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_B_XOR;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_C;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_C1;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_C2;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_C3;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_C4;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_C5;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_C6;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_CE;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_CLK;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_CMUX;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_CO5;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_CO6;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_CQ;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_C_CY;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_C_XOR;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_D;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_D1;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_D2;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_D3;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_D4;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_D5;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_D6;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_DO5;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_DO6;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_DQ;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_DX;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_D_CY;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_D_XOR;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_F7AMUX_O;
  wire [0:0] CLBLM_L_X62Y97_SLICE_X93Y97_SR;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_A;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_A1;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_A2;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_A3;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_A4;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_A5;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_A6;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_AO5;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_AO6;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_AQ;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_A_CY;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_A_XOR;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_B;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_B1;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_B2;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_B3;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_B4;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_B5;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_B6;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_BO5;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_BO6;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_BQ;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_B_CY;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_B_XOR;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_C;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_C1;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_C2;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_C3;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_C4;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_C5;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_C6;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_CE;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_CLK;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_CO5;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_CO6;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_CQ;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_C_CY;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_C_XOR;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_D;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_D1;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_D2;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_D3;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_D4;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_D5;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_D6;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_DO5;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_DO6;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_DQ;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_D_CY;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_D_XOR;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X92Y98_SR;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_A;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_A1;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_A2;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_A3;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_A4;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_A5;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_A6;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_AO5;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_AO6;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_AQ;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_A_CY;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_A_XOR;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_B;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_B1;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_B2;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_B3;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_B4;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_B5;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_B6;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_BO5;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_BO6;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_BQ;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_B_CY;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_B_XOR;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_C;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_C1;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_C2;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_C3;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_C4;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_C5;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_C6;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_CLK;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_CO5;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_CO6;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_C_CY;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_C_XOR;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_D;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_D1;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_D2;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_D3;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_D4;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_D5;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_D6;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_DO5;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_DO6;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_D_CY;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_D_XOR;
  wire [0:0] CLBLM_L_X62Y98_SLICE_X93Y98_SR;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_A;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_A1;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_A2;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_A3;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_A4;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_A5;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_A6;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_AMUX;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_AO5;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_AO6;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_A_CY;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_A_XOR;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_B;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_B1;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_B2;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_B3;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_B4;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_B5;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_B6;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_BO5;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_BO6;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_BQ;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_B_CY;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_B_XOR;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_C;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_C1;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_C2;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_C3;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_C4;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_C5;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_C6;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_CLK;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_CO5;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_CO6;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_C_CY;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_C_XOR;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_D;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_D1;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_D2;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_D3;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_D4;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_D5;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_D6;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_DO5;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_DO6;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_D_CY;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_D_XOR;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X92Y99_SR;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_A;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_A1;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_A2;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_A3;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_A4;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_A5;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_A6;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_AO5;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_AO6;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_AQ;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_AX;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_A_CY;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_A_XOR;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_B;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_B1;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_B2;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_B3;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_B4;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_B5;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_B6;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_BMUX;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_BO5;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_BO6;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_B_CY;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_B_XOR;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_C;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_C1;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_C2;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_C3;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_C4;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_C5;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_C6;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_CE;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_CLK;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_CO5;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_CO6;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_C_CY;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_C_XOR;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_D;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_D1;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_D2;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_D3;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_D4;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_D5;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_D6;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_DO5;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_DO6;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_D_CY;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_D_XOR;
  wire [0:0] CLBLM_L_X62Y99_SLICE_X93Y99_SR;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_A;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_A1;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_A2;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_A3;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_A4;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_A5;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_A6;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_AMUX;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_AO5;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_AO6;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_AX;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_A_CY;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_A_XOR;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_B;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_B1;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_B2;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_B3;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_B4;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_B5;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_B6;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_BMUX;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_BO5;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_BO6;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_BX;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_B_CY;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_B_XOR;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_C;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_C1;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_C2;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_C3;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_C4;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_C5;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_C6;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_CMUX;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_CO5;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_CO6;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_COUT;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_CX;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_C_CY;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_C_XOR;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_D;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_D1;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_D2;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_D3;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_D4;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_D5;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_D6;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_DMUX;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_DO5;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_DO6;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_DX;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_D_CY;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X96Y100_D_XOR;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_A;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_A1;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_A2;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_A3;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_A4;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_A5;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_A6;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_AMUX;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_AO5;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_AO6;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_AQ;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_AX;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_A_CY;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_A_XOR;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_B;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_B1;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_B2;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_B3;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_B4;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_B5;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_B6;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_BMUX;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_BO5;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_BO6;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_BQ;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_BX;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_B_CY;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_B_XOR;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_C;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_C1;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_C2;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_C3;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_C4;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_C5;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_C6;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_CE;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_CLK;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_CMUX;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_CO5;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_CO6;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_COUT;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_CX;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_C_CY;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_C_XOR;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_D;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_D1;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_D2;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_D3;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_D4;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_D5;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_D6;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_DMUX;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_DO5;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_DO6;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_DX;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_D_CY;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_D_XOR;
  wire [0:0] CLBLM_L_X64Y100_SLICE_X97Y100_SR;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_A;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_A1;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_A2;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_A3;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_A4;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_A5;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_A6;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_AMUX;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_AO5;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_AO6;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_AX;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_A_CY;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_A_XOR;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_B;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_B1;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_B2;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_B3;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_B4;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_B5;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_B6;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_BMUX;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_BO5;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_BO6;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_BX;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_B_CY;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_B_XOR;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_C;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_C1;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_C2;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_C3;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_C4;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_C5;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_C6;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_CIN;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_CMUX;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_CO5;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_CO6;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_COUT;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_CX;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_C_CY;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_C_XOR;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_D;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_D1;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_D2;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_D3;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_D4;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_D5;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_D6;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_DMUX;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_DO5;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_DO6;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_DX;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_D_CY;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X96Y101_D_XOR;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_A;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_A1;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_A2;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_A3;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_A4;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_A5;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_A6;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_AMUX;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_AO5;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_AO6;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_AX;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_A_CY;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_A_XOR;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_B;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_B1;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_B2;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_B3;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_B4;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_B5;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_B6;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_BMUX;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_BO5;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_BO6;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_BX;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_B_CY;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_B_XOR;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_C;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_C1;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_C2;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_C3;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_C4;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_C5;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_C6;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_CIN;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_CMUX;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_CO5;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_CO6;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_COUT;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_CX;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_C_CY;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_C_XOR;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_D;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_D1;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_D2;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_D3;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_D4;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_D5;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_D6;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_DMUX;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_DO5;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_DO6;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_DX;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_D_CY;
  wire [0:0] CLBLM_L_X64Y101_SLICE_X97Y101_D_XOR;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_A;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_A1;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_A2;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_A3;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_A4;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_A5;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_A6;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_AMUX;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_AO5;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_AO6;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_AX;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_A_CY;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_A_XOR;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_B;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_B1;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_B2;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_B3;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_B4;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_B5;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_B6;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_BMUX;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_BO5;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_BO6;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_BX;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_B_CY;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_B_XOR;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_C;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_C1;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_C2;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_C3;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_C4;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_C5;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_C6;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_CIN;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_CMUX;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_CO5;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_CO6;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_COUT;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_CX;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_C_CY;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_C_XOR;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_D;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_D1;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_D2;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_D3;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_D4;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_D5;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_D6;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_DMUX;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_DO5;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_DO6;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_DX;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_D_CY;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X96Y102_D_XOR;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_A;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_A1;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_A2;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_A3;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_A4;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_A5;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_A6;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_AMUX;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_AO5;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_AO6;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_AQ;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_AX;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_A_CY;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_A_XOR;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_B;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_B1;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_B2;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_B3;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_B4;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_B5;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_B6;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_BMUX;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_BO5;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_BO6;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_BQ;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_BX;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_B_CY;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_B_XOR;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_C;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_C1;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_C2;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_C3;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_C4;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_C5;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_C6;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_CE;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_CIN;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_CLK;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_CMUX;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_CO5;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_CO6;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_COUT;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_CQ;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_CX;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_C_CY;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_C_XOR;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_D;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_D1;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_D2;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_D3;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_D4;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_D5;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_D6;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_DMUX;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_DO5;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_DO6;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_D_CY;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_D_XOR;
  wire [0:0] CLBLM_L_X64Y102_SLICE_X97Y102_SR;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_A;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_A1;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_A2;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_A3;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_A4;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_A5;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_A6;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_AMUX;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_AO5;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_AO6;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_AX;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_A_CY;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_A_XOR;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_B;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_B1;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_B2;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_B3;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_B4;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_B5;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_B6;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_BMUX;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_BO5;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_BO6;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_BX;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_B_CY;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_B_XOR;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_C;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_C1;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_C2;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_C3;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_C4;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_C5;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_C6;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_CIN;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_CMUX;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_CO5;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_CO6;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_COUT;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_CX;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_C_CY;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_C_XOR;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_D;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_D1;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_D2;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_D3;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_D4;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_D5;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_D6;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_DMUX;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_DO5;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_DO6;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_DX;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_D_CY;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X96Y103_D_XOR;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_A;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_A1;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_A2;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_A3;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_A4;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_A5;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_A6;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_AMUX;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_AO5;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_AO6;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_AX;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_A_CY;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_A_XOR;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_B;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_B1;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_B2;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_B3;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_B4;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_B5;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_B6;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_BMUX;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_BO5;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_BO6;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_BX;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_B_CY;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_B_XOR;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_C;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_C1;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_C2;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_C3;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_C4;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_C5;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_C6;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_CIN;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_CMUX;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_CO5;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_CO6;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_COUT;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_CX;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_C_CY;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_C_XOR;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_D;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_D1;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_D2;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_D3;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_D4;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_D5;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_D6;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_DMUX;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_DO5;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_DO6;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_DX;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_D_CY;
  wire [0:0] CLBLM_L_X64Y103_SLICE_X97Y103_D_XOR;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_A;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_A1;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_A2;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_A3;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_A4;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_A5;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_A6;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_AMUX;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_AO5;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_AO6;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_AX;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_A_CY;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_A_XOR;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_B;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_B1;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_B2;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_B3;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_B4;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_B5;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_B6;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_BMUX;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_BO5;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_BO6;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_BX;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_B_CY;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_B_XOR;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_C;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_C1;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_C2;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_C3;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_C4;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_C5;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_C6;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_CIN;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_CO5;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_CO6;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_COUT;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_CX;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_C_CY;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_C_XOR;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_D;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_D1;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_D2;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_D3;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_D4;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_D5;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_D6;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_DO5;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_DO6;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_DX;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_D_CY;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X96Y104_D_XOR;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_A;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_A1;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_A2;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_A3;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_A4;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_A5;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_A6;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_AMUX;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_AO5;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_AO6;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_AX;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_A_CY;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_A_XOR;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_B;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_B1;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_B2;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_B3;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_B4;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_B5;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_B6;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_BMUX;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_BO5;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_BO6;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_BX;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_B_CY;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_B_XOR;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_C;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_C1;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_C2;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_C3;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_C4;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_C5;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_C6;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_CIN;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_CMUX;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_CO5;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_CO6;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_COUT;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_CX;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_C_CY;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_C_XOR;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_D;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_D1;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_D2;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_D3;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_D4;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_D5;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_D6;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_DO5;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_DO6;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_DX;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_D_CY;
  wire [0:0] CLBLM_L_X64Y104_SLICE_X97Y104_D_XOR;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_A;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_A1;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_A2;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_A3;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_A4;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_A5;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_A6;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_AO5;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_AO6;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_AQ;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_A_CY;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_A_XOR;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_B;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_B1;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_B2;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_B3;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_B4;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_B5;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_B6;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_BO5;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_BO6;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_B_CY;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_B_XOR;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_C;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_C1;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_C2;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_C3;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_C4;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_C5;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_C6;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_CE;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_CLK;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_CO5;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_CO6;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_C_CY;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_C_XOR;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_D;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_D1;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_D2;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_D3;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_D4;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_D5;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_D6;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_DO5;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_DO6;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_D_CY;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_D_XOR;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X96Y105_SR;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_A;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_A1;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_A2;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_A3;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_A4;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_A5;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_A6;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_AO5;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_AO6;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_AQ;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_A_CY;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_A_XOR;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_B;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_B1;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_B2;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_B3;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_B4;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_B5;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_B6;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_BO5;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_BO6;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_B_CY;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_B_XOR;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_C;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_C1;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_C2;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_C3;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_C4;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_C5;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_C6;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_CE;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_CLK;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_CO5;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_CO6;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_C_CY;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_C_XOR;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_D;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_D1;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_D2;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_D3;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_D4;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_D5;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_D6;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_DMUX;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_DO5;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_DO6;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_D_CY;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_D_XOR;
  wire [0:0] CLBLM_L_X64Y105_SLICE_X97Y105_SR;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_A;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_A1;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_A2;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_A3;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_A4;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_A5;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_A6;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_AO5;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_AO6;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_AQ;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_A_CY;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_A_XOR;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_B;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_B1;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_B2;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_B3;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_B4;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_B5;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_B6;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_BO5;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_BO6;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_BQ;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_B_CY;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_B_XOR;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_C;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_C1;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_C2;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_C3;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_C4;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_C5;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_C6;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_CE;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_CLK;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_CO5;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_CO6;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_C_CY;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_C_XOR;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_D;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_D1;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_D2;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_D3;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_D4;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_D5;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_D6;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_DMUX;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_DO5;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_DO6;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_D_CY;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_D_XOR;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X96Y106_SR;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_A;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_A1;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_A2;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_A3;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_A4;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_A5;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_A6;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_AO5;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_AO6;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_AQ;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_A_CY;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_A_XOR;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_B;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_B1;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_B2;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_B3;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_B4;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_B5;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_B6;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_BO5;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_BO6;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_BQ;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_B_CY;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_B_XOR;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_C;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_C1;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_C2;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_C3;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_C4;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_C5;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_C6;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_CE;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_CLK;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_CO5;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_CO6;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_CQ;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_C_CY;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_C_XOR;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_D;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_D1;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_D2;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_D3;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_D4;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_D5;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_D6;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_DO5;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_DO6;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_DQ;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_D_CY;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_D_XOR;
  wire [0:0] CLBLM_L_X64Y106_SLICE_X97Y106_SR;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_A;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_A1;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_A2;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_A3;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_A4;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_A5;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_A6;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_AO5;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_AO6;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_AQ;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_A_CY;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_A_XOR;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_B;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_B1;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_B2;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_B3;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_B4;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_B5;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_B6;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_BO5;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_BO6;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_BQ;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_B_CY;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_B_XOR;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_C;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_C1;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_C2;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_C3;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_C4;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_C5;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_C6;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_CE;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_CLK;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_CO5;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_CO6;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_C_CY;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_C_XOR;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_D;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_D1;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_D2;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_D3;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_D4;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_D5;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_D6;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_DO5;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_DO6;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_D_CY;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_D_XOR;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X96Y107_SR;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_A;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_A1;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_A2;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_A3;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_A4;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_A5;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_A6;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_AO5;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_AO6;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_AQ;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_A_CY;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_A_XOR;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_B;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_B1;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_B2;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_B3;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_B4;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_B5;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_B6;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_BO5;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_BO6;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_BQ;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_B_CY;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_B_XOR;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_C;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_C1;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_C2;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_C3;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_C4;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_C5;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_C6;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_CE;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_CLK;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_CO5;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_CO6;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_C_CY;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_C_XOR;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_D;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_D1;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_D2;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_D3;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_D4;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_D5;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_D6;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_DMUX;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_DO5;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_DO6;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_D_CY;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_D_XOR;
  wire [0:0] CLBLM_L_X64Y107_SLICE_X97Y107_SR;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_A;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_A1;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_A2;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_A3;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_A4;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_A5;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_A6;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_AO5;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_AO6;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_AQ;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_A_CY;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_A_XOR;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_B;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_B1;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_B2;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_B3;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_B4;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_B5;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_B6;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_BO5;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_BO6;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_BQ;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_B_CY;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_B_XOR;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_C;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_C1;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_C2;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_C3;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_C4;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_C5;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_C6;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_CE;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_CLK;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_CO5;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_CO6;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_C_CY;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_C_XOR;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_D;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_D1;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_D2;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_D3;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_D4;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_D5;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_D6;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_DO5;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_DO6;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_D_CY;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_D_XOR;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X96Y108_SR;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_A;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_A1;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_A2;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_A3;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_A4;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_A5;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_A6;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_AO5;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_AO6;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_AQ;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_A_CY;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_A_XOR;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_B;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_B1;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_B2;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_B3;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_B4;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_B5;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_B6;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_BO5;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_BO6;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_B_CY;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_B_XOR;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_C;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_C1;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_C2;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_C3;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_C4;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_C5;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_C6;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_CE;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_CLK;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_CO5;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_CO6;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_C_CY;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_C_XOR;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_D;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_D1;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_D2;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_D3;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_D4;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_D5;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_D6;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_DO5;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_DO6;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_D_CY;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_D_XOR;
  wire [0:0] CLBLM_L_X64Y108_SLICE_X97Y108_SR;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_A;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_A1;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_A2;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_A3;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_A4;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_A5;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_A5Q;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_A6;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_AMUX;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_AO5;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_AO6;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_AQ;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_A_CY;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_A_XOR;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_B;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_B1;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_B2;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_B3;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_B4;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_B5;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_B6;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_BO5;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_BO6;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_B_CY;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_B_XOR;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_C;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_C1;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_C2;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_C3;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_C4;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_C5;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_C6;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_CE;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_CLK;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_CO5;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_CO6;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_C_CY;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_C_XOR;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_D;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_D1;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_D2;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_D3;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_D4;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_D5;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_D6;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_DO5;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_DO6;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_D_CY;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_D_XOR;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X96Y109_SR;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_A;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_A1;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_A2;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_A3;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_A4;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_A5;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_A6;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_AO5;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_AO6;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_A_CY;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_A_XOR;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_B;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_B1;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_B2;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_B3;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_B4;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_B5;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_B6;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_BO5;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_BO6;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_B_CY;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_B_XOR;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_C;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_C1;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_C2;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_C3;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_C4;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_C5;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_C6;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_CO5;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_CO6;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_C_CY;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_C_XOR;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_D;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_D1;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_D2;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_D3;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_D4;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_D5;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_D6;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_DO5;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_DO6;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_D_CY;
  wire [0:0] CLBLM_L_X64Y109_SLICE_X97Y109_D_XOR;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_A;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_A1;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_A2;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_A3;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_A4;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_A5;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_A6;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_AI;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_AMUX;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_AO5;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_AO6;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_AX;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_B;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_B1;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_B2;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_B3;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_B4;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_B5;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_B6;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_BI;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_BMUX;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_BO5;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_BO6;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_BX;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_C;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_C1;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_C2;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_C3;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_C4;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_C5;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_C6;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_CE;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_CI;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_CLK;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_CMUX;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_CO5;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_CO6;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_CX;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_D;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_D1;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_D2;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_D3;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_D4;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_D5;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_D6;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_DI;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_DO5;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_DO6;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X96Y95_DX;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_A;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_A1;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_A2;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_A3;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_A4;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_A5;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_A6;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_AO5;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_AO6;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_A_CY;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_A_XOR;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_B;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_B1;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_B2;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_B3;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_B4;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_B5;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_B6;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_BO5;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_BO6;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_B_CY;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_B_XOR;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_C;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_C1;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_C2;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_C3;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_C4;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_C5;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_C6;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_CO5;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_CO6;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_C_CY;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_C_XOR;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_D;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_D1;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_D2;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_D3;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_D4;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_D5;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_D6;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_DO5;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_DO6;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_D_CY;
  wire [0:0] CLBLM_L_X64Y95_SLICE_X97Y95_D_XOR;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_A;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_A1;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_A2;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_A3;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_A4;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_A5;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_A6;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_AI;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_AMUX;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_AO5;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_AO6;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_AX;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_B;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_B1;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_B2;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_B3;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_B4;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_B5;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_B6;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_BI;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_BMUX;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_BO5;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_BO6;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_BX;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_C;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_C1;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_C2;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_C3;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_C4;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_C5;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_C6;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_CE;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_CI;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_CLK;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_CMUX;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_CO5;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_CO6;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_CX;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_D;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_D1;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_D2;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_D3;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_D4;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_D5;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_D6;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_DI;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_DO5;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_DO6;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X96Y96_DX;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_A;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_A1;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_A2;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_A3;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_A4;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_A5;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_A6;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_AO5;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_AO6;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_AQ;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_A_CY;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_A_XOR;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_B;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_B1;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_B2;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_B3;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_B4;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_B5;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_B6;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_BO5;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_BO6;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_BQ;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_B_CY;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_B_XOR;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_C;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_C1;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_C2;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_C3;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_C4;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_C5;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_C6;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_CE;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_CLK;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_CO5;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_CO6;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_CQ;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_C_CY;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_C_XOR;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_D;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_D1;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_D2;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_D3;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_D4;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_D5;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_D6;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_DO5;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_DO6;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_DQ;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_D_CY;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_D_XOR;
  wire [0:0] CLBLM_L_X64Y96_SLICE_X97Y96_SR;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_A;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_A1;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_A2;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_A3;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_A4;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_A5;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_A5Q;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_A6;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_AMUX;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_AO5;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_AO6;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_AQ;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_A_CY;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_A_XOR;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_B;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_B1;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_B2;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_B3;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_B4;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_B5;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_B5Q;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_B6;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_BMUX;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_BO5;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_BO6;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_BQ;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_B_CY;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_B_XOR;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_C;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_C1;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_C2;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_C3;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_C4;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_C5;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_C6;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_CE;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_CLK;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_CO5;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_CO6;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_C_CY;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_C_XOR;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_D;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_D1;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_D2;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_D3;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_D4;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_D5;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_D6;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_DO5;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_DO6;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_D_CY;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_D_XOR;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X96Y97_SR;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_A;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_A1;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_A2;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_A3;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_A4;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_A5;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_A6;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_AO5;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_AO6;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_AQ;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_A_CY;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_A_XOR;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_B;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_B1;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_B2;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_B3;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_B4;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_B5;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_B6;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_BO5;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_BO6;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_BQ;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_B_CY;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_B_XOR;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_C;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_C1;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_C2;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_C3;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_C4;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_C5;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_C6;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_CE;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_CLK;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_CMUX;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_CO5;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_CO6;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_C_CY;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_C_XOR;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_D;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_D1;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_D2;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_D3;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_D4;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_D5;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_D6;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_DO5;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_DO6;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_D_CY;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_D_XOR;
  wire [0:0] CLBLM_L_X64Y97_SLICE_X97Y97_SR;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_A;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_A1;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_A2;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_A3;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_A4;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_A5;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_A6;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_AO5;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_AO6;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_AQ;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_A_CY;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_A_XOR;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_B;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_B1;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_B2;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_B3;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_B4;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_B5;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_B6;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_BO5;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_BO6;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_B_CY;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_B_XOR;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_C;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_C1;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_C2;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_C3;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_C4;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_C5;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_C6;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_CE;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_CLK;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_CO5;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_CO6;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_C_CY;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_C_XOR;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_D;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_D1;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_D2;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_D3;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_D4;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_D5;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_D6;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_DO5;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_DO6;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_D_CY;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_D_XOR;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X96Y98_SR;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_A;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_A1;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_A2;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_A3;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_A4;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_A5;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_A6;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_AO5;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_AO6;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_AQ;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_A_CY;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_A_XOR;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_B;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_B1;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_B2;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_B3;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_B4;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_B5;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_B6;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_BO5;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_BO6;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_B_CY;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_B_XOR;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_C;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_C1;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_C2;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_C3;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_C4;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_C5;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_C6;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_CE;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_CLK;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_CO5;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_CO6;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_C_CY;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_C_XOR;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_D;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_D1;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_D2;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_D3;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_D4;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_D5;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_D6;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_DO5;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_DO6;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_D_CY;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_D_XOR;
  wire [0:0] CLBLM_L_X64Y98_SLICE_X97Y98_SR;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_A;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_A1;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_A2;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_A3;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_A4;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_A5;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_A6;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_AO5;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_AO6;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_AQ;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_A_CY;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_A_XOR;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_B;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_B1;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_B2;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_B3;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_B4;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_B5;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_B6;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_BO5;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_BO6;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_BQ;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_B_CY;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_B_XOR;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_C;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_C1;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_C2;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_C3;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_C4;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_C5;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_C6;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_CE;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_CLK;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_CO5;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_CO6;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_C_CY;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_C_XOR;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_D;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_D1;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_D2;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_D3;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_D4;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_D5;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_D6;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_DO5;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_DO6;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_D_CY;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_D_XOR;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X96Y99_SR;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_A;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_A1;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_A2;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_A3;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_A4;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_A5;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_A6;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_AO5;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_AO6;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_AQ;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_A_CY;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_A_XOR;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_B;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_B1;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_B2;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_B3;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_B4;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_B5;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_B6;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_BO5;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_BO6;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_B_CY;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_B_XOR;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_C;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_C1;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_C2;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_C3;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_C4;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_C5;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_C6;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_CE;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_CLK;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_CO5;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_CO6;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_C_CY;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_C_XOR;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_D;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_D1;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_D2;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_D3;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_D4;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_D5;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_D6;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_DO5;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_DO6;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_D_CY;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_D_XOR;
  wire [0:0] CLBLM_L_X64Y99_SLICE_X97Y99_SR;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_A;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_A1;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_A2;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_A3;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_A4;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_A5;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_A6;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_AO5;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_AO6;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_A_CY;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_A_XOR;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_B;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_B1;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_B2;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_B3;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_B4;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_B5;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_B6;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_BO5;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_BO6;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_B_CY;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_B_XOR;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_C;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_C1;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_C2;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_C3;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_C4;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_C5;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_C6;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_CO5;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_CO6;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_C_CY;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_C_XOR;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_D;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_D1;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_D2;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_D3;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_D4;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_D5;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_D6;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_DO5;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_DO6;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_D_CY;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_D_XOR;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_A;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_A1;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_A2;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_A3;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_A4;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_A5;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_A6;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_AO5;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_AO6;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_A_CY;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_A_XOR;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_B;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_B1;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_B2;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_B3;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_B4;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_B5;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_B6;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_BO5;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_BO6;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_B_CY;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_B_XOR;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_C;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_C1;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_C2;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_C3;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_C4;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_C5;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_C6;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_CO5;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_CO6;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_C_CY;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_C_XOR;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_D;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_D1;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_D2;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_D3;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_D4;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_D5;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_D6;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_DO5;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_DO6;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_D_CY;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_D_XOR;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_A;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_A1;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_A2;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_A3;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_A4;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_A5;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_A6;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_AO5;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_AO6;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_A_CY;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_A_XOR;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_B;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_B1;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_B2;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_B3;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_B4;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_B5;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_B6;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_BO5;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_BO6;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_B_CY;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_B_XOR;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_C;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_C1;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_C2;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_C3;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_C4;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_C5;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_C6;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_CO5;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_CO6;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_C_CY;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_C_XOR;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_D;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_D1;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_D2;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_D3;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_D4;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_D5;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_D6;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_DO5;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_DO6;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_D_CY;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X72Y119_D_XOR;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_A;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_A1;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_A2;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_A3;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_A4;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_A5;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_A6;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_AMUX;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_AO5;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_AO6;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_AQ;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_AX;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_A_CY;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_A_XOR;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_B;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_B1;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_B2;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_B3;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_B4;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_B5;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_B6;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_BO5;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_BO6;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_BQ;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_BX;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_B_CY;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_B_XOR;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_C;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_C1;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_C2;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_C3;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_C4;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_C5;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_C6;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_CLK;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_CO5;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_CO6;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_CQ;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_CX;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_C_CY;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_C_XOR;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_D;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_D1;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_D2;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_D3;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_D4;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_D5;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_D6;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_DO5;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_DO6;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_DQ;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_DX;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_D_CY;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_D_XOR;
  wire [0:0] CLBLM_R_X47Y119_SLICE_X73Y119_SR;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_A;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_A1;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_A2;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_A3;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_A4;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_A5;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_A6;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_AO5;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_AO6;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_AQ;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_AX;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_A_CY;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_A_XOR;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_B;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_B1;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_B2;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_B3;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_B4;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_B5;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_B6;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_BO5;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_BO6;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_BX;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_B_CY;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_B_XOR;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_C;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_C1;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_C2;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_C3;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_C4;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_C5;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_C6;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_CE;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_CLK;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_CO5;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_CO6;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_C_CY;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_C_XOR;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_D;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_D1;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_D2;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_D3;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_D4;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_D5;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_D6;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_DO5;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_DO6;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_D_CY;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_D_XOR;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X74Y104_SR;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_A;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_A1;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_A2;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_A3;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_A4;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_A5;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_A6;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_AO5;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_AO6;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_AQ;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_AX;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_A_CY;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_A_XOR;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_B;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_B1;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_B2;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_B3;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_B4;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_B5;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_B6;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_BO5;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_BO6;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_BQ;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_BX;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_B_CY;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_B_XOR;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_C;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_C1;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_C2;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_C3;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_C4;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_C5;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_C6;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_CE;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_CLK;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_CO5;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_CO6;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_CQ;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_CX;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_C_CY;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_C_XOR;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_D;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_D1;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_D2;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_D3;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_D4;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_D5;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_D6;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_DO5;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_DO6;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_DQ;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_DX;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_D_CY;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_D_XOR;
  wire [0:0] CLBLM_R_X49Y104_SLICE_X75Y104_SR;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_A;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_A1;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_A2;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_A3;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_A4;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_A5;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_A6;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_AO5;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_AO6;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_A_CY;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_A_XOR;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_B;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_B1;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_B2;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_B3;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_B4;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_B5;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_B6;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_BO5;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_BO6;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_B_CY;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_B_XOR;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_C;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_C1;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_C2;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_C3;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_C4;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_C5;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_C6;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_CO5;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_CO6;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_C_CY;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_C_XOR;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_D;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_D1;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_D2;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_D3;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_D4;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_D5;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_D6;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_DO5;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_DO6;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_D_CY;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X74Y105_D_XOR;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_A;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_A1;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_A2;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_A3;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_A4;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_A5;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_A6;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_AMUX;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_AO5;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_AO6;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_AX;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_A_CY;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_A_XOR;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_B;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_B1;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_B2;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_B3;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_B4;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_B5;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_B6;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_BO5;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_BO6;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_B_CY;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_B_XOR;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_C;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_C1;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_C2;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_C3;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_C4;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_C5;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_C6;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_CE;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_CLK;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_CO5;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_CO6;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_CQ;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_C_CY;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_C_XOR;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_D;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_D1;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_D2;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_D3;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_D4;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_D5;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_D6;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_DO5;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_DO6;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_D_CY;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_D_XOR;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_F7AMUX_O;
  wire [0:0] CLBLM_R_X49Y105_SLICE_X75Y105_SR;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_A;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_A1;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_A2;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_A3;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_A4;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_A5;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_A6;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_AO5;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_AO6;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_AQ;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_A_CY;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_A_XOR;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_B;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_B1;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_B2;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_B3;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_B4;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_B5;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_B6;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_BO5;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_BO6;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_B_CY;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_B_XOR;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_C;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_C1;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_C2;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_C3;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_C4;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_C5;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_C6;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_CE;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_CLK;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_CMUX;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_CO5;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_CO6;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_C_CY;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_C_XOR;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_D;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_D1;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_D2;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_D3;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_D4;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_D5;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_D6;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_DO5;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_DO6;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_D_CY;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_D_XOR;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X74Y106_SR;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_A;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_A1;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_A2;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_A3;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_A4;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_A5;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_A6;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_AMUX;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_AO5;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_AO6;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_AX;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_A_CY;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_A_XOR;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_B;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_B1;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_B2;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_B3;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_B4;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_B5;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_B6;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_BO5;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_BO6;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_BX;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_B_CY;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_B_XOR;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_C;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_C1;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_C2;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_C3;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_C4;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_C5;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_C6;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_CE;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_CLK;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_CO5;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_CO6;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_CQ;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_CX;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_C_CY;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_C_XOR;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_D;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_D1;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_D2;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_D3;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_D4;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_D5;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_D6;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_DMUX;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_DO5;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_DO6;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_DQ;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_DX;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_D_CY;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_D_XOR;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_F7AMUX_O;
  wire [0:0] CLBLM_R_X49Y106_SLICE_X75Y106_SR;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_A;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_A1;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_A2;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_A3;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_A4;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_A5;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_A6;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_AO5;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_AO6;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_AQ;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_A_CY;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_A_XOR;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_B;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_B1;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_B2;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_B3;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_B4;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_B5;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_B6;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_BO5;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_BO6;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_B_CY;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_B_XOR;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_C;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_C1;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_C2;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_C3;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_C4;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_C5;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_C6;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_CE;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_CLK;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_CO5;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_CO6;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_C_CY;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_C_XOR;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_D;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_D1;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_D2;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_D3;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_D4;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_D5;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_D6;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_DO5;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_DO6;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_D_CY;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_D_XOR;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X74Y107_SR;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_A;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_A1;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_A2;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_A3;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_A4;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_A5;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_A6;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_AMUX;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_AO5;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_AO6;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_AX;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_A_CY;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_A_XOR;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_B;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_B1;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_B2;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_B3;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_B4;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_B5;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_B6;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_BO5;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_BO6;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_BX;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_B_CY;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_B_XOR;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_C;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_C1;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_C2;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_C3;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_C4;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_C5;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_C6;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_CE;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_CLK;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_CMUX;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_CO5;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_CO6;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_CQ;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_CX;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_C_CY;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_C_XOR;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_D;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_D1;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_D2;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_D3;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_D4;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_D5;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_D6;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_DO5;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_DO6;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_DQ;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_DX;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_D_CY;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_D_XOR;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_F7AMUX_O;
  wire [0:0] CLBLM_R_X49Y107_SLICE_X75Y107_SR;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_A;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_A1;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_A2;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_A3;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_A4;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_A5;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_A5Q;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_A6;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_AMUX;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_AO5;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_AO6;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_AQ;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_A_CY;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_A_XOR;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_B;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_B1;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_B2;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_B3;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_B4;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_B5;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_B5Q;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_B6;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_BMUX;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_BO5;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_BO6;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_BQ;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_B_CY;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_B_XOR;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_C;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_C1;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_C2;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_C3;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_C4;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_C5;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_C5Q;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_C6;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_CE;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_CLK;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_CMUX;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_CO5;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_CO6;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_CQ;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_C_CY;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_C_XOR;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_D;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_D1;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_D2;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_D3;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_D4;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_D5;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_D6;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_DO5;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_DO6;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_D_CY;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_D_XOR;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X74Y108_SR;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_A;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_A1;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_A2;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_A3;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_A4;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_A5;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_A6;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_AMUX;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_AO5;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_AO6;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_AX;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_A_CY;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_A_XOR;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_B;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_B1;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_B2;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_B3;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_B4;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_B5;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_B6;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_BMUX;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_BO5;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_BO6;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_BX;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_B_CY;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_B_XOR;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_C;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_C1;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_C2;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_C3;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_C4;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_C5;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_C6;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_CE;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_CLK;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_CMUX;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_CO5;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_CO6;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_COUT;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_CX;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_C_CY;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_C_XOR;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_D;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_D1;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_D2;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_D3;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_D4;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_D5;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_D6;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_DMUX;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_DO5;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_DO6;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_DQ;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_DX;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_D_CY;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_D_XOR;
  wire [0:0] CLBLM_R_X49Y108_SLICE_X75Y108_SR;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_A;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_A1;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_A2;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_A3;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_A4;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_A5;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_A6;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_AO5;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_AO6;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_AQ;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_A_CY;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_A_XOR;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_B;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_B1;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_B2;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_B3;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_B4;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_B5;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_B6;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_BO5;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_BO6;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_BQ;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_B_CY;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_B_XOR;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_C;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_C1;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_C2;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_C3;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_C4;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_C5;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_C6;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_CE;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_CLK;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_CO5;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_CO6;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_CQ;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_C_CY;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_C_XOR;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_D;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_D1;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_D2;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_D3;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_D4;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_D5;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_D6;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_DO5;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_DO6;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_DQ;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_D_CY;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_D_XOR;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X74Y109_SR;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_A;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_A1;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_A2;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_A3;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_A4;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_A5;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_A6;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_AMUX;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_AO5;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_AO6;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_AX;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_A_CY;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_A_XOR;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_B;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_B1;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_B2;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_B3;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_B4;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_B5;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_B6;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_BMUX;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_BO5;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_BO6;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_BX;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_B_CY;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_B_XOR;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_C;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_C1;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_C2;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_C3;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_C4;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_C5;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_C6;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_CIN;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_CMUX;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_CO5;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_CO6;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_COUT;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_CX;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_C_CY;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_C_XOR;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_D;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_D1;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_D2;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_D3;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_D4;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_D5;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_D6;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_DMUX;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_DO5;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_DO6;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_DX;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_D_CY;
  wire [0:0] CLBLM_R_X49Y109_SLICE_X75Y109_D_XOR;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_A;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_A1;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_A2;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_A3;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_A4;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_A5;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_A5Q;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_A6;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_AMUX;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_AO5;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_AO6;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_AQ;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_A_CY;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_A_XOR;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_B;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_B1;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_B2;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_B3;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_B4;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_B5;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_B6;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_BO5;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_BO6;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_B_CY;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_B_XOR;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_C;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_C1;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_C2;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_C3;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_C4;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_C5;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_C6;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_CE;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_CLK;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_CO5;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_CO6;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_C_CY;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_C_XOR;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_D;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_D1;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_D2;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_D3;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_D4;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_D5;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_D6;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_DO5;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_DO6;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_D_CY;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_D_XOR;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X74Y110_SR;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_A;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_A1;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_A2;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_A3;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_A4;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_A5;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_A6;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_AMUX;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_AO5;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_AO6;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_AX;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_A_CY;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_A_XOR;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_B;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_B1;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_B2;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_B3;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_B4;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_B5;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_B6;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_BO5;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_BO6;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_BX;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_B_CY;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_B_XOR;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_C;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_C1;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_C2;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_C3;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_C4;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_C5;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_C6;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_CIN;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_CO5;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_CO6;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_COUT;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_CX;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_C_CY;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_C_XOR;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_D;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_D1;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_D2;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_D3;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_D4;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_D5;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_D6;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_DO5;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_DO6;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_DX;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_D_CY;
  wire [0:0] CLBLM_R_X49Y110_SLICE_X75Y110_D_XOR;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_A;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_A1;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_A2;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_A3;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_A4;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_A5;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_A6;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_AO5;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_AO6;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_AQ;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_A_CY;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_A_XOR;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_B;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_B1;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_B2;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_B3;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_B4;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_B5;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_B6;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_BO5;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_BO6;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_BQ;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_B_CY;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_B_XOR;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_C;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_C1;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_C2;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_C3;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_C4;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_C5;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_C6;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_CE;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_CLK;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_CO5;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_CO6;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_CQ;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_C_CY;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_C_XOR;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_D;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_D1;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_D2;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_D3;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_D4;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_D5;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_D6;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_DO5;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_DO6;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_D_CY;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_D_XOR;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X74Y111_SR;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_A;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_A1;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_A2;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_A3;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_A4;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_A5;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_A5Q;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_A6;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_AMUX;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_AO5;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_AO6;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_AQ;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_A_CY;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_A_XOR;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_B;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_B1;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_B2;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_B3;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_B4;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_B5;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_B6;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_BMUX;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_BO5;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_BO6;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_B_CY;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_B_XOR;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_C;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_C1;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_C2;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_C3;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_C4;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_C5;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_C6;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_CE;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_CLK;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_CO5;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_CO6;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_C_CY;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_C_XOR;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_D;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_D1;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_D2;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_D3;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_D4;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_D5;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_D6;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_DO5;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_DO6;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_D_CY;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_D_XOR;
  wire [0:0] CLBLM_R_X49Y111_SLICE_X75Y111_SR;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_A;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_A1;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_A2;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_A3;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_A4;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_A5;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_A6;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_AO5;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_AO6;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_AQ;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_A_CY;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_A_XOR;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_B;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_B1;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_B2;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_B3;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_B4;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_B5;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_B6;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_BO5;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_BO6;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_BQ;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_B_CY;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_B_XOR;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_C;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_C1;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_C2;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_C3;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_C4;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_C5;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_C6;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_CLK;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_CO5;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_CO6;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_C_CY;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_C_XOR;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_D;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_D1;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_D2;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_D3;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_D4;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_D5;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_D6;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_DO5;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_DO6;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_D_CY;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_D_XOR;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X74Y119_SR;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_A;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_A1;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_A2;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_A3;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_A4;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_A5;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_A6;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_AO5;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_AO6;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_A_CY;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_A_XOR;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_B;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_B1;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_B2;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_B3;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_B4;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_B5;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_B6;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_BO5;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_BO6;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_B_CY;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_B_XOR;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_C;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_C1;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_C2;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_C3;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_C4;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_C5;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_C6;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_CO5;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_CO6;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_C_CY;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_C_XOR;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_D;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_D1;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_D2;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_D3;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_D4;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_D5;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_D6;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_DO5;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_DO6;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_D_CY;
  wire [0:0] CLBLM_R_X49Y119_SLICE_X75Y119_D_XOR;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_A;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_A1;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_A2;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_A3;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_A4;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_A5;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_A5Q;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_A6;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_AMUX;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_AO5;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_AO6;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_AQ;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_A_CY;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_A_XOR;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_B;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_B1;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_B2;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_B3;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_B4;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_B5;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_B6;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_BMUX;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_BO5;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_BO6;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_B_CY;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_B_XOR;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_C;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_C1;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_C2;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_C3;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_C4;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_C5;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_C6;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_CE;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_CLK;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_CMUX;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_CO5;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_CO6;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_C_CY;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_C_XOR;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_D;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_D1;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_D2;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_D3;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_D4;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_D5;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_D6;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_DO5;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_DO6;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_D_CY;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_D_XOR;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X80Y100_SR;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_A;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_A1;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_A2;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_A3;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_A4;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_A5;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_A6;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_AMUX;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_AO5;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_AO6;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_AQ;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_A_CY;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_A_XOR;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_B;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_B1;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_B2;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_B3;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_B4;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_B5;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_B6;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_BO5;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_BO6;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_B_CY;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_B_XOR;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_C;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_C1;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_C2;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_C3;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_C4;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_C5;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_C6;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_CE;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_CLK;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_CO5;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_CO6;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_C_CY;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_C_XOR;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_D;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_D1;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_D2;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_D3;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_D4;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_D5;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_D6;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_DO5;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_DO6;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_D_CY;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_D_XOR;
  wire [0:0] CLBLM_R_X53Y100_SLICE_X81Y100_SR;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_A;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_A1;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_A2;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_A3;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_A4;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_A5;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_A6;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_AMUX;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_AO5;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_AO6;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_A_CY;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_A_XOR;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_B;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_B1;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_B2;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_B3;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_B4;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_B5;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_B6;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_BO5;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_BO6;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_BQ;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_B_CY;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_B_XOR;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_C;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_C1;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_C2;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_C3;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_C4;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_C5;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_C6;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_CE;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_CLK;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_CO5;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_CO6;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_C_CY;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_C_XOR;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_D;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_D1;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_D2;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_D3;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_D4;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_D5;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_D6;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_DO5;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_DO6;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_D_CY;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_D_XOR;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X80Y101_SR;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_A;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_A1;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_A2;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_A3;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_A4;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_A5;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_A6;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_AO5;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_AO6;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_AQ;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_A_CY;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_A_XOR;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_B;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_B1;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_B2;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_B3;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_B4;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_B5;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_B6;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_BMUX;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_BO5;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_BO6;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_B_CY;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_B_XOR;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_C;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_C1;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_C2;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_C3;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_C4;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_C5;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_C6;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_CE;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_CLK;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_CO5;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_CO6;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_C_CY;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_C_XOR;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_D;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_D1;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_D2;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_D3;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_D4;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_D5;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_D6;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_DO5;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_DO6;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_D_CY;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_D_XOR;
  wire [0:0] CLBLM_R_X53Y101_SLICE_X81Y101_SR;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_A;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_A1;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_A2;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_A3;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_A4;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_A5;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_A6;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_AO5;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_AO6;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_A_CY;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_A_XOR;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_B;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_B1;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_B2;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_B3;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_B4;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_B5;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_B6;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_BO5;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_BO6;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_B_CY;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_B_XOR;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_C;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_C1;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_C2;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_C3;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_C4;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_C5;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_C6;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_CO5;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_CO6;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_C_CY;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_C_XOR;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_D;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_D1;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_D2;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_D3;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_D4;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_D5;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_D6;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_DO5;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_DO6;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_D_CY;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X80Y102_D_XOR;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_A;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_A1;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_A2;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_A3;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_A4;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_A5;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_A6;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_AO5;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_AO6;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_A_CY;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_A_XOR;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_B;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_B1;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_B2;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_B3;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_B4;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_B5;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_B6;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_BO5;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_BO6;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_B_CY;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_B_XOR;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_C;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_C1;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_C2;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_C3;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_C4;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_C5;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_C6;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_CO5;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_CO6;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_C_CY;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_C_XOR;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_D;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_D1;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_D2;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_D3;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_D4;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_D5;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_D6;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_DO5;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_DO6;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_D_CY;
  wire [0:0] CLBLM_R_X53Y102_SLICE_X81Y102_D_XOR;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_A;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_A1;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_A2;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_A3;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_A4;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_A5;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_A6;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_AO5;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_AO6;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_A_CY;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_A_XOR;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_B;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_B1;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_B2;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_B3;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_B4;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_B5;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_B6;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_BO5;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_BO6;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_B_CY;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_B_XOR;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_C;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_C1;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_C2;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_C3;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_C4;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_C5;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_C6;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_CO5;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_CO6;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_C_CY;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_C_XOR;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_D;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_D1;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_D2;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_D3;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_D4;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_D5;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_D6;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_DO5;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_DO6;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_D_CY;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X80Y103_D_XOR;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_A;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_A1;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_A2;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_A3;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_A4;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_A5;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_A6;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_AMUX;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_AO5;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_AO6;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_AX;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_A_CY;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_A_XOR;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_B;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_B1;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_B2;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_B3;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_B4;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_B5;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_B6;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_BMUX;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_BO5;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_BO6;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_B_CY;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_B_XOR;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_C;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_C1;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_C2;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_C3;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_C4;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_C5;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_C6;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_CMUX;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_CO5;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_CO6;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_COUT;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_CX;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_C_CY;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_C_XOR;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_D;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_D1;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_D2;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_D3;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_D4;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_D5;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_D6;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_DMUX;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_DO5;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_DO6;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_DX;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_D_CY;
  wire [0:0] CLBLM_R_X53Y103_SLICE_X81Y103_D_XOR;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_A;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_A1;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_A2;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_A3;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_A4;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_A5;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_A6;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_AMUX;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_AO5;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_AO6;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_A_CY;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_A_XOR;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_B;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_B1;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_B2;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_B3;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_B4;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_B5;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_B6;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_BO5;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_BO6;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_B_CY;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_B_XOR;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_C;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_C1;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_C2;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_C3;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_C4;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_C5;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_C6;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_CMUX;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_CO5;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_CO6;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_C_CY;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_C_XOR;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_D;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_D1;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_D2;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_D3;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_D4;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_D5;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_D6;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_DMUX;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_DO5;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_DO6;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_D_CY;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X80Y104_D_XOR;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_A;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_A1;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_A2;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_A3;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_A4;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_A5;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_A6;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_AMUX;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_AO5;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_AO6;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_AX;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_A_CY;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_A_XOR;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_B;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_B1;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_B2;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_B3;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_B4;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_B5;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_B6;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_BMUX;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_BO5;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_BO6;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_BX;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_B_CY;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_B_XOR;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_C;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_C1;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_C2;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_C3;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_C4;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_C5;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_C6;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_CIN;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_CMUX;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_CO5;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_CO6;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_COUT;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_CX;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_C_CY;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_C_XOR;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_D;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_D1;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_D2;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_D3;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_D4;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_D5;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_D6;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_DMUX;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_DO5;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_DO6;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_DX;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_D_CY;
  wire [0:0] CLBLM_R_X53Y104_SLICE_X81Y104_D_XOR;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_A;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_A1;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_A2;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_A3;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_A4;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_A5;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_A6;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_AO5;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_AO6;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_A_CY;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_A_XOR;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_B;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_B1;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_B2;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_B3;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_B4;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_B5;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_B6;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_BO5;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_BO6;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_B_CY;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_B_XOR;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_C;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_C1;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_C2;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_C3;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_C4;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_C5;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_C6;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_CO5;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_CO6;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_C_CY;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_C_XOR;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_D;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_D1;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_D2;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_D3;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_D4;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_D5;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_D6;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_DO5;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_DO6;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_D_CY;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X80Y105_D_XOR;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_A;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_A1;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_A2;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_A3;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_A4;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_A5;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_A6;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_AMUX;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_AO5;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_AO6;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_AX;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_A_CY;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_A_XOR;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_B;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_B1;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_B2;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_B3;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_B4;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_B5;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_B6;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_BMUX;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_BO5;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_BO6;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_B_CY;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_B_XOR;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_C;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_C1;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_C2;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_C3;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_C4;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_C5;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_C6;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_CIN;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_CMUX;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_CO5;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_CO6;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_COUT;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_CX;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_C_CY;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_C_XOR;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_D;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_D1;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_D2;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_D3;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_D4;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_D5;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_D6;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_DO5;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_DO6;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_DX;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_D_CY;
  wire [0:0] CLBLM_R_X53Y105_SLICE_X81Y105_D_XOR;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_A;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_A1;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_A2;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_A3;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_A4;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_A5;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_A6;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_AMUX;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_AO5;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_AO6;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_A_CY;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_A_XOR;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_B;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_B1;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_B2;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_B3;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_B4;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_B5;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_B6;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_BO5;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_BO6;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_B_CY;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_B_XOR;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_C;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_C1;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_C2;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_C3;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_C4;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_C5;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_C6;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_CO5;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_CO6;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_C_CY;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_C_XOR;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_D;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_D1;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_D2;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_D3;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_D4;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_D5;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_D6;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_DO5;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_DO6;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_D_CY;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X80Y106_D_XOR;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_A;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_A1;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_A2;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_A3;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_A4;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_A5;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_A6;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_AMUX;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_AO5;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_AO6;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_AX;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_A_CY;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_A_XOR;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_B;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_B1;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_B2;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_B3;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_B4;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_B5;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_B6;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_BMUX;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_BO5;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_BO6;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_B_CY;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_B_XOR;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_C;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_C1;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_C2;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_C3;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_C4;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_C5;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_C6;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_CMUX;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_CO5;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_CO6;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_COUT;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_CX;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_C_CY;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_C_XOR;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_D;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_D1;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_D2;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_D3;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_D4;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_D5;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_D6;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_DMUX;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_DO5;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_DO6;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_DX;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_D_CY;
  wire [0:0] CLBLM_R_X53Y106_SLICE_X81Y106_D_XOR;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_A;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_A1;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_A2;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_A3;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_A4;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_A5;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_A6;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_AMUX;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_AO5;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_AO6;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_A_CY;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_A_XOR;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_B;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_B1;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_B2;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_B3;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_B4;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_B5;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_B6;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_BMUX;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_BO5;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_BO6;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_B_CY;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_B_XOR;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_C;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_C1;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_C2;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_C3;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_C4;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_C5;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_C6;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_CO5;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_CO6;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_C_CY;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_C_XOR;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_D;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_D1;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_D2;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_D3;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_D4;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_D5;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_D6;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_DO5;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_DO6;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_D_CY;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X80Y107_D_XOR;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_A;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_A1;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_A2;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_A3;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_A4;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_A5;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_A6;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_AMUX;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_AO5;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_AO6;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_AX;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_A_CY;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_A_XOR;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_B;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_B1;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_B2;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_B3;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_B4;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_B5;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_B6;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_BMUX;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_BO5;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_BO6;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_BX;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_B_CY;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_B_XOR;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_C;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_C1;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_C2;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_C3;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_C4;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_C5;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_C6;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_CIN;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_CMUX;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_CO5;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_CO6;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_COUT;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_CX;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_C_CY;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_C_XOR;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_D;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_D1;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_D2;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_D3;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_D4;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_D5;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_D6;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_DMUX;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_DO5;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_DO6;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_DX;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_D_CY;
  wire [0:0] CLBLM_R_X53Y107_SLICE_X81Y107_D_XOR;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_A;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_A1;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_A2;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_A3;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_A4;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_A5;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_A6;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_AO5;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_AO6;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_A_CY;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_A_XOR;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_B;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_B1;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_B2;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_B3;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_B4;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_B5;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_B6;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_BO5;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_BO6;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_B_CY;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_B_XOR;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_C;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_C1;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_C2;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_C3;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_C4;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_C5;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_C6;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_CMUX;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_CO5;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_CO6;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_C_CY;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_C_XOR;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_D;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_D1;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_D2;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_D3;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_D4;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_D5;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_D6;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_DO5;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_DO6;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_D_CY;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X80Y108_D_XOR;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_A;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_A1;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_A2;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_A3;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_A4;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_A5;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_A6;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_AMUX;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_AO5;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_AO6;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_AX;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_A_CY;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_A_XOR;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_B;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_B1;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_B2;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_B3;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_B4;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_B5;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_B6;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_BMUX;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_BO5;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_BO6;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_B_CY;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_B_XOR;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_C;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_C1;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_C2;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_C3;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_C4;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_C5;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_C6;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_CIN;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_CMUX;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_CO5;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_CO6;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_COUT;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_CX;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_C_CY;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_C_XOR;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_D;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_D1;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_D2;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_D3;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_D4;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_D5;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_D6;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_DO5;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_DO6;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_DX;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_D_CY;
  wire [0:0] CLBLM_R_X53Y108_SLICE_X81Y108_D_XOR;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_A;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_A1;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_A2;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_A3;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_A4;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_A5;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_A6;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_AO5;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_AO6;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_A_CY;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_A_XOR;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_B;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_B1;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_B2;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_B3;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_B4;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_B5;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_B6;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_BO5;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_BO6;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_B_CY;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_B_XOR;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_C;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_C1;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_C2;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_C3;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_C4;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_C5;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_C6;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_CO5;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_CO6;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_C_CY;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_C_XOR;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_D;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_D1;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_D2;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_D3;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_D4;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_D5;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_D6;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_DO5;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_DO6;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_D_CY;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X80Y98_D_XOR;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_A;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_A1;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_A2;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_A3;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_A4;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_A5;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_A6;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_AO5;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_AO6;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_A_CY;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_A_XOR;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_B;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_B1;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_B2;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_B3;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_B4;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_B5;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_B6;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_BO5;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_BO6;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_B_CY;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_B_XOR;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_C;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_C1;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_C2;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_C3;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_C4;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_C5;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_C6;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_CO5;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_CO6;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_C_CY;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_C_XOR;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_D;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_D1;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_D2;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_D3;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_D4;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_D5;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_D6;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_DO5;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_DO6;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_D_CY;
  wire [0:0] CLBLM_R_X53Y98_SLICE_X81Y98_D_XOR;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_A;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_A1;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_A2;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_A3;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_A4;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_A5;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_A6;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_AMUX;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_AO5;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_AO6;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_A_CY;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_A_XOR;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_B;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_B1;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_B2;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_B3;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_B4;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_B5;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_B6;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_BMUX;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_BO5;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_BO6;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_B_CY;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_B_XOR;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_C;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_C1;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_C2;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_C3;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_C4;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_C5;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_C6;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_CO5;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_CO6;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_C_CY;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_C_XOR;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_D;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_D1;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_D2;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_D3;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_D4;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_D5;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_D6;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_DMUX;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_DO5;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_DO6;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_D_CY;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X80Y99_D_XOR;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_A;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_A1;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_A2;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_A3;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_A4;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_A5;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_A6;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_AMUX;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_AO5;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_AO6;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_AQ;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_AX;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_A_CY;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_A_XOR;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_B;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_B1;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_B2;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_B3;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_B4;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_B5;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_B6;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_BO5;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_BO6;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_BQ;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_B_CY;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_B_XOR;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_C;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_C1;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_C2;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_C3;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_C4;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_C5;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_C6;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_CE;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_CLK;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_CO5;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_CO6;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_C_CY;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_C_XOR;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_D;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_D1;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_D2;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_D3;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_D4;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_D5;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_D6;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_DO5;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_DO6;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_D_CY;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_D_XOR;
  wire [0:0] CLBLM_R_X53Y99_SLICE_X81Y99_SR;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_A;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_A1;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_A2;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_A3;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_A4;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_A5;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_A6;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_AMUX;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_AO5;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_AO6;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_AQ;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_AX;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_A_CY;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_A_XOR;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_B;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_B1;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_B2;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_B3;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_B4;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_B5;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_B5Q;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_B6;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_BMUX;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_BO5;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_BO6;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_BQ;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_BX;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_B_CY;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_B_XOR;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_C;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_C1;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_C2;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_C3;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_C4;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_C5;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_C5Q;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_C6;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_CE;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_CLK;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_CMUX;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_CO5;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_CO6;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_CQ;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_CX;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_C_CY;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_C_XOR;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_D;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_D1;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_D2;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_D3;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_D4;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_D5;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_D6;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_DO5;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_DO6;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_DQ;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_DX;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_D_CY;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_D_XOR;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X88Y100_SR;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_A;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_A1;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_A2;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_A3;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_A4;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_A5;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_A6;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_AO5;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_AO6;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_AQ;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_A_CY;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_A_XOR;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_B;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_B1;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_B2;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_B3;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_B4;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_B5;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_B6;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_BO5;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_BO6;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_BQ;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_B_CY;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_B_XOR;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_C;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_C1;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_C2;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_C3;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_C4;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_C5;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_C6;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_CE;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_CLK;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_CO5;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_CO6;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_CQ;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_C_CY;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_C_XOR;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_D;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_D1;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_D2;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_D3;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_D4;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_D5;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_D6;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_DO5;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_DO6;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_DQ;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_D_CY;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_D_XOR;
  wire [0:0] CLBLM_R_X59Y100_SLICE_X89Y100_SR;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_A;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_A1;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_A2;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_A3;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_A4;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_A5;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_A6;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_AO5;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_AO6;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_A_CY;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_A_XOR;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_B;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_B1;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_B2;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_B3;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_B4;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_B5;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_B6;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_BO5;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_BO6;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_B_CY;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_B_XOR;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_C;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_C1;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_C2;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_C3;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_C4;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_C5;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_C6;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_CO5;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_CO6;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_C_CY;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_C_XOR;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_D;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_D1;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_D2;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_D3;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_D4;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_D5;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_D6;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_DMUX;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_DO5;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_DO6;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_D_CY;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X88Y101_D_XOR;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_A;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_A1;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_A2;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_A3;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_A4;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_A5;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_A6;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_AO5;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_AO6;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_AQ;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_A_CY;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_A_XOR;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_B;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_B1;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_B2;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_B3;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_B4;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_B5;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_B6;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_BMUX;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_BO5;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_BO6;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_B_CY;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_B_XOR;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_C;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_C1;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_C2;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_C3;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_C4;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_C5;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_C6;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_CE;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_CLK;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_CO5;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_CO6;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_C_CY;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_C_XOR;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_D;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_D1;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_D2;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_D3;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_D4;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_D5;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_D6;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_DO5;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_DO6;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_D_CY;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_D_XOR;
  wire [0:0] CLBLM_R_X59Y101_SLICE_X89Y101_SR;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_A;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_A1;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_A2;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_A3;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_A4;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_A5;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_A6;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_AO5;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_AO6;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_AQ;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_A_CY;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_A_XOR;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_B;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_B1;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_B2;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_B3;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_B4;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_B5;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_B6;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_BO5;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_BO6;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_B_CY;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_B_XOR;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_C;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_C1;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_C2;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_C3;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_C4;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_C5;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_C6;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_CE;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_CLK;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_CO5;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_CO6;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_C_CY;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_C_XOR;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_D;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_D1;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_D2;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_D3;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_D4;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_D5;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_D6;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_DO5;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_DO6;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_D_CY;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_D_XOR;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X88Y102_SR;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_A;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_A1;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_A2;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_A3;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_A4;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_A5;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_A6;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_AO5;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_AO6;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_AQ;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_A_CY;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_A_XOR;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_B;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_B1;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_B2;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_B3;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_B4;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_B5;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_B6;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_BO5;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_BO6;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_B_CY;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_B_XOR;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_C;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_C1;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_C2;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_C3;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_C4;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_C5;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_C6;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_CE;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_CLK;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_CO5;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_CO6;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_C_CY;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_C_XOR;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_D;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_D1;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_D2;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_D3;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_D4;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_D5;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_D6;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_DMUX;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_DO5;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_DO6;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_D_CY;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_D_XOR;
  wire [0:0] CLBLM_R_X59Y102_SLICE_X89Y102_SR;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_A;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_A1;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_A2;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_A3;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_A4;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_A5;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_A6;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_AMUX;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_AO5;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_AO6;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_AX;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_A_CY;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_A_XOR;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_B;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_B1;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_B2;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_B3;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_B4;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_B5;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_B6;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_BO5;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_BO6;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_BQ;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_BX;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_B_CY;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_B_XOR;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_C;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_C1;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_C2;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_C3;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_C4;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_C5;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_C6;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_CE;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_CLK;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_CO5;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_CO6;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_CQ;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_CX;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_C_CY;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_C_XOR;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_D;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_D1;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_D2;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_D3;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_D4;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_D5;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_D6;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_DO5;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_DO6;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_DQ;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_DX;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_D_CY;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_D_XOR;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_F7AMUX_O;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X88Y103_SR;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_A;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_A1;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_A2;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_A3;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_A4;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_A5;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_A5Q;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_A6;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_AMUX;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_AO5;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_AO6;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_AX;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_A_CY;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_A_XOR;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_B;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_B1;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_B2;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_B3;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_B4;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_B5;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_B6;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_BO5;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_BO6;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_B_CY;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_B_XOR;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_C;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_C1;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_C2;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_C3;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_C4;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_C5;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_C6;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_CE;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_CLK;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_CO5;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_CO6;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_CQ;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_C_CY;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_C_XOR;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_D;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_D1;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_D2;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_D3;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_D4;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_D5;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_D6;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_DO5;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_DO6;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_DQ;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_D_CY;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_D_XOR;
  wire [0:0] CLBLM_R_X59Y103_SLICE_X89Y103_SR;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_A;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_A1;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_A2;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_A3;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_A4;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_A5;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_A6;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_AMUX;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_AO5;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_AO6;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_AQ;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_AX;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_A_CY;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_A_XOR;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_B;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_B1;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_B2;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_B3;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_B4;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_B5;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_B6;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_BMUX;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_BO5;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_BO6;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_BQ;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_BX;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_B_CY;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_B_XOR;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_C;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_C1;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_C2;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_C3;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_C4;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_C5;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_C6;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_CE;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_CLK;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_CMUX;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_CO5;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_CO6;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_C_CY;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_C_XOR;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_D;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_D1;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_D2;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_D3;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_D4;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_D5;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_D6;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_DO5;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_DO6;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_D_CY;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_D_XOR;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X88Y104_SR;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_A;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_A1;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_A2;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_A3;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_A4;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_A5;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_A6;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_AMUX;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_AO5;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_AO6;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_AX;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_A_CY;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_A_XOR;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_B;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_B1;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_B2;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_B3;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_B4;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_B5;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_B6;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_BO5;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_BO6;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_B_CY;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_B_XOR;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_C;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_C1;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_C2;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_C3;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_C4;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_C5;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_C6;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_CE;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_CLK;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_CO5;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_CO6;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_CQ;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_C_CY;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_C_XOR;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_D;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_D1;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_D2;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_D3;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_D4;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_D5;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_D6;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_DO5;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_DO6;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_D_CY;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_D_XOR;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_F7AMUX_O;
  wire [0:0] CLBLM_R_X59Y104_SLICE_X89Y104_SR;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_A;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_A1;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_A2;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_A3;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_A4;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_A5;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_A6;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_AMUX;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_AO5;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_AO6;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_AX;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_A_CY;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_A_XOR;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_B;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_B1;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_B2;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_B3;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_B4;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_B5;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_B6;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_BO5;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_BO6;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_BQ;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_BX;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_B_CY;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_B_XOR;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_C;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_C1;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_C2;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_C3;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_C4;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_C5;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_C6;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_CE;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_CLK;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_CO5;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_CO6;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_C_CY;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_C_XOR;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_D;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_D1;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_D2;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_D3;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_D4;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_D5;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_D6;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_DO5;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_DO6;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_D_CY;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_D_XOR;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_F7AMUX_O;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X88Y105_SR;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_A;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_A1;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_A2;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_A3;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_A4;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_A5;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_A6;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_AMUX;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_AO5;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_AO6;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_AX;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_A_CY;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_A_XOR;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_B;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_B1;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_B2;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_B3;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_B4;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_B5;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_B6;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_BO5;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_BO6;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_B_CY;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_B_XOR;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_C;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_C1;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_C2;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_C3;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_C4;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_C5;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_C6;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_CE;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_CLK;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_CO5;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_CO6;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_CQ;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_C_CY;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_C_XOR;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_D;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_D1;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_D2;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_D3;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_D4;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_D5;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_D6;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_DO5;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_DO6;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_D_CY;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_D_XOR;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_F7AMUX_O;
  wire [0:0] CLBLM_R_X59Y105_SLICE_X89Y105_SR;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_A;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_A1;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_A2;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_A3;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_A4;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_A5;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_A6;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_AO5;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_AO6;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_AQ;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_A_CY;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_A_XOR;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_B;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_B1;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_B2;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_B3;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_B4;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_B5;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_B6;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_BO5;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_BO6;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_BQ;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_B_CY;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_B_XOR;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_C;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_C1;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_C2;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_C3;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_C4;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_C5;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_C6;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_CE;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_CLK;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_CO5;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_CO6;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_C_CY;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_C_XOR;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_D;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_D1;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_D2;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_D3;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_D4;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_D5;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_D6;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_DO5;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_DO6;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_D_CY;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_D_XOR;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X88Y106_SR;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_A;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_A1;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_A2;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_A3;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_A4;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_A5;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_A6;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_AMUX;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_AO5;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_AO6;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_A_CY;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_A_XOR;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_B;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_B1;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_B2;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_B3;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_B4;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_B5;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_B6;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_BO5;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_BO6;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_BQ;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_B_CY;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_B_XOR;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_C;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_C1;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_C2;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_C3;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_C4;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_C5;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_C6;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_CE;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_CLK;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_CO5;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_CO6;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_CQ;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_C_CY;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_C_XOR;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_D;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_D1;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_D2;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_D3;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_D4;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_D5;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_D6;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_DO5;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_DO6;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_D_CY;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_D_XOR;
  wire [0:0] CLBLM_R_X59Y106_SLICE_X89Y106_SR;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_A;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_A1;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_A2;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_A3;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_A4;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_A5;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_A6;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_AO5;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_AO6;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_AQ;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_AX;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_A_CY;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_A_XOR;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_B;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_B1;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_B2;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_B3;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_B4;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_B5;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_B6;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_BO5;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_BO6;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_B_CY;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_B_XOR;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_C;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_C1;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_C2;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_C3;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_C4;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_C5;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_C6;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_CE;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_CLK;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_CO5;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_CO6;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_C_CY;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_C_XOR;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_D;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_D1;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_D2;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_D3;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_D4;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_D5;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_D6;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_DO5;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_DO6;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_D_CY;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_D_XOR;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X88Y107_SR;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_A;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_A1;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_A2;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_A3;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_A4;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_A5;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_A6;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_AMUX;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_AO5;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_AO6;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_AX;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_A_CY;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_A_XOR;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_B;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_B1;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_B2;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_B3;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_B4;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_B5;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_B6;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_BMUX;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_BO5;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_BO6;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_BQ;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_BX;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_B_CY;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_B_XOR;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_C;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_C1;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_C2;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_C3;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_C4;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_C5;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_C6;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_CE;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_CLK;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_CMUX;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_CO5;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_CO6;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_COUT;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_CX;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_C_CY;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_C_XOR;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_D;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_D1;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_D2;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_D3;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_D4;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_D5;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_D6;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_DMUX;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_DO5;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_DO6;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_DX;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_D_CY;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_D_XOR;
  wire [0:0] CLBLM_R_X59Y107_SLICE_X89Y107_SR;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_A;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_A1;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_A2;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_A3;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_A4;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_A5;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_A6;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_AMUX;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_AO5;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_AO6;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_AQ;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_AX;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_A_CY;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_A_XOR;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_B;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_B1;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_B2;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_B3;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_B4;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_B5;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_B6;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_BMUX;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_BO5;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_BO6;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_BX;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_B_CY;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_B_XOR;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_C;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_C1;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_C2;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_C3;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_C4;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_C5;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_C6;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_CE;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_CLK;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_CMUX;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_CO5;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_CO6;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_COUT;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_CX;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_C_CY;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_C_XOR;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_D;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_D1;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_D2;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_D3;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_D4;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_D5;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_D6;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_DMUX;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_DO5;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_DO6;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_DX;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_D_CY;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_D_XOR;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X88Y108_SR;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_A;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_A1;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_A2;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_A3;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_A4;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_A5;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_A6;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_AMUX;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_AO5;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_AO6;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_AQ;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_AX;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_A_CY;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_A_XOR;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_B;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_B1;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_B2;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_B3;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_B4;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_B5;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_B6;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_BMUX;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_BO5;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_BO6;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_BX;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_B_CY;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_B_XOR;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_C;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_C1;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_C2;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_C3;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_C4;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_C5;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_C6;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_CE;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_CIN;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_CLK;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_CMUX;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_CO5;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_CO6;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_COUT;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_CX;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_C_CY;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_C_XOR;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_D;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_D1;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_D2;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_D3;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_D4;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_D5;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_D6;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_DMUX;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_DO5;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_DO6;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_DX;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_D_CY;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_D_XOR;
  wire [0:0] CLBLM_R_X59Y108_SLICE_X89Y108_SR;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_A;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_A1;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_A2;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_A3;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_A4;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_A5;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_A6;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_AMUX;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_AO5;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_AO6;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_AX;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_A_CY;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_A_XOR;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_B;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_B1;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_B2;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_B3;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_B4;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_B5;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_B6;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_BMUX;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_BO5;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_BO6;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_BX;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_B_CY;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_B_XOR;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_C;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_C1;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_C2;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_C3;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_C4;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_C5;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_C6;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_CIN;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_CMUX;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_CO5;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_CO6;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_COUT;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_CX;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_C_CY;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_C_XOR;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_D;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_D1;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_D2;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_D3;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_D4;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_D5;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_D6;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_DMUX;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_DO5;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_DO6;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_DX;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_D_CY;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X88Y109_D_XOR;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_A;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_A1;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_A2;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_A3;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_A4;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_A5;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_A6;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_AMUX;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_AO5;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_AO6;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_AX;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_A_CY;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_A_XOR;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_B;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_B1;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_B2;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_B3;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_B4;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_B5;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_B6;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_BMUX;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_BO5;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_BO6;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_BX;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_B_CY;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_B_XOR;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_C;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_C1;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_C2;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_C3;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_C4;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_C5;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_C6;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_CIN;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_CMUX;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_CO5;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_CO6;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_COUT;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_CX;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_C_CY;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_C_XOR;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_D;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_D1;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_D2;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_D3;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_D4;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_D5;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_D6;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_DO5;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_DO6;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_DX;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_D_CY;
  wire [0:0] CLBLM_R_X59Y109_SLICE_X89Y109_D_XOR;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_A;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_A1;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_A2;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_A3;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_A4;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_A5;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_A6;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_AMUX;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_AO5;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_AO6;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_AX;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_A_CY;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_A_XOR;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_B;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_B1;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_B2;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_B3;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_B4;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_B5;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_B6;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_BMUX;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_BO5;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_BO6;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_BX;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_B_CY;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_B_XOR;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_C;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_C1;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_C2;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_C3;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_C4;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_C5;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_C6;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_CIN;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_CMUX;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_CO5;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_CO6;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_COUT;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_CX;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_C_CY;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_C_XOR;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_D;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_D1;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_D2;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_D3;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_D4;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_D5;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_D6;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_DMUX;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_DO5;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_DO6;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_DX;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_D_CY;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X88Y110_D_XOR;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_A;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_A1;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_A2;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_A3;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_A4;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_A5;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_A6;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_AO5;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_AO6;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_AQ;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_A_CY;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_A_XOR;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_B;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_B1;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_B2;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_B3;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_B4;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_B5;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_B6;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_BO5;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_BO6;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_B_CY;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_B_XOR;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_C;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_C1;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_C2;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_C3;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_C4;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_C5;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_C6;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_CE;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_CLK;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_CO5;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_CO6;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_C_CY;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_C_XOR;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_D;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_D1;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_D2;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_D3;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_D4;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_D5;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_D6;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_DMUX;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_DO5;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_DO6;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_D_CY;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_D_XOR;
  wire [0:0] CLBLM_R_X59Y110_SLICE_X89Y110_SR;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_A;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_A1;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_A2;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_A3;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_A4;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_A5;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_A6;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_AMUX;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_AO5;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_AO6;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_A_CY;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_A_XOR;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_B;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_B1;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_B2;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_B3;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_B4;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_B5;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_B6;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_BO5;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_BO6;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_B_CY;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_B_XOR;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_C;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_C1;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_C2;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_C3;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_C4;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_C5;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_C6;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_CO5;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_CO6;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_C_CY;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_C_XOR;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_D;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_D1;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_D2;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_D3;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_D4;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_D5;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_D6;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_DO5;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_DO6;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_D_CY;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X88Y111_D_XOR;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_A;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_A1;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_A2;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_A3;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_A4;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_A5;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_A6;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_AO5;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_AO6;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_AQ;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_A_CY;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_A_XOR;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_B;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_B1;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_B2;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_B3;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_B4;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_B5;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_B6;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_BO5;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_BO6;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_BQ;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_B_CY;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_B_XOR;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_C;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_C1;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_C2;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_C3;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_C4;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_C5;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_C6;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_CE;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_CLK;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_CO5;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_CO6;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_CQ;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_C_CY;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_C_XOR;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_D;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_D1;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_D2;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_D3;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_D4;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_D5;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_D6;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_DO5;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_DO6;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_D_CY;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_D_XOR;
  wire [0:0] CLBLM_R_X59Y111_SLICE_X89Y111_SR;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_A;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_A1;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_A2;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_A3;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_A4;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_A5;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_A6;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_AO5;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_AO6;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_A_CY;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_A_XOR;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_B;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_B1;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_B2;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_B3;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_B4;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_B5;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_B6;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_BO5;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_BO6;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_B_CY;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_B_XOR;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_C;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_C1;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_C2;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_C3;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_C4;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_C5;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_C6;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_CO5;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_CO6;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_C_CY;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_C_XOR;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_D;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_D1;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_D2;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_D3;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_D4;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_D5;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_D6;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_DO5;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_DO6;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_D_CY;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X88Y112_D_XOR;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_A;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_A1;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_A2;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_A3;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_A4;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_A5;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_A6;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_AO5;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_AO6;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_AQ;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_A_CY;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_A_XOR;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_B;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_B1;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_B2;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_B3;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_B4;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_B5;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_B6;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_BO5;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_BO6;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_BQ;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_B_CY;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_B_XOR;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_C;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_C1;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_C2;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_C3;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_C4;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_C5;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_C6;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_CE;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_CLK;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_CO5;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_CO6;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_C_CY;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_C_XOR;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_D;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_D1;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_D2;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_D3;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_D4;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_D5;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_D6;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_DO5;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_DO6;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_D_CY;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_D_XOR;
  wire [0:0] CLBLM_R_X59Y112_SLICE_X89Y112_SR;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_A;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_A1;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_A2;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_A3;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_A4;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_A5;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_A6;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_AO5;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_AO6;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_AQ;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_A_CY;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_A_XOR;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_B;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_B1;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_B2;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_B3;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_B4;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_B5;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_B6;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_BO5;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_BO6;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_BQ;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_B_CY;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_B_XOR;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_C;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_C1;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_C2;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_C3;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_C4;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_C5;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_C6;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_CLK;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_CO5;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_CO6;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_C_CY;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_C_XOR;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_D;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_D1;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_D2;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_D3;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_D4;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_D5;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_D6;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_DMUX;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_DO5;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_DO6;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_D_CY;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_D_XOR;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X88Y96_SR;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_A;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_A1;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_A2;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_A3;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_A4;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_A5;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_A5Q;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_A6;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_AMUX;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_AO5;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_AO6;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_AQ;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_A_CY;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_A_XOR;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_B;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_B1;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_B2;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_B3;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_B4;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_B5;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_B6;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_BO5;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_BO6;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_B_CY;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_B_XOR;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_C;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_C1;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_C2;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_C3;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_C4;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_C5;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_C6;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_CE;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_CLK;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_CO5;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_CO6;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_C_CY;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_C_XOR;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_D;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_D1;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_D2;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_D3;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_D4;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_D5;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_D6;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_DO5;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_DO6;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_D_CY;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_D_XOR;
  wire [0:0] CLBLM_R_X59Y96_SLICE_X89Y96_SR;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_A;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_A1;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_A2;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_A3;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_A4;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_A5;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_A6;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_AO5;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_AO6;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_AQ;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_A_CY;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_A_XOR;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_B;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_B1;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_B2;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_B3;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_B4;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_B5;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_B6;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_BO5;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_BO6;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_BQ;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_B_CY;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_B_XOR;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_C;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_C1;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_C2;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_C3;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_C4;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_C5;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_C6;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_CLK;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_CO5;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_CO6;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_C_CY;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_C_XOR;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_D;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_D1;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_D2;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_D3;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_D4;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_D5;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_D6;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_DO5;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_DO6;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_D_CY;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_D_XOR;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X88Y97_SR;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_A;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_A1;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_A2;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_A3;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_A4;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_A5;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_A5Q;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_A6;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_AMUX;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_AO5;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_AO6;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_AQ;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_AX;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_A_CY;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_A_XOR;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_B;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_B1;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_B2;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_B3;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_B4;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_B5;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_B5Q;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_B6;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_BMUX;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_BO5;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_BO6;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_BQ;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_BX;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_B_CY;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_B_XOR;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_C;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_C1;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_C2;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_C3;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_C4;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_C5;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_C5Q;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_C6;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_CE;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_CLK;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_CMUX;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_CO5;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_CO6;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_CQ;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_CX;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_C_CY;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_C_XOR;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_D;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_D1;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_D2;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_D3;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_D4;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_D5;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_D5Q;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_D6;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_DMUX;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_DO5;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_DO6;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_DQ;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_DX;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_D_CY;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_D_XOR;
  wire [0:0] CLBLM_R_X59Y97_SLICE_X89Y97_SR;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_A;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_A1;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_A2;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_A3;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_A4;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_A5;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_A6;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_AO5;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_AO6;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_AQ;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_A_CY;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_A_XOR;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_B;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_B1;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_B2;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_B3;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_B4;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_B5;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_B6;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_BO5;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_BO6;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_BQ;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_B_CY;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_B_XOR;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_C;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_C1;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_C2;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_C3;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_C4;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_C5;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_C6;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_CE;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_CLK;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_CO5;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_CO6;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_CQ;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_C_CY;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_C_XOR;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_D;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_D1;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_D2;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_D3;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_D4;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_D5;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_D6;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_DO5;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_DO6;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_DQ;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_D_CY;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_D_XOR;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X88Y98_SR;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_A;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_A1;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_A2;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_A3;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_A4;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_A5;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_A5Q;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_A6;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_AMUX;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_AO5;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_AO6;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_AQ;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_A_CY;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_A_XOR;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_B;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_B1;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_B2;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_B3;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_B4;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_B5;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_B5Q;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_B6;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_BMUX;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_BO5;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_BO6;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_BQ;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_B_CY;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_B_XOR;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_C;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_C1;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_C2;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_C3;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_C4;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_C5;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_C5Q;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_C6;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_CE;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_CLK;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_CMUX;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_CO5;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_CO6;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_CQ;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_C_CY;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_C_XOR;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_D;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_D1;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_D2;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_D3;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_D4;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_D5;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_D6;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_DMUX;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_DO5;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_DO6;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_D_CY;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_D_XOR;
  wire [0:0] CLBLM_R_X59Y98_SLICE_X89Y98_SR;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_A;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_A1;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_A2;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_A3;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_A4;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_A5;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_A6;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_AO5;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_AO6;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_AQ;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_A_CY;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_A_XOR;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_B;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_B1;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_B2;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_B3;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_B4;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_B5;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_B5Q;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_B6;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_BMUX;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_BO5;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_BO6;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_BQ;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_B_CY;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_B_XOR;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_C;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_C1;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_C2;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_C3;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_C4;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_C5;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_C6;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_CE;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_CLK;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_CO5;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_CO6;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_CQ;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_C_CY;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_C_XOR;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_D;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_D1;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_D2;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_D3;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_D4;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_D5;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_D6;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_DO5;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_DO6;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_DQ;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_D_CY;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_D_XOR;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X88Y99_SR;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_A;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_A1;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_A2;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_A3;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_A4;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_A5;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_A5Q;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_A6;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_AMUX;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_AO5;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_AO6;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_AQ;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_A_CY;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_A_XOR;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_B;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_B1;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_B2;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_B3;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_B4;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_B5;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_B6;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_BO5;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_BO6;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_BQ;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_B_CY;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_B_XOR;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_C;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_C1;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_C2;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_C3;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_C4;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_C5;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_C6;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_CE;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_CLK;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_CO5;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_CO6;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_C_CY;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_C_XOR;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_D;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_D1;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_D2;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_D3;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_D4;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_D5;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_D6;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_DO5;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_DO6;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_D_CY;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_D_XOR;
  wire [0:0] CLBLM_R_X59Y99_SLICE_X89Y99_SR;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_A;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_A1;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_A2;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_A3;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_A4;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_A5;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_A6;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_AO5;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_AO6;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_AQ;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_A_CY;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_A_XOR;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_B;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_B1;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_B2;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_B3;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_B4;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_B5;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_B6;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_BO5;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_BO6;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_B_CY;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_B_XOR;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_C;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_C1;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_C2;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_C3;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_C4;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_C5;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_C6;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_CLK;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_CO5;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_CO6;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_C_CY;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_C_XOR;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_D;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_D1;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_D2;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_D3;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_D4;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_D5;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_D6;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_DO5;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_DO6;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_D_CY;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_D_XOR;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X94Y100_SR;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_A;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_A1;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_A2;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_A3;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_A4;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_A5;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_A5Q;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_A6;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_AMUX;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_AO5;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_AO6;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_AQ;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_A_CY;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_A_XOR;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_B;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_B1;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_B2;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_B3;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_B4;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_B5;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_B6;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_BO5;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_BO6;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_B_CY;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_B_XOR;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_C;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_C1;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_C2;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_C3;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_C4;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_C5;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_C6;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_CE;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_CLK;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_CO5;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_CO6;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_C_CY;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_C_XOR;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_D;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_D1;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_D2;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_D3;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_D4;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_D5;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_D6;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_DO5;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_DO6;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_D_CY;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_D_XOR;
  wire [0:0] CLBLM_R_X63Y100_SLICE_X95Y100_SR;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_A;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_A1;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_A2;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_A3;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_A4;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_A5;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_A6;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_AO5;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_AO6;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_A_CY;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_A_XOR;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_B;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_B1;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_B2;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_B3;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_B4;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_B5;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_B6;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_BO5;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_BO6;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_B_CY;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_B_XOR;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_C;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_C1;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_C2;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_C3;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_C4;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_C5;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_C6;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_CO5;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_CO6;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_C_CY;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_C_XOR;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_D;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_D1;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_D2;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_D3;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_D4;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_D5;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_D6;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_DO5;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_DO6;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_D_CY;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X94Y101_D_XOR;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_A;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_A1;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_A2;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_A3;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_A4;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_A5;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_A6;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_AO5;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_AO6;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_AQ;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_A_CY;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_A_XOR;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_B;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_B1;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_B2;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_B3;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_B4;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_B5;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_B6;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_BO5;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_BO6;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_B_CY;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_B_XOR;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_C;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_C1;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_C2;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_C3;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_C4;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_C5;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_C6;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_CE;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_CLK;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_CO5;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_CO6;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_C_CY;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_C_XOR;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_D;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_D1;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_D2;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_D3;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_D4;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_D5;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_D6;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_DO5;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_DO6;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_D_CY;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_D_XOR;
  wire [0:0] CLBLM_R_X63Y101_SLICE_X95Y101_SR;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_A;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_A1;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_A2;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_A3;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_A4;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_A5;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_A6;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_AO5;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_AO6;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_A_CY;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_A_XOR;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_B;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_B1;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_B2;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_B3;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_B4;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_B5;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_B6;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_BO5;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_BO6;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_B_CY;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_B_XOR;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_C;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_C1;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_C2;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_C3;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_C4;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_C5;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_C6;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_CO5;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_CO6;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_C_CY;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_C_XOR;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_D;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_D1;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_D2;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_D3;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_D4;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_D5;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_D6;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_DO5;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_DO6;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_D_CY;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X94Y102_D_XOR;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_A;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_A1;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_A2;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_A3;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_A4;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_A5;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_A6;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_AO5;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_AO6;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_A_CY;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_A_XOR;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_B;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_B1;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_B2;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_B3;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_B4;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_B5;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_B6;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_BO5;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_BO6;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_B_CY;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_B_XOR;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_C;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_C1;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_C2;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_C3;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_C4;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_C5;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_C6;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_CO5;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_CO6;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_C_CY;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_C_XOR;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_D;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_D1;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_D2;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_D3;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_D4;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_D5;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_D6;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_DO5;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_DO6;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_D_CY;
  wire [0:0] CLBLM_R_X63Y102_SLICE_X95Y102_D_XOR;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_A;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_A1;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_A2;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_A3;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_A4;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_A5;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_A6;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_AO5;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_AO6;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_A_CY;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_A_XOR;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_B;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_B1;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_B2;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_B3;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_B4;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_B5;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_B6;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_BO5;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_BO6;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_B_CY;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_B_XOR;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_C;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_C1;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_C2;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_C3;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_C4;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_C5;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_C6;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_CO5;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_CO6;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_C_CY;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_C_XOR;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_D;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_D1;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_D2;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_D3;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_D4;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_D5;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_D6;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_DO5;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_DO6;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_D_CY;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X94Y103_D_XOR;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_A;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_A1;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_A2;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_A3;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_A4;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_A5;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_A6;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_AO5;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_AO6;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_AQ;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_A_CY;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_A_XOR;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_B;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_B1;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_B2;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_B3;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_B4;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_B5;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_B6;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_BO5;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_BO6;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_BQ;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_B_CY;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_B_XOR;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_C;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_C1;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_C2;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_C3;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_C4;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_C5;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_C6;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_CE;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_CLK;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_CO5;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_CO6;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_CQ;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_C_CY;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_C_XOR;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_D;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_D1;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_D2;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_D3;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_D4;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_D5;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_D6;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_DO5;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_DO6;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_D_CY;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_D_XOR;
  wire [0:0] CLBLM_R_X63Y103_SLICE_X95Y103_SR;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_A;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_A1;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_A2;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_A3;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_A4;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_A5;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_A6;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_AO5;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_AO6;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_AQ;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_A_CY;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_A_XOR;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_B;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_B1;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_B2;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_B3;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_B4;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_B5;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_B6;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_BO5;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_BO6;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_BQ;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_B_CY;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_B_XOR;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_C;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_C1;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_C2;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_C3;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_C4;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_C5;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_C6;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_CE;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_CLK;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_CMUX;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_CO5;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_CO6;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_C_CY;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_C_XOR;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_D;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_D1;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_D2;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_D3;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_D4;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_D5;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_D6;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_DO5;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_DO6;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_D_CY;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_D_XOR;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X94Y104_SR;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_A;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_A1;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_A2;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_A3;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_A4;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_A5;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_A6;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_AO5;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_AO6;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_A_CY;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_A_XOR;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_B;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_B1;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_B2;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_B3;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_B4;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_B5;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_B6;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_BO5;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_BO6;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_B_CY;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_B_XOR;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_C;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_C1;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_C2;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_C3;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_C4;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_C5;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_C6;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_CO5;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_CO6;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_C_CY;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_C_XOR;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_D;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_D1;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_D2;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_D3;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_D4;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_D5;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_D6;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_DO5;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_DO6;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_D_CY;
  wire [0:0] CLBLM_R_X63Y104_SLICE_X95Y104_D_XOR;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_A;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_A1;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_A2;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_A3;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_A4;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_A5;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_A6;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_AMUX;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_AO5;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_AO6;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_AQ;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_AX;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_A_CY;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_A_XOR;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_B;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_B1;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_B2;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_B3;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_B4;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_B5;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_B6;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_BMUX;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_BO5;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_BO6;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_BX;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_B_CY;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_B_XOR;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_C;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_C1;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_C2;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_C3;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_C4;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_C5;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_C6;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_CE;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_CLK;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_CMUX;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_CO5;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_CO6;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_COUT;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_CX;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_C_CY;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_C_XOR;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_D;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_D1;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_D2;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_D3;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_D4;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_D5;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_D6;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_DMUX;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_DO5;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_DO6;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_DX;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_D_CY;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_D_XOR;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X94Y105_SR;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_A;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_A1;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_A2;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_A3;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_A4;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_A5;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_A6;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_AMUX;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_AO5;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_AO6;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_AX;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_A_CY;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_A_XOR;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_B;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_B1;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_B2;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_B3;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_B4;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_B5;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_B6;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_BMUX;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_BO5;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_BO6;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_BX;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_B_CY;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_B_XOR;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_C;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_C1;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_C2;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_C3;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_C4;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_C5;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_C6;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_CMUX;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_CO5;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_CO6;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_COUT;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_CX;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_C_CY;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_C_XOR;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_D;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_D1;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_D2;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_D3;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_D4;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_D5;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_D6;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_DMUX;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_DO5;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_DO6;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_DX;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_D_CY;
  wire [0:0] CLBLM_R_X63Y105_SLICE_X95Y105_D_XOR;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_A;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_A1;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_A2;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_A3;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_A4;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_A5;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_A6;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_AMUX;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_AO5;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_AO6;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_AX;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_A_CY;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_A_XOR;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_B;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_B1;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_B2;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_B3;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_B4;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_B5;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_B6;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_BMUX;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_BO5;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_BO6;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_BX;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_B_CY;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_B_XOR;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_C;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_C1;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_C2;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_C3;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_C4;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_C5;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_C6;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_CIN;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_CMUX;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_CO5;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_CO6;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_COUT;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_CX;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_C_CY;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_C_XOR;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_D;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_D1;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_D2;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_D3;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_D4;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_D5;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_D6;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_DMUX;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_DO5;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_DO6;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_DX;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_D_CY;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X94Y106_D_XOR;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_A;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_A1;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_A2;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_A3;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_A4;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_A5;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_A6;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_AMUX;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_AO5;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_AO6;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_AX;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_A_CY;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_A_XOR;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_B;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_B1;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_B2;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_B3;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_B4;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_B5;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_B6;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_BMUX;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_BO5;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_BO6;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_BX;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_B_CY;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_B_XOR;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_C;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_C1;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_C2;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_C3;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_C4;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_C5;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_C6;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_CIN;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_CMUX;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_CO5;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_CO6;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_COUT;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_CX;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_C_CY;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_C_XOR;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_D;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_D1;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_D2;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_D3;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_D4;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_D5;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_D6;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_DMUX;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_DO5;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_DO6;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_DX;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_D_CY;
  wire [0:0] CLBLM_R_X63Y106_SLICE_X95Y106_D_XOR;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_A;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_A1;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_A2;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_A3;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_A4;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_A5;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_A6;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_AMUX;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_AO5;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_AO6;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_AX;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_A_CY;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_A_XOR;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_B;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_B1;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_B2;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_B3;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_B4;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_B5;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_B6;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_BMUX;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_BO5;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_BO6;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_BX;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_B_CY;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_B_XOR;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_C;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_C1;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_C2;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_C3;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_C4;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_C5;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_C6;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_CIN;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_CMUX;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_CO5;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_CO6;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_COUT;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_CX;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_C_CY;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_C_XOR;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_D;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_D1;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_D2;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_D3;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_D4;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_D5;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_D6;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_DMUX;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_DO5;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_DO6;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_DX;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_D_CY;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X94Y107_D_XOR;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_A;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_A1;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_A2;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_A3;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_A4;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_A5;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_A6;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_AMUX;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_AO5;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_AO6;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_AX;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_A_CY;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_A_XOR;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_B;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_B1;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_B2;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_B3;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_B4;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_B5;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_B6;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_BMUX;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_BO5;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_BO6;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_BX;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_B_CY;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_B_XOR;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_C;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_C1;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_C2;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_C3;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_C4;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_C5;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_C6;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_CIN;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_CMUX;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_CO5;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_CO6;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_COUT;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_CX;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_C_CY;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_C_XOR;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_D;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_D1;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_D2;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_D3;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_D4;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_D5;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_D6;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_DMUX;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_DO5;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_DO6;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_DX;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_D_CY;
  wire [0:0] CLBLM_R_X63Y107_SLICE_X95Y107_D_XOR;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_A;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_A1;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_A2;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_A3;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_A4;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_A5;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_A6;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_AMUX;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_AO5;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_AO6;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_AX;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_A_CY;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_A_XOR;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_B;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_B1;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_B2;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_B3;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_B4;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_B5;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_B6;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_BMUX;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_BO5;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_BO6;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_BX;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_B_CY;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_B_XOR;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_C;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_C1;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_C2;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_C3;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_C4;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_C5;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_C6;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_CIN;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_CMUX;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_CO5;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_CO6;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_COUT;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_CX;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_C_CY;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_C_XOR;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_D;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_D1;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_D2;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_D3;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_D4;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_D5;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_D6;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_DMUX;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_DO5;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_DO6;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_DX;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_D_CY;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X94Y108_D_XOR;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_A;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_A1;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_A2;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_A3;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_A4;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_A5;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_A6;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_AMUX;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_AO5;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_AO6;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_AX;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_A_CY;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_A_XOR;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_B;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_B1;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_B2;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_B3;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_B4;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_B5;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_B6;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_BMUX;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_BO5;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_BO6;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_BX;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_B_CY;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_B_XOR;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_C;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_C1;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_C2;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_C3;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_C4;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_C5;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_C6;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_CIN;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_CMUX;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_CO5;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_CO6;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_COUT;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_CX;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_C_CY;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_C_XOR;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_D;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_D1;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_D2;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_D3;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_D4;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_D5;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_D6;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_DMUX;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_DO5;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_DO6;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_DX;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_D_CY;
  wire [0:0] CLBLM_R_X63Y108_SLICE_X95Y108_D_XOR;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_A;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_A1;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_A2;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_A3;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_A4;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_A5;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_A6;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_AMUX;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_AO5;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_AO6;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_AX;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_A_CY;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_A_XOR;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_B;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_B1;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_B2;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_B3;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_B4;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_B5;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_B6;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_BMUX;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_BO5;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_BO6;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_BX;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_B_CY;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_B_XOR;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_C;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_C1;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_C2;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_C3;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_C4;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_C5;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_C6;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_CIN;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_CMUX;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_CO5;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_CO6;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_COUT;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_CX;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_C_CY;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_C_XOR;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_D;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_D1;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_D2;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_D3;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_D4;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_D5;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_D6;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_DMUX;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_DO5;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_DO6;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_DX;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_D_CY;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X94Y109_D_XOR;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_A;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_A1;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_A2;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_A3;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_A4;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_A5;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_A6;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_AMUX;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_AO5;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_AO6;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_AX;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_A_CY;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_A_XOR;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_B;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_B1;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_B2;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_B3;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_B4;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_B5;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_B6;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_BMUX;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_BO5;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_BO6;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_BX;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_B_CY;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_B_XOR;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_C;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_C1;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_C2;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_C3;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_C4;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_C5;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_C6;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_CIN;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_CMUX;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_CO5;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_CO6;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_COUT;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_CX;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_C_CY;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_C_XOR;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_D;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_D1;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_D2;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_D3;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_D4;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_D5;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_D6;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_DO5;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_DO6;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_DX;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_D_CY;
  wire [0:0] CLBLM_R_X63Y109_SLICE_X95Y109_D_XOR;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_A;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_A1;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_A2;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_A3;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_A4;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_A5;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_A6;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_AO5;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_AO6;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_AQ;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_A_CY;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_A_XOR;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_B;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_B1;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_B2;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_B3;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_B4;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_B5;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_B6;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_BO5;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_BO6;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_B_CY;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_B_XOR;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_C;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_C1;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_C2;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_C3;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_C4;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_C5;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_C6;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_CE;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_CLK;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_CO5;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_CO6;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_C_CY;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_C_XOR;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_D;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_D1;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_D2;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_D3;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_D4;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_D5;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_D6;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_DO5;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_DO6;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_D_CY;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_D_XOR;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X94Y110_SR;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_A;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_A1;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_A2;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_A3;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_A4;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_A5;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_A6;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_AO5;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_AO6;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_A_CY;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_A_XOR;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_B;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_B1;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_B2;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_B3;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_B4;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_B5;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_B6;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_BO5;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_BO6;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_B_CY;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_B_XOR;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_C;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_C1;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_C2;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_C3;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_C4;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_C5;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_C6;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_CO5;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_CO6;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_C_CY;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_C_XOR;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_D;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_D1;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_D2;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_D3;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_D4;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_D5;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_D6;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_DO5;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_DO6;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_D_CY;
  wire [0:0] CLBLM_R_X63Y110_SLICE_X95Y110_D_XOR;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_A;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_A1;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_A2;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_A3;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_A4;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_A5;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_A6;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_AO5;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_AO6;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_AQ;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_A_CY;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_A_XOR;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_B;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_B1;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_B2;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_B3;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_B4;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_B5;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_B6;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_BO5;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_BO6;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_B_CY;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_B_XOR;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_C;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_C1;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_C2;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_C3;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_C4;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_C5;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_C6;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_CE;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_CLK;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_CO5;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_CO6;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_C_CY;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_C_XOR;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_D;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_D1;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_D2;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_D3;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_D4;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_D5;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_D6;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_DO5;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_DO6;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_D_CY;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_D_XOR;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X94Y94_SR;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_A;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_A1;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_A2;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_A3;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_A4;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_A5;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_A6;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_AO5;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_AO6;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_AQ;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_A_CY;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_A_XOR;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_B;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_B1;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_B2;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_B3;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_B4;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_B5;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_B6;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_BO5;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_BO6;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_B_CY;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_B_XOR;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_C;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_C1;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_C2;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_C3;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_C4;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_C5;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_C6;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_CE;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_CLK;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_CO5;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_CO6;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_C_CY;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_C_XOR;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_D;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_D1;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_D2;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_D3;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_D4;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_D5;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_D6;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_DO5;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_DO6;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_D_CY;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_D_XOR;
  wire [0:0] CLBLM_R_X63Y94_SLICE_X95Y94_SR;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_A;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_A1;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_A2;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_A3;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_A4;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_A5;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_A6;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_AI;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_AMUX;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_AO5;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_AO6;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_AX;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_B;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_B1;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_B2;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_B3;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_B4;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_B5;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_B6;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_BO5;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_BO6;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_BX;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_C;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_C1;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_C2;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_C3;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_C4;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_C5;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_C6;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_CE;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_CLK;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_CO5;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_CO6;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_CX;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_D;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_D1;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_D2;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_D3;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_D4;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_D5;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_D6;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_DI;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_DO5;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_DO6;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X94Y95_DX;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_A;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_A1;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_A2;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_A3;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_A4;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_A5;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_A6;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_AMUX;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_AO5;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_AO6;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_AQ;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_AX;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_A_CY;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_A_XOR;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_B;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_B1;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_B2;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_B3;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_B4;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_B5;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_B5Q;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_B6;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_BMUX;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_BO5;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_BO6;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_BQ;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_BX;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_B_CY;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_B_XOR;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_C;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_C1;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_C2;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_C3;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_C4;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_C5;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_C5Q;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_C6;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_CE;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_CLK;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_CMUX;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_CO5;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_CO6;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_CQ;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_CX;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_C_CY;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_C_XOR;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_D;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_D1;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_D2;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_D3;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_D4;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_D5;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_D5Q;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_D6;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_DMUX;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_DO5;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_DO6;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_DQ;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_DX;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_D_CY;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_D_XOR;
  wire [0:0] CLBLM_R_X63Y95_SLICE_X95Y95_SR;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_A;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_A1;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_A2;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_A3;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_A4;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_A5;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_A6;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_AI;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_AMUX;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_AO5;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_AO6;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_AX;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_B;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_B1;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_B2;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_B3;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_B4;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_B5;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_B6;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_BI;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_BMUX;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_BO5;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_BO6;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_BX;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_C;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_C1;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_C2;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_C3;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_C4;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_C5;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_C6;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_CE;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_CI;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_CLK;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_CMUX;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_CO5;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_CO6;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_CX;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_D;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_D1;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_D2;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_D3;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_D4;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_D5;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_D6;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_DI;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_DO5;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_DO6;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X94Y96_DX;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_A;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_A1;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_A2;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_A3;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_A4;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_A5;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_A6;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_AMUX;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_AO5;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_AO6;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_AQ;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_AX;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_A_CY;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_A_XOR;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_B;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_B1;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_B2;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_B3;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_B4;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_B5;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_B6;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_BO5;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_BO6;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_BQ;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_B_CY;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_B_XOR;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_C;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_C1;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_C2;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_C3;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_C4;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_C5;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_C6;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_CE;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_CLK;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_CO5;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_CO6;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_C_CY;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_C_XOR;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_D;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_D1;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_D2;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_D3;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_D4;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_D5;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_D6;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_DO5;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_DO6;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_D_CY;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_D_XOR;
  wire [0:0] CLBLM_R_X63Y96_SLICE_X95Y96_SR;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_A;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_A1;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_A2;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_A3;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_A4;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_A5;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_A6;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_AMUX;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_AO5;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_AO6;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_AX;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_A_CY;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_A_XOR;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_B;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_B1;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_B2;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_B3;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_B4;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_B5;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_B6;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_BO5;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_BO6;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_BQ;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_BX;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_B_CY;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_B_XOR;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_C;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_C1;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_C2;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_C3;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_C4;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_C5;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_C6;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_CE;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_CLK;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_CMUX;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_CO5;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_CO6;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_CQ;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_CX;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_C_CY;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_C_XOR;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_D;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_D1;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_D2;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_D3;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_D4;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_D5;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_D6;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_DO5;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_DO6;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_DQ;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_D_CY;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_D_XOR;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_F7AMUX_O;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X94Y97_SR;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_A;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_A1;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_A2;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_A3;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_A4;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_A5;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_A6;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_AMUX;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_AO5;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_AO6;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_AX;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_A_CY;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_A_XOR;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_B;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_B1;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_B2;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_B3;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_B4;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_B5;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_B6;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_BO5;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_BO6;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_B_CY;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_B_XOR;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_C;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_C1;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_C2;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_C3;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_C4;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_C5;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_C5Q;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_C6;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_CE;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_CLK;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_CMUX;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_CO5;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_CO6;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_CQ;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_C_CY;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_C_XOR;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_D;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_D1;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_D2;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_D3;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_D4;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_D5;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_D5Q;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_D6;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_DMUX;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_DO5;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_DO6;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_DQ;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_D_CY;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_D_XOR;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_F7AMUX_O;
  wire [0:0] CLBLM_R_X63Y97_SLICE_X95Y97_SR;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_A;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_A1;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_A2;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_A3;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_A4;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_A5;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_A6;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_AMUX;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_AO5;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_AO6;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_AX;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_A_CY;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_A_XOR;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_B;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_B1;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_B2;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_B3;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_B4;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_B5;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_B6;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_BO5;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_BO6;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_B_CY;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_B_XOR;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_C;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_C1;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_C2;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_C3;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_C4;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_C5;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_C5Q;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_C6;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_CE;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_CLK;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_CMUX;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_CO5;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_CO6;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_CQ;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_C_CY;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_C_XOR;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_D;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_D1;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_D2;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_D3;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_D4;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_D5;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_D6;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_DO5;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_DO6;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_D_CY;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_D_XOR;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_F7AMUX_O;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X94Y98_SR;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_A;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_A1;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_A2;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_A3;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_A4;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_A5;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_A5Q;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_A6;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_AMUX;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_AO5;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_AO6;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_AQ;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_A_CY;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_A_XOR;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_B;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_B1;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_B2;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_B3;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_B4;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_B5;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_B5Q;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_B6;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_BMUX;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_BO5;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_BO6;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_BQ;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_B_CY;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_B_XOR;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_C;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_C1;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_C2;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_C3;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_C4;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_C5;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_C5Q;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_C6;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_CE;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_CLK;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_CMUX;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_CO5;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_CO6;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_CQ;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_C_CY;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_C_XOR;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_D;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_D1;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_D2;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_D3;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_D4;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_D5;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_D5Q;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_D6;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_DMUX;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_DO5;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_DO6;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_DQ;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_D_CY;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_D_XOR;
  wire [0:0] CLBLM_R_X63Y98_SLICE_X95Y98_SR;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_A;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_A1;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_A2;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_A3;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_A4;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_A5;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_A6;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_AMUX;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_AO5;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_AO6;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_AX;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_A_CY;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_A_XOR;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_B;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_B1;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_B2;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_B3;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_B4;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_B5;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_B6;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_BO5;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_BO6;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_B_CY;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_B_XOR;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_C;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_C1;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_C2;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_C3;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_C4;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_C5;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_C5Q;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_C6;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_CE;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_CLK;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_CMUX;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_CO5;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_CO6;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_CQ;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_C_CY;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_C_XOR;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_D;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_D1;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_D2;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_D3;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_D4;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_D5;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_D6;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_DMUX;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_DO5;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_DO6;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_D_CY;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_D_XOR;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_F7AMUX_O;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X94Y99_SR;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_A;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_A1;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_A2;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_A3;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_A4;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_A5;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_A5Q;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_A6;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_AMUX;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_AO5;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_AO6;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_AQ;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_A_CY;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_A_XOR;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_B;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_B1;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_B2;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_B3;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_B4;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_B5;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_B5Q;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_B6;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_BMUX;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_BO5;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_BO6;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_BQ;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_B_CY;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_B_XOR;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_C;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_C1;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_C2;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_C3;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_C4;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_C5;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_C5Q;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_C6;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_CE;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_CLK;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_CMUX;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_CO5;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_CO6;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_CQ;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_C_CY;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_C_XOR;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_D;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_D1;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_D2;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_D3;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_D4;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_D5;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_D6;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_DO5;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_DO6;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_D_CY;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_D_XOR;
  wire [0:0] CLBLM_R_X63Y99_SLICE_X95Y99_SR;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_A;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_A1;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_A2;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_A3;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_A4;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_A5;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_A6;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_AO5;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_AO6;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_AX;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_A_CY;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_A_XOR;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_B;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_B1;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_B2;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_B3;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_B4;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_B5;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_B6;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_BMUX;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_BO5;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_BO6;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_BX;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_B_CY;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_B_XOR;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_C;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_C1;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_C2;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_C3;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_C4;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_C5;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_C6;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_CMUX;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_CO5;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_CO6;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_COUT;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_CX;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_C_CY;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_C_XOR;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_D;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_D1;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_D2;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_D3;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_D4;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_D5;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_D6;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_DMUX;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_DO5;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_DO6;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_DX;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_D_CY;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X98Y100_D_XOR;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_A;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_A1;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_A2;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_A3;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_A4;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_A5;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_A6;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_AO5;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_AO6;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_AQ;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_A_CY;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_A_XOR;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_B;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_B1;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_B2;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_B3;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_B4;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_B5;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_B6;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_BO5;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_BO6;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_BQ;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_B_CY;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_B_XOR;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_C;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_C1;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_C2;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_C3;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_C4;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_C5;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_C6;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_CE;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_CLK;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_CO5;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_CO6;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_CQ;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_C_CY;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_C_XOR;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_D;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_D1;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_D2;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_D3;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_D4;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_D5;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_D6;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_DO5;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_DO6;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_D_CY;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_D_XOR;
  wire [0:0] CLBLM_R_X65Y100_SLICE_X99Y100_SR;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_A;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_A1;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_A2;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_A3;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_A4;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_A5;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_A6;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_AMUX;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_AO5;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_AO6;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_AX;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_A_CY;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_A_XOR;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_B;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_B1;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_B2;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_B3;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_B4;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_B5;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_B6;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_BMUX;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_BO5;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_BO6;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_BX;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_B_CY;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_B_XOR;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_C;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_C1;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_C2;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_C3;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_C4;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_C5;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_C6;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_CIN;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_CMUX;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_CO5;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_CO6;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_COUT;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_CX;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_C_CY;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_C_XOR;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_D;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_D1;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_D2;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_D3;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_D4;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_D5;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_D6;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_DMUX;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_DO5;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_DO6;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_DX;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_D_CY;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X98Y101_D_XOR;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_A;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_A1;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_A2;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_A3;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_A4;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_A5;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_A6;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_AO5;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_AO6;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_AQ;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_A_CY;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_A_XOR;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_B;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_B1;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_B2;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_B3;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_B4;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_B5;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_B6;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_BO5;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_BO6;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_B_CY;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_B_XOR;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_C;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_C1;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_C2;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_C3;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_C4;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_C5;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_C6;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_CE;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_CLK;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_CO5;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_CO6;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_C_CY;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_C_XOR;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_D;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_D1;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_D2;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_D3;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_D4;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_D5;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_D6;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_DO5;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_DO6;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_D_CY;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_D_XOR;
  wire [0:0] CLBLM_R_X65Y101_SLICE_X99Y101_SR;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_A;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_A1;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_A2;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_A3;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_A4;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_A5;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_A6;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_AMUX;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_AO5;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_AO6;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_A_CY;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_A_XOR;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_B;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_B1;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_B2;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_B3;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_B4;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_B5;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_B6;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_BMUX;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_BO5;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_BO6;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_BX;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_B_CY;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_B_XOR;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_C;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_C1;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_C2;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_C3;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_C4;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_C5;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_C6;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_CIN;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_CMUX;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_CO5;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_CO6;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_COUT;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_CX;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_C_CY;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_C_XOR;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_D;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_D1;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_D2;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_D3;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_D4;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_D5;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_D6;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_DMUX;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_DO5;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_DO6;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_DX;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_D_CY;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X98Y102_D_XOR;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_A;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_A1;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_A2;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_A3;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_A4;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_A5;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_A6;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_AO5;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_AO6;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_AQ;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_A_CY;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_A_XOR;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_B;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_B1;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_B2;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_B3;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_B4;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_B5;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_B6;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_BO5;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_BO6;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_B_CY;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_B_XOR;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_C;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_C1;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_C2;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_C3;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_C4;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_C5;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_C6;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_CE;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_CLK;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_CO5;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_CO6;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_C_CY;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_C_XOR;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_D;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_D1;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_D2;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_D3;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_D4;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_D5;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_D6;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_DO5;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_DO6;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_D_CY;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_D_XOR;
  wire [0:0] CLBLM_R_X65Y102_SLICE_X99Y102_SR;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_A;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_A1;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_A2;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_A3;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_A4;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_A5;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_A6;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_AMUX;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_AO5;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_AO6;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_AX;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_A_CY;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_A_XOR;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_B;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_B1;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_B2;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_B3;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_B4;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_B5;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_B6;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_BMUX;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_BO5;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_BO6;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_BX;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_B_CY;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_B_XOR;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_C;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_C1;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_C2;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_C3;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_C4;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_C5;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_C6;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_CIN;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_CMUX;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_CO5;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_CO6;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_COUT;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_CX;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_C_CY;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_C_XOR;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_D;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_D1;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_D2;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_D3;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_D4;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_D5;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_D6;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_DMUX;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_DO5;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_DO6;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_DX;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_D_CY;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X98Y103_D_XOR;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_A;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_A1;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_A2;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_A3;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_A4;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_A5;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_A6;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_AO5;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_AO6;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_AQ;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_A_CY;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_A_XOR;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_B;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_B1;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_B2;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_B3;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_B4;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_B5;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_B6;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_BO5;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_BO6;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_BQ;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_B_CY;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_B_XOR;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_C;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_C1;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_C2;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_C3;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_C4;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_C5;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_C6;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_CE;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_CLK;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_CMUX;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_CO5;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_CO6;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_C_CY;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_C_XOR;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_D;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_D1;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_D2;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_D3;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_D4;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_D5;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_D6;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_DO5;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_DO6;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_D_CY;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_D_XOR;
  wire [0:0] CLBLM_R_X65Y103_SLICE_X99Y103_SR;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_A;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_A1;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_A2;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_A3;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_A4;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_A5;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_A6;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_AMUX;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_AO5;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_AO6;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_AX;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_A_CY;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_A_XOR;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_B;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_B1;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_B2;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_B3;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_B4;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_B5;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_B6;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_BMUX;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_BO5;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_BO6;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_BX;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_B_CY;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_B_XOR;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_C;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_C1;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_C2;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_C3;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_C4;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_C5;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_C6;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_CIN;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_CMUX;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_CO5;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_CO6;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_COUT;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_CX;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_C_CY;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_C_XOR;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_D;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_D1;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_D2;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_D3;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_D4;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_D5;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_D6;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_DO5;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_DO6;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_DX;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_D_CY;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X98Y104_D_XOR;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_A;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_A1;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_A2;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_A3;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_A4;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_A5;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_A6;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_AO5;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_AO6;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_AQ;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_A_CY;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_A_XOR;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_B;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_B1;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_B2;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_B3;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_B4;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_B5;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_B6;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_BO5;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_BO6;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_BQ;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_B_CY;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_B_XOR;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_C;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_C1;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_C2;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_C3;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_C4;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_C5;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_C6;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_CE;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_CLK;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_CO5;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_CO6;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_C_CY;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_C_XOR;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_D;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_D1;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_D2;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_D3;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_D4;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_D5;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_D6;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_DO5;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_DO6;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_D_CY;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_D_XOR;
  wire [0:0] CLBLM_R_X65Y104_SLICE_X99Y104_SR;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_A;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_A1;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_A2;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_A3;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_A4;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_A5;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_A6;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_AO5;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_AO6;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_AQ;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_A_CY;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_A_XOR;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_B;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_B1;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_B2;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_B3;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_B4;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_B5;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_B6;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_BO5;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_BO6;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_BQ;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_B_CY;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_B_XOR;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_C;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_C1;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_C2;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_C3;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_C4;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_C5;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_C6;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_CE;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_CLK;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_CO5;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_CO6;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_C_CY;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_C_XOR;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_D;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_D1;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_D2;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_D3;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_D4;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_D5;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_D6;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_DO5;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_DO6;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_D_CY;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_D_XOR;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X98Y105_SR;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_A;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_A1;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_A2;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_A3;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_A4;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_A5;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_A6;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_AO5;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_AO6;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_AQ;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_A_CY;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_A_XOR;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_B;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_B1;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_B2;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_B3;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_B4;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_B5;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_B6;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_BO5;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_BO6;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_B_CY;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_B_XOR;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_C;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_C1;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_C2;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_C3;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_C4;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_C5;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_C6;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_CE;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_CLK;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_CO5;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_CO6;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_C_CY;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_C_XOR;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_D;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_D1;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_D2;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_D3;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_D4;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_D5;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_D6;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_DO5;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_DO6;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_D_CY;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_D_XOR;
  wire [0:0] CLBLM_R_X65Y105_SLICE_X99Y105_SR;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_A;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_A1;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_A2;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_A3;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_A4;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_A5;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_A6;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_AO5;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_AO6;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_AQ;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_A_CY;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_A_XOR;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_B;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_B1;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_B2;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_B3;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_B4;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_B5;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_B6;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_BO5;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_BO6;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_BQ;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_B_CY;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_B_XOR;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_C;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_C1;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_C2;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_C3;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_C4;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_C5;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_C6;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_CE;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_CLK;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_CO5;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_CO6;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_CQ;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_C_CY;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_C_XOR;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_D;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_D1;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_D2;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_D3;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_D4;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_D5;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_D6;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_DO5;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_DO6;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_DQ;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_D_CY;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_D_XOR;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X98Y106_SR;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_A;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_A1;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_A2;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_A3;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_A4;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_A5;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_A6;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_AO5;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_AO6;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_A_CY;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_A_XOR;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_B;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_B1;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_B2;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_B3;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_B4;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_B5;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_B6;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_BO5;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_BO6;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_B_CY;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_B_XOR;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_C;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_C1;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_C2;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_C3;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_C4;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_C5;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_C6;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_CO5;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_CO6;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_C_CY;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_C_XOR;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_D;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_D1;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_D2;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_D3;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_D4;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_D5;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_D6;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_DO5;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_DO6;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_D_CY;
  wire [0:0] CLBLM_R_X65Y106_SLICE_X99Y106_D_XOR;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_A;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_A1;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_A2;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_A3;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_A4;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_A5;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_A6;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_AO5;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_AO6;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_AQ;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_A_CY;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_A_XOR;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_B;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_B1;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_B2;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_B3;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_B4;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_B5;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_B6;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_BO5;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_BO6;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_BQ;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_B_CY;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_B_XOR;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_C;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_C1;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_C2;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_C3;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_C4;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_C5;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_C6;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_CE;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_CLK;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_CO5;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_CO6;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_CQ;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_C_CY;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_C_XOR;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_D;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_D1;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_D2;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_D3;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_D4;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_D5;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_D6;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_DO5;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_DO6;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_DQ;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_D_CY;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_D_XOR;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X98Y107_SR;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_A;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_A1;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_A2;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_A3;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_A4;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_A5;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_A6;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_AO5;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_AO6;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_A_CY;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_A_XOR;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_B;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_B1;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_B2;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_B3;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_B4;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_B5;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_B6;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_BO5;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_BO6;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_B_CY;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_B_XOR;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_C;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_C1;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_C2;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_C3;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_C4;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_C5;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_C6;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_CO5;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_CO6;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_C_CY;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_C_XOR;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_D;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_D1;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_D2;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_D3;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_D4;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_D5;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_D6;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_DO5;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_DO6;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_D_CY;
  wire [0:0] CLBLM_R_X65Y107_SLICE_X99Y107_D_XOR;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_A;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_A1;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_A2;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_A3;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_A4;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_A5;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_A6;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_AO5;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_AO6;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_A_CY;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_A_XOR;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_B;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_B1;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_B2;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_B3;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_B4;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_B5;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_B6;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_BO5;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_BO6;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_B_CY;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_B_XOR;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_C;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_C1;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_C2;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_C3;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_C4;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_C5;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_C6;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_CO5;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_CO6;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_C_CY;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_C_XOR;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_D;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_D1;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_D2;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_D3;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_D4;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_D5;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_D6;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_DO5;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_DO6;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_D_CY;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X98Y96_D_XOR;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_A;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_A1;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_A2;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_A3;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_A4;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_A5;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_A6;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_AO5;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_AO6;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_A_CY;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_A_XOR;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_B;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_B1;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_B2;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_B3;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_B4;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_B5;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_B6;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_BO5;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_BO6;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_B_CY;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_B_XOR;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_C;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_C1;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_C2;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_C3;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_C4;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_C5;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_C6;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_CO5;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_CO6;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_C_CY;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_C_XOR;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_D;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_D1;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_D2;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_D3;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_D4;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_D5;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_D6;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_DO5;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_DO6;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_D_CY;
  wire [0:0] CLBLM_R_X65Y96_SLICE_X99Y96_D_XOR;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_A;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_A1;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_A2;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_A3;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_A4;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_A5;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_A6;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_AMUX;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_AO5;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_AO6;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_A_CY;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_A_XOR;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_B;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_B1;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_B2;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_B3;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_B4;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_B5;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_B6;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_BO5;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_BO6;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_B_CY;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_B_XOR;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_C;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_C1;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_C2;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_C3;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_C4;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_C5;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_C6;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_CO5;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_CO6;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_C_CY;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_C_XOR;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_D;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_D1;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_D2;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_D3;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_D4;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_D5;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_D6;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_DO5;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_DO6;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_D_CY;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X98Y97_D_XOR;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_A;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_A1;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_A2;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_A3;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_A4;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_A5;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_A6;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_AO5;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_AO6;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_A_CY;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_A_XOR;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_B;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_B1;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_B2;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_B3;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_B4;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_B5;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_B6;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_BO5;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_BO6;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_B_CY;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_B_XOR;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_C;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_C1;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_C2;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_C3;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_C4;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_C5;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_C6;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_CO5;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_CO6;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_C_CY;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_C_XOR;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_D;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_D1;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_D2;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_D3;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_D4;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_D5;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_D6;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_DO5;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_DO6;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_D_CY;
  wire [0:0] CLBLM_R_X65Y97_SLICE_X99Y97_D_XOR;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_A;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_A1;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_A2;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_A3;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_A4;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_A5;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_A6;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_AO5;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_AO6;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_AQ;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_A_CY;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_A_XOR;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_B;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_B1;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_B2;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_B3;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_B4;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_B5;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_B6;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_BO5;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_BO6;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_BQ;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_B_CY;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_B_XOR;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_C;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_C1;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_C2;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_C3;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_C4;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_C5;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_C6;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_CE;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_CLK;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_CMUX;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_CO5;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_CO6;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_C_CY;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_C_XOR;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_D;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_D1;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_D2;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_D3;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_D4;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_D5;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_D6;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_DO5;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_DO6;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_D_CY;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_D_XOR;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X98Y98_SR;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_A;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_A1;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_A2;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_A3;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_A4;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_A5;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_A6;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_AO5;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_AO6;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_AQ;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_A_CY;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_A_XOR;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_B;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_B1;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_B2;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_B3;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_B4;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_B5;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_B6;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_BO5;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_BO6;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_B_CY;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_B_XOR;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_C;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_C1;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_C2;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_C3;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_C4;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_C5;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_C6;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_CE;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_CLK;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_CO5;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_CO6;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_C_CY;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_C_XOR;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_D;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_D1;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_D2;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_D3;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_D4;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_D5;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_D6;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_DO5;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_DO6;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_D_CY;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_D_XOR;
  wire [0:0] CLBLM_R_X65Y98_SLICE_X99Y98_SR;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_A;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_A1;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_A2;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_A3;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_A4;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_A5;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_A6;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_AO5;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_AO6;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_AQ;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_A_CY;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_A_XOR;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_B;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_B1;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_B2;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_B3;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_B4;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_B5;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_B6;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_BO5;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_BO6;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_B_CY;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_B_XOR;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_C;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_C1;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_C2;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_C3;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_C4;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_C5;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_C6;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_CE;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_CLK;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_CO5;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_CO6;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_C_CY;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_C_XOR;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_D;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_D1;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_D2;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_D3;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_D4;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_D5;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_D6;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_DO5;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_DO6;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_D_CY;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_D_XOR;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X98Y99_SR;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_A;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_A1;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_A2;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_A3;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_A4;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_A5;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_A6;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_AO5;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_AO6;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_AQ;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_A_CY;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_A_XOR;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_B;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_B1;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_B2;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_B3;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_B4;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_B5;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_B6;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_BO5;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_BO6;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_B_CY;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_B_XOR;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_C;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_C1;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_C2;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_C3;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_C4;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_C5;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_C6;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_CE;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_CLK;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_CO5;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_CO6;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_C_CY;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_C_XOR;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_D;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_D1;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_D2;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_D3;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_D4;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_D5;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_D6;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_DO5;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_DO6;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_D_CY;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_D_XOR;
  wire [0:0] CLBLM_R_X65Y99_SLICE_X99Y99_SR;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_CE;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_I;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  wire [0:0] CLK_HROW_BOT_R_X139Y78_BUFHCE_X0Y20_CE;
  wire [0:0] CLK_HROW_BOT_R_X139Y78_BUFHCE_X0Y20_I;
  wire [0:0] CLK_HROW_BOT_R_X139Y78_BUFHCE_X0Y20_O;
  wire [0:0] CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_CE;
  wire [0:0] CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_I;
  wire [0:0] CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_I;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_I;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_I;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_I;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_I;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_I;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_I;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_O;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_O;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_D;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_O;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y119_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y119_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_O;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_O;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_D;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_O;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y118_D;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y118_O;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y121_D;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y121_O;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y122_D;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y122_O;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y123_D;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y123_O;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_TQ;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_O;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_O;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_O;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_O;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_O;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_O;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_O;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y114_O;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y115_O;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y116_O;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y117_O;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y118_O;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y119_O;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y120_O;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y121_O;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y122_O;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y123_O;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y124_O;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y125_O;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y126_O;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y127_O;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y128_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y129_O;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y130_O;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y131_O;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y132_O;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y133_O;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y134_O;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y135_O;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y136_O;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y137_O;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y138_O;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y139_O;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y140_O;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y141_O;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y142_O;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y143_O;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y144_O;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y145_O;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_D;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_TQ;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_O;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y109_D1;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y109_OQ;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y109_T1;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y109_TQ;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y110_D1;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y110_OQ;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y110_T1;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y110_TQ;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y111_D1;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y111_OQ;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y111_T1;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y111_TQ;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y112_D1;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y112_OQ;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y112_T1;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y112_TQ;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y115_D1;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y115_OQ;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y115_T1;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y115_TQ;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y116_D1;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y116_OQ;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y116_T1;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y116_TQ;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y117_D1;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y117_OQ;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y117_T1;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y117_TQ;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y118_D1;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y118_OQ;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y118_T1;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y118_TQ;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y121_D1;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y121_OQ;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y121_T1;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y121_TQ;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y122_D1;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y122_OQ;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y122_T1;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y122_TQ;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y123_D1;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y123_OQ;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y123_T1;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y123_TQ;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y124_D1;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y124_OQ;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y124_T1;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y124_TQ;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y125_D1;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y125_OQ;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y125_T1;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y125_TQ;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y126_D1;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y126_OQ;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y126_T1;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y126_TQ;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_O;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_D1;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_OQ;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_T1;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_TQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_D1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_OQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_T1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_TQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_D1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_OQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_T1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_TQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_D1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_OQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_T1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_TQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_D1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_OQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_T1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_TQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_D1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_OQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_T1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_TQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_D1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_OQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_T1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_TQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_D1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_OQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_T1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_TQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_D1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_OQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_T1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_TQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_D1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_OQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_T1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_TQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_D1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_OQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_T1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_TQ;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_D1;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_OQ;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_T1;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_TQ;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y99_SLICE_X78Y99_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y99_SLICE_X78Y99_DO5),
.O6(CLBLL_L_X52Y99_SLICE_X78Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y99_SLICE_X78Y99_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y99_SLICE_X78Y99_CO5),
.O6(CLBLL_L_X52Y99_SLICE_X78Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y99_SLICE_X78Y99_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y99_SLICE_X78Y99_BO5),
.O6(CLBLL_L_X52Y99_SLICE_X78Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0022010001000002)
  ) CLBLL_L_X52Y99_SLICE_X78Y99_ALUT (
.I0(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.I1(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I2(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.I3(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.I4(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.I5(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.O5(CLBLL_L_X52Y99_SLICE_X78Y99_AO5),
.O6(CLBLL_L_X52Y99_SLICE_X78Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0040000000000100)
  ) CLBLL_L_X52Y99_SLICE_X79Y99_DLUT (
.I0(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I1(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.I2(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.I3(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.I4(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.I5(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.O5(CLBLL_L_X52Y99_SLICE_X79Y99_DO5),
.O6(CLBLL_L_X52Y99_SLICE_X79Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000040000004000)
  ) CLBLL_L_X52Y99_SLICE_X79Y99_CLUT (
.I0(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I1(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.I2(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.I3(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.I4(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.I5(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.O5(CLBLL_L_X52Y99_SLICE_X79Y99_CO5),
.O6(CLBLL_L_X52Y99_SLICE_X79Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha330073003300330)
  ) CLBLL_L_X52Y99_SLICE_X79Y99_BLUT (
.I0(CLBLM_R_X49Y108_SLICE_X75Y108_DQ),
.I1(CLBLM_R_X53Y99_SLICE_X80Y99_AO6),
.I2(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.I3(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I4(CLBLM_R_X49Y107_SLICE_X75Y107_DQ),
.I5(CLBLM_L_X56Y97_SLICE_X84Y97_CO5),
.O5(CLBLL_L_X52Y99_SLICE_X79Y99_BO5),
.O6(CLBLL_L_X52Y99_SLICE_X79Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffba)
  ) CLBLL_L_X52Y99_SLICE_X79Y99_ALUT (
.I0(CLBLL_L_X52Y99_SLICE_X79Y99_DO6),
.I1(CLBLM_R_X53Y99_SLICE_X80Y99_AO5),
.I2(CLBLM_L_X56Y97_SLICE_X84Y97_AO6),
.I3(CLBLL_L_X52Y99_SLICE_X79Y99_BO6),
.I4(CLBLL_L_X52Y101_SLICE_X79Y101_AO6),
.I5(CLBLL_L_X52Y99_SLICE_X79Y99_CO6),
.O5(CLBLL_L_X52Y99_SLICE_X79Y99_AO5),
.O6(CLBLL_L_X52Y99_SLICE_X79Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y101_SLICE_X78Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y101_SLICE_X78Y101_DO5),
.O6(CLBLL_L_X52Y101_SLICE_X78Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y101_SLICE_X78Y101_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y101_SLICE_X78Y101_CO5),
.O6(CLBLL_L_X52Y101_SLICE_X78Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y101_SLICE_X78Y101_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y101_SLICE_X78Y101_BO5),
.O6(CLBLL_L_X52Y101_SLICE_X78Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y101_SLICE_X78Y101_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y101_SLICE_X78Y101_AO5),
.O6(CLBLL_L_X52Y101_SLICE_X78Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y101_SLICE_X79Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y101_SLICE_X79Y101_DO5),
.O6(CLBLL_L_X52Y101_SLICE_X79Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y101_SLICE_X79Y101_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y101_SLICE_X79Y101_CO5),
.O6(CLBLL_L_X52Y101_SLICE_X79Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y101_SLICE_X79Y101_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y101_SLICE_X79Y101_BO5),
.O6(CLBLL_L_X52Y101_SLICE_X79Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000010000)
  ) CLBLL_L_X52Y101_SLICE_X79Y101_ALUT (
.I0(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.I1(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.I2(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I3(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I4(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.I5(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.O5(CLBLL_L_X52Y101_SLICE_X79Y101_AO5),
.O6(CLBLL_L_X52Y101_SLICE_X79Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y105_SLICE_X78Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y105_SLICE_X78Y105_DO5),
.O6(CLBLL_L_X52Y105_SLICE_X78Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf500ffffe400ffff)
  ) CLBLL_L_X52Y105_SLICE_X78Y105_CLUT (
.I0(CLBLM_R_X53Y101_SLICE_X80Y101_BQ),
.I1(CLBLL_L_X52Y106_SLICE_X78Y106_AO5),
.I2(CLBLL_R_X57Y97_SLICE_X86Y97_AQ),
.I3(CLBLL_L_X52Y105_SLICE_X78Y105_AO5),
.I4(CLBLM_R_X53Y101_SLICE_X81Y101_AQ),
.I5(CLBLL_R_X57Y99_SLICE_X86Y99_BQ),
.O5(CLBLL_L_X52Y105_SLICE_X78Y105_CO5),
.O6(CLBLL_L_X52Y105_SLICE_X78Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0000ff0f0f)
  ) CLBLL_L_X52Y105_SLICE_X78Y105_BLUT (
.I0(CLBLL_R_X57Y100_SLICE_X86Y100_BQ),
.I1(1'b1),
.I2(CLBLL_R_X57Y100_SLICE_X86Y100_DQ),
.I3(CLBLM_L_X56Y101_SLICE_X85Y101_CQ),
.I4(CLBLL_L_X54Y100_SLICE_X82Y100_BQ),
.I5(1'b1),
.O5(CLBLL_L_X52Y105_SLICE_X78Y105_BO5),
.O6(CLBLL_L_X52Y105_SLICE_X78Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8080a0000000aaaa)
  ) CLBLL_L_X52Y105_SLICE_X78Y105_ALUT (
.I0(CLBLM_R_X53Y100_SLICE_X81Y100_AQ),
.I1(CLBLL_R_X57Y100_SLICE_X86Y100_DQ),
.I2(CLBLM_R_X53Y101_SLICE_X80Y101_BQ),
.I3(CLBLL_R_X57Y99_SLICE_X86Y99_BQ),
.I4(CLBLL_L_X54Y100_SLICE_X82Y100_BQ),
.I5(1'b1),
.O5(CLBLL_L_X52Y105_SLICE_X78Y105_AO5),
.O6(CLBLL_L_X52Y105_SLICE_X78Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y105_SLICE_X79Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y105_SLICE_X79Y105_DO5),
.O6(CLBLL_L_X52Y105_SLICE_X79Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y105_SLICE_X79Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y105_SLICE_X79Y105_CO5),
.O6(CLBLL_L_X52Y105_SLICE_X79Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y105_SLICE_X79Y105_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y105_SLICE_X79Y105_BO5),
.O6(CLBLL_L_X52Y105_SLICE_X79Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y105_SLICE_X79Y105_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y105_SLICE_X79Y105_AO5),
.O6(CLBLL_L_X52Y105_SLICE_X79Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y106_SLICE_X78Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y106_SLICE_X78Y106_DO5),
.O6(CLBLL_L_X52Y106_SLICE_X78Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y106_SLICE_X78Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y106_SLICE_X78Y106_CO5),
.O6(CLBLL_L_X52Y106_SLICE_X78Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y106_SLICE_X78Y106_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y106_SLICE_X78Y106_BO5),
.O6(CLBLL_L_X52Y106_SLICE_X78Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000fffafffa)
  ) CLBLL_L_X52Y106_SLICE_X78Y106_ALUT (
.I0(CLBLM_L_X50Y106_SLICE_X76Y106_BO5),
.I1(1'b1),
.I2(CLBLL_R_X57Y101_SLICE_X87Y101_DQ),
.I3(CLBLM_L_X56Y101_SLICE_X85Y101_DQ),
.I4(CLBLL_R_X57Y99_SLICE_X86Y99_AQ),
.I5(1'b1),
.O5(CLBLL_L_X52Y106_SLICE_X78Y106_AO5),
.O6(CLBLL_L_X52Y106_SLICE_X78Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y106_SLICE_X79Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y106_SLICE_X79Y106_DO5),
.O6(CLBLL_L_X52Y106_SLICE_X79Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y106_SLICE_X79Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y106_SLICE_X79Y106_CO5),
.O6(CLBLL_L_X52Y106_SLICE_X79Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aaaaaaff000000)
  ) CLBLL_L_X52Y106_SLICE_X79Y106_BLUT (
.I0(CLBLL_R_X57Y101_SLICE_X87Y101_CQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X56Y101_SLICE_X85Y101_DQ),
.I4(CLBLL_R_X57Y100_SLICE_X86Y100_AQ),
.I5(CLBLL_R_X57Y100_SLICE_X86Y100_BQ),
.O5(CLBLL_L_X52Y106_SLICE_X79Y106_BO5),
.O6(CLBLL_L_X52Y106_SLICE_X79Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0fe329292)
  ) CLBLL_L_X52Y106_SLICE_X79Y106_ALUT (
.I0(CLBLL_R_X57Y101_SLICE_X87Y101_CQ),
.I1(CLBLL_L_X54Y100_SLICE_X82Y100_BQ),
.I2(CLBLL_R_X57Y101_SLICE_X87Y101_AQ),
.I3(CLBLL_R_X57Y100_SLICE_X86Y100_DQ),
.I4(CLBLM_R_X53Y101_SLICE_X80Y101_BQ),
.I5(1'b1),
.O5(CLBLL_L_X52Y106_SLICE_X79Y106_AO5),
.O6(CLBLL_L_X52Y106_SLICE_X79Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y107_SLICE_X78Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y107_SLICE_X78Y107_DO5),
.O6(CLBLL_L_X52Y107_SLICE_X78Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y107_SLICE_X78Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y107_SLICE_X78Y107_CO5),
.O6(CLBLL_L_X52Y107_SLICE_X78Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000acf3a0cc)
  ) CLBLL_L_X52Y107_SLICE_X78Y107_BLUT (
.I0(CLBLM_L_X56Y101_SLICE_X85Y101_CQ),
.I1(CLBLL_R_X57Y100_SLICE_X87Y100_BQ),
.I2(CLBLM_R_X53Y101_SLICE_X80Y101_BQ),
.I3(CLBLL_L_X54Y100_SLICE_X82Y100_BQ),
.I4(CLBLL_R_X57Y101_SLICE_X87Y101_DQ),
.I5(1'b1),
.O5(CLBLL_L_X52Y107_SLICE_X78Y107_BO5),
.O6(CLBLL_L_X52Y107_SLICE_X78Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00f9e23922)
  ) CLBLL_L_X52Y107_SLICE_X78Y107_ALUT (
.I0(CLBLM_L_X56Y101_SLICE_X85Y101_DQ),
.I1(CLBLL_L_X54Y100_SLICE_X82Y100_BQ),
.I2(CLBLM_R_X53Y101_SLICE_X80Y101_BQ),
.I3(CLBLM_L_X56Y101_SLICE_X85Y101_BQ),
.I4(CLBLL_R_X57Y100_SLICE_X86Y100_CQ),
.I5(1'b1),
.O5(CLBLL_L_X52Y107_SLICE_X78Y107_AO5),
.O6(CLBLL_L_X52Y107_SLICE_X78Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y107_SLICE_X79Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y107_SLICE_X79Y107_DO5),
.O6(CLBLL_L_X52Y107_SLICE_X79Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y107_SLICE_X79Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y107_SLICE_X79Y107_CO5),
.O6(CLBLL_L_X52Y107_SLICE_X79Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y107_SLICE_X79Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y107_SLICE_X79Y107_BO5),
.O6(CLBLL_L_X52Y107_SLICE_X79Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y107_SLICE_X79Y107_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y107_SLICE_X79Y107_AO5),
.O6(CLBLL_L_X52Y107_SLICE_X79Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y97_SLICE_X82Y97_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y97_SLICE_X82Y97_DO5),
.O6(CLBLL_L_X54Y97_SLICE_X82Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y97_SLICE_X82Y97_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y97_SLICE_X82Y97_CO5),
.O6(CLBLL_L_X54Y97_SLICE_X82Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y97_SLICE_X82Y97_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y97_SLICE_X82Y97_BO5),
.O6(CLBLL_L_X54Y97_SLICE_X82Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y97_SLICE_X82Y97_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y97_SLICE_X82Y97_AO5),
.O6(CLBLL_L_X54Y97_SLICE_X82Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y97_SLICE_X83Y97_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y97_SLICE_X83Y97_DO5),
.O6(CLBLL_L_X54Y97_SLICE_X83Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y97_SLICE_X83Y97_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y97_SLICE_X83Y97_CO5),
.O6(CLBLL_L_X54Y97_SLICE_X83Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000002000000000)
  ) CLBLL_L_X54Y97_SLICE_X83Y97_BLUT (
.I0(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.I1(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I2(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.I3(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I4(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.I5(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.O5(CLBLL_L_X54Y97_SLICE_X83Y97_BO5),
.O6(CLBLL_L_X54Y97_SLICE_X83Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0045000000000000)
  ) CLBLL_L_X54Y97_SLICE_X83Y97_ALUT (
.I0(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.I1(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I2(CLBLM_R_X49Y107_SLICE_X75Y107_DQ),
.I3(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I4(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.I5(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.O5(CLBLL_L_X54Y97_SLICE_X83Y97_AO5),
.O6(CLBLL_L_X54Y97_SLICE_X83Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0004000000f00000)
  ) CLBLL_L_X54Y98_SLICE_X82Y98_DLUT (
.I0(CLBLM_R_X49Y107_SLICE_X75Y107_DQ),
.I1(CLBLL_L_X54Y99_SLICE_X83Y99_BO5),
.I2(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I3(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.I4(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.I5(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.O5(CLBLL_L_X54Y98_SLICE_X82Y98_DO5),
.O6(CLBLL_L_X54Y98_SLICE_X82Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0002c0c000000000)
  ) CLBLL_L_X54Y98_SLICE_X82Y98_CLUT (
.I0(CLBLM_R_X49Y107_SLICE_X75Y107_DQ),
.I1(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.I2(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I3(CLBLM_R_X53Y100_SLICE_X81Y100_AO5),
.I4(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.I5(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.O5(CLBLL_L_X54Y98_SLICE_X82Y98_CO5),
.O6(CLBLL_L_X54Y98_SLICE_X82Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000020006040000)
  ) CLBLL_L_X54Y98_SLICE_X82Y98_BLUT (
.I0(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.I1(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.I2(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I3(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.I4(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I5(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.O5(CLBLL_L_X54Y98_SLICE_X82Y98_BO5),
.O6(CLBLL_L_X54Y98_SLICE_X82Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0011001100110010)
  ) CLBLL_L_X54Y98_SLICE_X82Y98_ALUT (
.I0(CLBLL_L_X54Y98_SLICE_X82Y98_BO6),
.I1(CLBLM_R_X53Y100_SLICE_X81Y100_DO6),
.I2(CLBLM_R_X53Y99_SLICE_X80Y99_AO5),
.I3(CLBLM_R_X53Y98_SLICE_X81Y98_AO6),
.I4(CLBLM_R_X49Y107_SLICE_X75Y107_DQ),
.I5(CLBLM_R_X53Y100_SLICE_X81Y100_AO5),
.O5(CLBLL_L_X54Y98_SLICE_X82Y98_AO5),
.O6(CLBLL_L_X54Y98_SLICE_X82Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLL_L_X54Y98_SLICE_X83Y98_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X0Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_L_X54Y98_SLICE_X83Y98_AO6),
.Q(CLBLL_L_X54Y98_SLICE_X83Y98_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLL_L_X54Y98_SLICE_X83Y98_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X0Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_L_X54Y98_SLICE_X83Y98_BO6),
.Q(CLBLL_L_X54Y98_SLICE_X83Y98_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000040000000)
  ) CLBLL_L_X54Y98_SLICE_X83Y98_DLUT (
.I0(CLBLM_R_X49Y107_SLICE_X75Y107_DQ),
.I1(CLBLL_L_X54Y99_SLICE_X83Y99_BO5),
.I2(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I3(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.I4(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.I5(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.O5(CLBLL_L_X54Y98_SLICE_X83Y98_DO5),
.O6(CLBLL_L_X54Y98_SLICE_X83Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffcfcffcfcfcfc)
  ) CLBLL_L_X54Y98_SLICE_X83Y98_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.I2(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I3(1'b1),
.I4(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.I5(1'b1),
.O5(CLBLL_L_X54Y98_SLICE_X83Y98_CO5),
.O6(CLBLL_L_X54Y98_SLICE_X83Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfdfcfcfffdfffc)
  ) CLBLL_L_X54Y98_SLICE_X83Y98_BLUT (
.I0(CLBLM_R_X53Y99_SLICE_X80Y99_AO5),
.I1(CLBLM_R_X53Y99_SLICE_X81Y99_CO6),
.I2(CLBLL_L_X54Y97_SLICE_X83Y97_BO6),
.I3(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.I4(CLBLM_L_X56Y98_SLICE_X84Y98_AO6),
.I5(CLBLL_L_X54Y98_SLICE_X83Y98_CO6),
.O5(CLBLL_L_X54Y98_SLICE_X83Y98_BO5),
.O6(CLBLL_L_X54Y98_SLICE_X83Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffafffefffafffa)
  ) CLBLL_L_X54Y98_SLICE_X83Y98_ALUT (
.I0(CLBLM_R_X53Y99_SLICE_X81Y99_AO6),
.I1(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.I2(CLBLL_L_X54Y97_SLICE_X83Y97_AO6),
.I3(CLBLL_L_X54Y98_SLICE_X82Y98_CO6),
.I4(CLBLL_L_X54Y98_SLICE_X83Y98_CO5),
.I5(CLBLL_L_X54Y99_SLICE_X83Y99_BO5),
.O5(CLBLL_L_X54Y98_SLICE_X83Y98_AO5),
.O6(CLBLL_L_X54Y98_SLICE_X83Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLL_L_X54Y99_SLICE_X82Y99_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X0Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_L_X54Y99_SLICE_X82Y99_BO5),
.Q(CLBLL_L_X54Y99_SLICE_X82Y99_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLL_L_X54Y99_SLICE_X82Y99_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X0Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_L_X54Y99_SLICE_X82Y99_CO6),
.Q(CLBLL_L_X54Y99_SLICE_X82Y99_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3030ffff6068)
  ) CLBLL_L_X54Y99_SLICE_X82Y99_DLUT (
.I0(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.I1(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.I2(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I3(CLBLM_R_X53Y100_SLICE_X81Y100_AO5),
.I4(CLBLM_R_X53Y99_SLICE_X81Y99_AO6),
.I5(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.O5(CLBLL_L_X54Y99_SLICE_X82Y99_DO5),
.O6(CLBLL_L_X54Y99_SLICE_X82Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffefffc)
  ) CLBLL_L_X54Y99_SLICE_X82Y99_CLUT (
.I0(CLBLM_L_X56Y97_SLICE_X84Y97_CO5),
.I1(CLBLM_R_X53Y99_SLICE_X80Y99_DO6),
.I2(CLBLL_L_X54Y99_SLICE_X82Y99_AO5),
.I3(CLBLL_L_X54Y98_SLICE_X82Y98_DO6),
.I4(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I5(CLBLM_R_X53Y98_SLICE_X81Y98_AO6),
.O5(CLBLL_L_X54Y99_SLICE_X82Y99_CO5),
.O6(CLBLL_L_X54Y99_SLICE_X82Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffaffffdccceece)
  ) CLBLL_L_X54Y99_SLICE_X82Y99_BLUT (
.I0(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I1(CLBLM_R_X53Y99_SLICE_X81Y99_CO6),
.I2(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.I3(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.I4(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.I5(1'b1),
.O5(CLBLL_L_X54Y99_SLICE_X82Y99_BO5),
.O6(CLBLL_L_X54Y99_SLICE_X82Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbfffbf40024002)
  ) CLBLL_L_X54Y99_SLICE_X82Y99_ALUT (
.I0(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I1(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.I2(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.I3(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y99_SLICE_X82Y99_AO5),
.O6(CLBLL_L_X54Y99_SLICE_X82Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLL_L_X54Y99_SLICE_X83Y99_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X0Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_L_X54Y99_SLICE_X83Y99_AQ),
.Q(CLBLL_L_X54Y99_SLICE_X83Y99_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLL_L_X54Y99_SLICE_X83Y99_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X0Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_L_X54Y99_SLICE_X83Y99_AO6),
.Q(CLBLL_L_X54Y99_SLICE_X83Y99_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000030007c)
  ) CLBLL_L_X54Y99_SLICE_X83Y99_DLUT (
.I0(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.I1(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.I2(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.I3(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I4(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I5(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.O5(CLBLL_L_X54Y99_SLICE_X83Y99_DO5),
.O6(CLBLL_L_X54Y99_SLICE_X83Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000550100000000)
  ) CLBLL_L_X54Y99_SLICE_X83Y99_CLUT (
.I0(CLBLL_L_X54Y98_SLICE_X83Y98_CO5),
.I1(CLBLM_R_X49Y108_SLICE_X75Y108_DQ),
.I2(CLBLM_R_X49Y107_SLICE_X75Y107_DQ),
.I3(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.I4(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.I5(CLBLL_L_X54Y99_SLICE_X83Y99_BO6),
.O5(CLBLL_L_X54Y99_SLICE_X83Y99_CO5),
.O6(CLBLL_L_X54Y99_SLICE_X83Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0c0c0cc0c0c0c0)
  ) CLBLL_L_X54Y99_SLICE_X83Y99_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I2(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y99_SLICE_X83Y99_BO5),
.O6(CLBLL_L_X54Y99_SLICE_X83Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffbfafafa)
  ) CLBLL_L_X54Y99_SLICE_X83Y99_ALUT (
.I0(CLBLL_L_X54Y99_SLICE_X83Y99_DO6),
.I1(CLBLM_R_X53Y99_SLICE_X80Y99_AO5),
.I2(CLBLL_L_X52Y99_SLICE_X79Y99_AO6),
.I3(CLBLL_L_X54Y99_SLICE_X83Y99_BO6),
.I4(CLBLM_R_X49Y107_SLICE_X75Y107_DQ),
.I5(CLBLL_L_X54Y100_SLICE_X83Y100_AO5),
.O5(CLBLL_L_X54Y99_SLICE_X83Y99_AO5),
.O6(CLBLL_L_X54Y99_SLICE_X83Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLL_L_X54Y100_SLICE_X82Y100_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_L_X54Y100_SLICE_X82Y100_BO6),
.Q(CLBLL_L_X54Y100_SLICE_X82Y100_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfccfffdcdcfcfc)
  ) CLBLL_L_X54Y100_SLICE_X82Y100_DLUT (
.I0(CLBLL_L_X54Y99_SLICE_X82Y99_BO6),
.I1(CLBLL_L_X54Y100_SLICE_X83Y100_CO6),
.I2(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I3(CLBLL_L_X54Y100_SLICE_X82Y100_AO5),
.I4(CLBLL_L_X54Y99_SLICE_X82Y99_AO6),
.I5(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.O5(CLBLL_L_X54Y100_SLICE_X82Y100_DO5),
.O6(CLBLL_L_X54Y100_SLICE_X82Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff05c5ffff0000)
  ) CLBLL_L_X54Y100_SLICE_X82Y100_CLUT (
.I0(CLBLL_L_X54Y100_SLICE_X82Y100_AO6),
.I1(CLBLM_R_X49Y107_SLICE_X75Y107_DQ),
.I2(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I3(CLBLM_R_X53Y99_SLICE_X80Y99_AO5),
.I4(CLBLL_L_X54Y99_SLICE_X82Y99_DO6),
.I5(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.O5(CLBLL_L_X54Y100_SLICE_X82Y100_CO5),
.O6(CLBLL_L_X54Y100_SLICE_X82Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffefffe)
  ) CLBLL_L_X54Y100_SLICE_X82Y100_BLUT (
.I0(CLBLL_L_X54Y100_SLICE_X82Y100_DO6),
.I1(CLBLL_L_X54Y100_SLICE_X83Y100_BO6),
.I2(CLBLL_L_X54Y100_SLICE_X83Y100_AO6),
.I3(CLBLM_L_X56Y99_SLICE_X84Y99_CO6),
.I4(1'b1),
.I5(CLBLL_L_X54Y100_SLICE_X82Y100_CO6),
.O5(CLBLL_L_X54Y100_SLICE_X82Y100_BO5),
.O6(CLBLL_L_X54Y100_SLICE_X82Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffefffefffbfffbf)
  ) CLBLL_L_X54Y100_SLICE_X82Y100_ALUT (
.I0(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.I1(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.I2(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.I3(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y100_SLICE_X82Y100_AO5),
.O6(CLBLL_L_X54Y100_SLICE_X82Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y100_SLICE_X83Y100_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y100_SLICE_X83Y100_DO5),
.O6(CLBLL_L_X54Y100_SLICE_X83Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f0f3f0f0f3f3)
  ) CLBLL_L_X54Y100_SLICE_X83Y100_CLUT (
.I0(CLBLL_L_X54Y99_SLICE_X82Y99_AO6),
.I1(CLBLM_R_X53Y99_SLICE_X80Y99_AO5),
.I2(CLBLL_L_X54Y99_SLICE_X83Y99_CO6),
.I3(CLBLM_R_X49Y107_SLICE_X75Y107_DQ),
.I4(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I5(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.O5(CLBLL_L_X54Y100_SLICE_X83Y100_CO5),
.O6(CLBLL_L_X54Y100_SLICE_X83Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000103000000)
  ) CLBLL_L_X54Y100_SLICE_X83Y100_BLUT (
.I0(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I1(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.I2(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I3(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.I4(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.I5(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.O5(CLBLL_L_X54Y100_SLICE_X83Y100_BO5),
.O6(CLBLL_L_X54Y100_SLICE_X83Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2088000022200000)
  ) CLBLL_L_X54Y100_SLICE_X83Y100_ALUT (
.I0(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I1(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.I2(CLBLM_R_X49Y107_SLICE_X75Y107_DQ),
.I3(CLBLM_R_X49Y108_SLICE_X75Y108_DQ),
.I4(CLBLM_L_X56Y97_SLICE_X84Y97_CO5),
.I5(1'b1),
.O5(CLBLL_L_X54Y100_SLICE_X83Y100_AO5),
.O6(CLBLL_L_X54Y100_SLICE_X83Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLL_L_X54Y101_SLICE_X82Y101_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X56Y98_SLICE_X84Y98_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_L_X54Y101_SLICE_X82Y101_AO6),
.Q(CLBLL_L_X54Y101_SLICE_X82Y101_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLL_L_X54Y101_SLICE_X82Y101_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X56Y98_SLICE_X84Y98_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_L_X54Y101_SLICE_X82Y101_AO5),
.Q(CLBLL_L_X54Y101_SLICE_X82Y101_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y101_SLICE_X82Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y101_SLICE_X82Y101_DO5),
.O6(CLBLL_L_X54Y101_SLICE_X82Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y101_SLICE_X82Y101_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y101_SLICE_X82Y101_CO5),
.O6(CLBLL_L_X54Y101_SLICE_X82Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y101_SLICE_X82Y101_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y101_SLICE_X82Y101_BO5),
.O6(CLBLL_L_X54Y101_SLICE_X82Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0404040402020202)
  ) CLBLL_L_X54Y101_SLICE_X82Y101_ALUT (
.I0(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I1(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.I2(CLBLM_R_X49Y107_SLICE_X75Y107_DQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y101_SLICE_X82Y101_AO5),
.O6(CLBLL_L_X54Y101_SLICE_X82Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y101_SLICE_X83Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y101_SLICE_X83Y101_DO5),
.O6(CLBLL_L_X54Y101_SLICE_X83Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0030003000000000)
  ) CLBLL_L_X54Y101_SLICE_X83Y101_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X53Y100_SLICE_X80Y100_A5Q),
.I2(CLBLM_R_X53Y100_SLICE_X80Y100_AQ),
.I3(CLBLM_R_X53Y101_SLICE_X80Y101_BQ),
.I4(1'b1),
.I5(CLBLM_R_X53Y101_SLICE_X81Y101_AQ),
.O5(CLBLL_L_X54Y101_SLICE_X83Y101_CO5),
.O6(CLBLL_L_X54Y101_SLICE_X83Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff7fffffff)
  ) CLBLL_L_X54Y101_SLICE_X83Y101_BLUT (
.I0(CLBLM_R_X53Y100_SLICE_X80Y100_AQ),
.I1(CLBLM_R_X53Y101_SLICE_X81Y101_AQ),
.I2(CLBLM_R_X53Y100_SLICE_X81Y100_AQ),
.I3(CLBLL_L_X54Y100_SLICE_X82Y100_BQ),
.I4(CLBLM_R_X53Y101_SLICE_X80Y101_BQ),
.I5(CLBLM_R_X53Y100_SLICE_X80Y100_A5Q),
.O5(CLBLL_L_X54Y101_SLICE_X83Y101_BO5),
.O6(CLBLL_L_X54Y101_SLICE_X83Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000008000000)
  ) CLBLL_L_X54Y101_SLICE_X83Y101_ALUT (
.I0(CLBLM_R_X53Y100_SLICE_X80Y100_AQ),
.I1(CLBLM_R_X53Y101_SLICE_X81Y101_AQ),
.I2(CLBLM_R_X53Y101_SLICE_X80Y101_BQ),
.I3(CLBLL_L_X54Y100_SLICE_X82Y100_BQ),
.I4(CLBLM_R_X53Y100_SLICE_X81Y100_AQ),
.I5(CLBLM_R_X53Y100_SLICE_X80Y100_A5Q),
.O5(CLBLL_L_X54Y101_SLICE_X83Y101_AO5),
.O6(CLBLL_L_X54Y101_SLICE_X83Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y102_SLICE_X82Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y102_SLICE_X82Y102_DO5),
.O6(CLBLL_L_X54Y102_SLICE_X82Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000040)
  ) CLBLL_L_X54Y102_SLICE_X82Y102_CLUT (
.I0(CLBLM_R_X49Y107_SLICE_X75Y107_DQ),
.I1(CLBLM_L_X56Y97_SLICE_X84Y97_CO5),
.I2(CLBLM_R_X49Y104_SLICE_X75Y104_DQ),
.I3(CLBLM_R_X49Y108_SLICE_X75Y108_DQ),
.I4(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I5(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.O5(CLBLL_L_X54Y102_SLICE_X82Y102_CO5),
.O6(CLBLL_L_X54Y102_SLICE_X82Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000100000000)
  ) CLBLL_L_X54Y102_SLICE_X82Y102_BLUT (
.I0(CLBLM_R_X49Y106_SLICE_X75Y106_DQ),
.I1(CLBLM_R_X49Y106_SLICE_X75Y106_CQ),
.I2(CLBLM_R_X49Y107_SLICE_X75Y107_CQ),
.I3(CLBLM_R_X49Y104_SLICE_X75Y104_CQ),
.I4(CLBLM_R_X49Y104_SLICE_X75Y104_BQ),
.I5(CLBLL_L_X54Y102_SLICE_X82Y102_CO6),
.O5(CLBLL_L_X54Y102_SLICE_X82Y102_BO5),
.O6(CLBLL_L_X54Y102_SLICE_X82Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3ffffffffffffefe)
  ) CLBLL_L_X54Y102_SLICE_X82Y102_ALUT (
.I0(CLBLM_R_X49Y106_SLICE_X75Y106_DQ),
.I1(CLBLM_R_X49Y104_SLICE_X75Y104_BQ),
.I2(CLBLM_R_X49Y107_SLICE_X75Y107_CQ),
.I3(CLBLM_R_X49Y106_SLICE_X75Y106_CQ),
.I4(CLBLM_R_X49Y104_SLICE_X75Y104_CQ),
.I5(1'b1),
.O5(CLBLL_L_X54Y102_SLICE_X82Y102_AO5),
.O6(CLBLL_L_X54Y102_SLICE_X82Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y102_SLICE_X83Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y102_SLICE_X83Y102_DO5),
.O6(CLBLL_L_X54Y102_SLICE_X83Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y102_SLICE_X83Y102_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y102_SLICE_X83Y102_CO5),
.O6(CLBLL_L_X54Y102_SLICE_X83Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y102_SLICE_X83Y102_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y102_SLICE_X83Y102_BO5),
.O6(CLBLL_L_X54Y102_SLICE_X83Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y102_SLICE_X83Y102_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y102_SLICE_X83Y102_AO5),
.O6(CLBLL_L_X54Y102_SLICE_X83Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLL_L_X54Y103_SLICE_X82Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(CLBLM_R_X15Y122_SLICE_X20Y122_AO6),
.D(CLBLL_L_X54Y103_SLICE_X82Y103_AO6),
.Q(CLBLL_L_X54Y103_SLICE_X82Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y103_SLICE_X82Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y103_SLICE_X82Y103_DO5),
.O6(CLBLL_L_X54Y103_SLICE_X82Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y103_SLICE_X82Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y103_SLICE_X82Y103_CO5),
.O6(CLBLL_L_X54Y103_SLICE_X82Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y103_SLICE_X82Y103_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y103_SLICE_X82Y103_BO5),
.O6(CLBLL_L_X54Y103_SLICE_X82Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff007f00ff00ff)
  ) CLBLL_L_X54Y103_SLICE_X82Y103_ALUT (
.I0(CLBLM_R_X49Y104_SLICE_X75Y104_AQ),
.I1(CLBLM_R_X49Y104_SLICE_X74Y104_AQ),
.I2(CLBLM_R_X49Y106_SLICE_X75Y106_DQ),
.I3(CLBLM_L_X56Y104_SLICE_X84Y104_AQ),
.I4(CLBLL_L_X54Y102_SLICE_X82Y102_AO6),
.I5(CLBLL_L_X54Y102_SLICE_X82Y102_CO6),
.O5(CLBLL_L_X54Y103_SLICE_X82Y103_AO5),
.O6(CLBLL_L_X54Y103_SLICE_X82Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y103_SLICE_X83Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y103_SLICE_X83Y103_DO5),
.O6(CLBLL_L_X54Y103_SLICE_X83Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y103_SLICE_X83Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y103_SLICE_X83Y103_CO5),
.O6(CLBLL_L_X54Y103_SLICE_X83Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y103_SLICE_X83Y103_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y103_SLICE_X83Y103_BO5),
.O6(CLBLL_L_X54Y103_SLICE_X83Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y103_SLICE_X83Y103_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y103_SLICE_X83Y103_AO5),
.O6(CLBLL_L_X54Y103_SLICE_X83Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y104_SLICE_X82Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y104_SLICE_X82Y104_DO5),
.O6(CLBLL_L_X54Y104_SLICE_X82Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y104_SLICE_X82Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y104_SLICE_X82Y104_CO5),
.O6(CLBLL_L_X54Y104_SLICE_X82Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hec808080a0000000)
  ) CLBLL_L_X54Y104_SLICE_X82Y104_BLUT (
.I0(CLBLM_L_X56Y101_SLICE_X85Y101_BQ),
.I1(CLBLM_L_X56Y101_SLICE_X85Y101_CQ),
.I2(CLBLL_R_X57Y100_SLICE_X86Y100_CQ),
.I3(CLBLL_R_X57Y100_SLICE_X87Y100_BQ),
.I4(CLBLL_R_X57Y100_SLICE_X86Y100_DQ),
.I5(CLBLL_R_X57Y101_SLICE_X87Y101_AQ),
.O5(CLBLL_L_X54Y104_SLICE_X82Y104_BO5),
.O6(CLBLL_L_X54Y104_SLICE_X82Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he888a000c0000000)
  ) CLBLL_L_X54Y104_SLICE_X82Y104_ALUT (
.I0(CLBLM_L_X56Y101_SLICE_X85Y101_BQ),
.I1(CLBLM_L_X56Y101_SLICE_X85Y101_CQ),
.I2(CLBLL_R_X57Y100_SLICE_X86Y100_CQ),
.I3(CLBLL_R_X57Y101_SLICE_X87Y101_AQ),
.I4(CLBLL_R_X57Y100_SLICE_X87Y100_AQ),
.I5(CLBLL_R_X57Y100_SLICE_X86Y100_DQ),
.O5(CLBLL_L_X54Y104_SLICE_X82Y104_AO5),
.O6(CLBLL_L_X54Y104_SLICE_X82Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y104_SLICE_X83Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y104_SLICE_X83Y104_DO5),
.O6(CLBLL_L_X54Y104_SLICE_X83Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y104_SLICE_X83Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y104_SLICE_X83Y104_CO5),
.O6(CLBLL_L_X54Y104_SLICE_X83Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y104_SLICE_X83Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y104_SLICE_X83Y104_BO5),
.O6(CLBLL_L_X54Y104_SLICE_X83Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y104_SLICE_X83Y104_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y104_SLICE_X83Y104_AO5),
.O6(CLBLL_L_X54Y104_SLICE_X83Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_L_X54Y105_SLICE_X82Y105_CARRY4 (
.CI(1'b0),
.CO({CLBLL_L_X54Y105_SLICE_X82Y105_D_CY, CLBLL_L_X54Y105_SLICE_X82Y105_C_CY, CLBLL_L_X54Y105_SLICE_X82Y105_B_CY, CLBLL_L_X54Y105_SLICE_X82Y105_A_CY}),
.CYINIT(1'b0),
.DI({CLBLL_L_X54Y105_SLICE_X82Y105_DO5, CLBLM_R_X53Y104_SLICE_X81Y104_B_XOR, CLBLM_R_X53Y104_SLICE_X81Y104_A_XOR, CLBLM_R_X53Y103_SLICE_X81Y103_D_XOR}),
.O({CLBLL_L_X54Y105_SLICE_X82Y105_D_XOR, CLBLL_L_X54Y105_SLICE_X82Y105_C_XOR, CLBLL_L_X54Y105_SLICE_X82Y105_B_XOR, CLBLL_L_X54Y105_SLICE_X82Y105_A_XOR}),
.S({CLBLL_L_X54Y105_SLICE_X82Y105_DO6, CLBLL_L_X54Y105_SLICE_X82Y105_CO6, CLBLL_L_X54Y105_SLICE_X82Y105_BO6, CLBLL_L_X54Y105_SLICE_X82Y105_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9666966666666666)
  ) CLBLL_L_X54Y105_SLICE_X82Y105_DLUT (
.I0(CLBLM_R_X53Y104_SLICE_X81Y104_C_XOR),
.I1(CLBLM_R_X53Y106_SLICE_X81Y106_D_XOR),
.I2(CLBLL_R_X57Y100_SLICE_X86Y100_AQ),
.I3(CLBLL_R_X57Y101_SLICE_X87Y101_DQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y105_SLICE_X82Y105_DO5),
.O6(CLBLL_L_X54Y105_SLICE_X82Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5a5a5a5a5a)
  ) CLBLL_L_X54Y105_SLICE_X82Y105_CLUT (
.I0(CLBLM_R_X53Y104_SLICE_X81Y104_B_XOR),
.I1(1'b1),
.I2(CLBLM_R_X53Y106_SLICE_X81Y106_C_XOR),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y105_SLICE_X82Y105_CO5),
.O6(CLBLL_L_X54Y105_SLICE_X82Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa55aa55aa55aa)
  ) CLBLL_L_X54Y105_SLICE_X82Y105_BLUT (
.I0(CLBLM_R_X53Y106_SLICE_X81Y106_B_XOR),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X53Y104_SLICE_X81Y104_A_XOR),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y105_SLICE_X82Y105_BO5),
.O6(CLBLL_L_X54Y105_SLICE_X82Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffffffff0000)
  ) CLBLL_L_X54Y105_SLICE_X82Y105_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X53Y103_SLICE_X81Y103_D_XOR),
.I5(CLBLM_R_X53Y106_SLICE_X81Y106_A_XOR),
.O5(CLBLL_L_X54Y105_SLICE_X82Y105_AO5),
.O6(CLBLL_L_X54Y105_SLICE_X82Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y105_SLICE_X83Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y105_SLICE_X83Y105_DO5),
.O6(CLBLL_L_X54Y105_SLICE_X83Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y105_SLICE_X83Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y105_SLICE_X83Y105_CO5),
.O6(CLBLL_L_X54Y105_SLICE_X83Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y105_SLICE_X83Y105_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y105_SLICE_X83Y105_BO5),
.O6(CLBLL_L_X54Y105_SLICE_X83Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y105_SLICE_X83Y105_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y105_SLICE_X83Y105_AO5),
.O6(CLBLL_L_X54Y105_SLICE_X83Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_L_X54Y106_SLICE_X82Y106_CARRY4 (
.CI(CLBLL_L_X54Y105_SLICE_X82Y105_COUT),
.CO({CLBLL_L_X54Y106_SLICE_X82Y106_D_CY, CLBLL_L_X54Y106_SLICE_X82Y106_C_CY, CLBLL_L_X54Y106_SLICE_X82Y106_B_CY, CLBLL_L_X54Y106_SLICE_X82Y106_A_CY}),
.CYINIT(1'b0),
.DI({CLBLL_L_X54Y106_SLICE_X83Y106_BO6, CLBLM_R_X53Y105_SLICE_X80Y105_AO6, CLBLM_R_X53Y106_SLICE_X80Y106_BO6, CLBLL_L_X54Y106_SLICE_X83Y106_CO6}),
.O({CLBLL_L_X54Y106_SLICE_X82Y106_D_XOR, CLBLL_L_X54Y106_SLICE_X82Y106_C_XOR, CLBLL_L_X54Y106_SLICE_X82Y106_B_XOR, CLBLL_L_X54Y106_SLICE_X82Y106_A_XOR}),
.S({CLBLL_L_X54Y106_SLICE_X82Y106_DO6, CLBLL_L_X54Y106_SLICE_X82Y106_CO6, CLBLL_L_X54Y106_SLICE_X82Y106_BO6, CLBLL_L_X54Y106_SLICE_X82Y106_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h963c69c3963c69c3)
  ) CLBLL_L_X54Y106_SLICE_X82Y106_DLUT (
.I0(CLBLL_R_X57Y101_SLICE_X87Y101_AQ),
.I1(CLBLL_L_X54Y106_SLICE_X83Y106_AO5),
.I2(CLBLL_L_X54Y106_SLICE_X83Y106_BO6),
.I3(CLBLL_R_X57Y101_SLICE_X87Y101_DQ),
.I4(CLBLM_R_X53Y107_SLICE_X80Y107_BO5),
.I5(1'b1),
.O5(CLBLL_L_X54Y106_SLICE_X82Y106_DO5),
.O6(CLBLL_L_X54Y106_SLICE_X82Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9696666669699999)
  ) CLBLL_L_X54Y106_SLICE_X82Y106_CLUT (
.I0(CLBLM_R_X53Y105_SLICE_X80Y105_AO6),
.I1(CLBLL_L_X54Y106_SLICE_X83Y106_AO6),
.I2(CLBLL_R_X57Y101_SLICE_X87Y101_DQ),
.I3(1'b1),
.I4(CLBLL_R_X57Y100_SLICE_X87Y100_AQ),
.I5(CLBLM_R_X53Y106_SLICE_X80Y106_AO6),
.O5(CLBLL_L_X54Y106_SLICE_X82Y106_CO5),
.O6(CLBLL_L_X54Y106_SLICE_X82Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f780f7878f078f0)
  ) CLBLL_L_X54Y106_SLICE_X82Y106_BLUT (
.I0(CLBLL_R_X57Y99_SLICE_X86Y99_BQ),
.I1(CLBLL_R_X57Y100_SLICE_X86Y100_AQ),
.I2(CLBLM_R_X53Y106_SLICE_X80Y106_BO6),
.I3(CLBLM_R_X53Y104_SLICE_X81Y104_D_XOR),
.I4(1'b1),
.I5(CLBLM_R_X53Y107_SLICE_X81Y107_A_XOR),
.O5(CLBLL_L_X54Y106_SLICE_X82Y106_BO5),
.O6(CLBLL_L_X54Y106_SLICE_X82Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h965a3cf0965a3cf0)
  ) CLBLL_L_X54Y106_SLICE_X82Y106_ALUT (
.I0(CLBLM_R_X53Y106_SLICE_X81Y106_D_XOR),
.I1(CLBLL_R_X57Y101_SLICE_X87Y101_DQ),
.I2(CLBLL_L_X54Y106_SLICE_X83Y106_CO6),
.I3(CLBLL_R_X57Y100_SLICE_X86Y100_BQ),
.I4(CLBLM_R_X53Y104_SLICE_X81Y104_C_XOR),
.I5(1'b1),
.O5(CLBLL_L_X54Y106_SLICE_X82Y106_AO5),
.O6(CLBLL_L_X54Y106_SLICE_X82Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0fc00f0c0fc00f0)
  ) CLBLL_L_X54Y106_SLICE_X83Y106_DLUT (
.I0(1'b1),
.I1(CLBLL_R_X57Y101_SLICE_X87Y101_DQ),
.I2(CLBLM_R_X53Y107_SLICE_X80Y107_BO5),
.I3(CLBLL_L_X54Y106_SLICE_X83Y106_AO5),
.I4(CLBLL_R_X57Y101_SLICE_X87Y101_AQ),
.I5(1'b1),
.O5(CLBLL_L_X54Y106_SLICE_X83Y106_DO5),
.O6(CLBLL_L_X54Y106_SLICE_X83Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h939393936c6c6c6c)
  ) CLBLL_L_X54Y106_SLICE_X83Y106_CLUT (
.I0(CLBLL_R_X57Y100_SLICE_X86Y100_AQ),
.I1(CLBLM_R_X53Y107_SLICE_X81Y107_A_XOR),
.I2(CLBLL_R_X57Y99_SLICE_X86Y99_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X53Y104_SLICE_X81Y104_D_XOR),
.O5(CLBLL_L_X54Y106_SLICE_X83Y106_CO5),
.O6(CLBLL_L_X54Y106_SLICE_X83Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb332200bb332200)
  ) CLBLL_L_X54Y106_SLICE_X83Y106_BLUT (
.I0(CLBLL_R_X57Y101_SLICE_X87Y101_DQ),
.I1(CLBLM_R_X53Y106_SLICE_X80Y106_AO6),
.I2(1'b1),
.I3(CLBLL_R_X57Y100_SLICE_X87Y100_AQ),
.I4(CLBLL_L_X54Y106_SLICE_X83Y106_AO6),
.I5(1'b1),
.O5(CLBLL_L_X54Y106_SLICE_X83Y106_BO5),
.O6(CLBLL_L_X54Y106_SLICE_X83Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc33c0ff0033f0fff)
  ) CLBLL_L_X54Y106_SLICE_X83Y106_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X56Y101_SLICE_X85Y101_AQ),
.I2(CLBLM_R_X53Y107_SLICE_X81Y107_C_XOR),
.I3(CLBLM_R_X53Y105_SLICE_X81Y105_B_XOR),
.I4(CLBLL_R_X57Y99_SLICE_X86Y99_BQ),
.I5(1'b1),
.O5(CLBLL_L_X54Y106_SLICE_X83Y106_AO5),
.O6(CLBLL_L_X54Y106_SLICE_X83Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_L_X54Y107_SLICE_X82Y107_CARRY4 (
.CI(CLBLL_L_X54Y106_SLICE_X82Y106_COUT),
.CO({CLBLL_L_X54Y107_SLICE_X82Y107_D_CY, CLBLL_L_X54Y107_SLICE_X82Y107_C_CY, CLBLL_L_X54Y107_SLICE_X82Y107_B_CY, CLBLL_L_X54Y107_SLICE_X82Y107_A_CY}),
.CYINIT(1'b0),
.DI({CLBLL_L_X54Y107_SLICE_X83Y107_BO6, CLBLL_L_X54Y107_SLICE_X83Y107_CO6, CLBLL_L_X54Y107_SLICE_X83Y107_DO6, CLBLL_L_X54Y106_SLICE_X83Y106_DO6}),
.O({CLBLL_L_X54Y107_SLICE_X82Y107_D_XOR, CLBLL_L_X54Y107_SLICE_X82Y107_C_XOR, CLBLL_L_X54Y107_SLICE_X82Y107_B_XOR, CLBLL_L_X54Y107_SLICE_X82Y107_A_XOR}),
.S({CLBLL_L_X54Y107_SLICE_X82Y107_DO6, CLBLL_L_X54Y107_SLICE_X82Y107_CO6, CLBLL_L_X54Y107_SLICE_X82Y107_BO6, CLBLL_L_X54Y107_SLICE_X82Y107_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb236fcf0246cc000)
  ) CLBLL_L_X54Y107_SLICE_X82Y107_DLUT (
.I0(CLBLL_R_X57Y101_SLICE_X87Y101_DQ),
.I1(CLBLL_R_X57Y99_SLICE_X86Y99_BQ),
.I2(CLBLL_L_X54Y107_SLICE_X83Y107_AO6),
.I3(CLBLL_R_X57Y100_SLICE_X87Y100_BQ),
.I4(CLBLL_R_X57Y99_SLICE_X86Y99_AQ),
.I5(CLBLM_R_X53Y108_SLICE_X81Y108_C_CY),
.O5(CLBLL_L_X54Y107_SLICE_X82Y107_DO5),
.O6(CLBLL_L_X54Y107_SLICE_X82Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999999996666666)
  ) CLBLL_L_X54Y107_SLICE_X82Y107_CLUT (
.I0(CLBLL_L_X52Y106_SLICE_X78Y106_AO6),
.I1(CLBLL_L_X54Y107_SLICE_X83Y107_CO6),
.I2(CLBLM_R_X53Y108_SLICE_X81Y108_B_XOR),
.I3(CLBLL_R_X57Y99_SLICE_X86Y99_BQ),
.I4(CLBLM_L_X56Y101_SLICE_X85Y101_BQ),
.I5(CLBLL_L_X54Y108_SLICE_X83Y108_AO6),
.O5(CLBLL_L_X54Y107_SLICE_X82Y107_CO5),
.O6(CLBLL_L_X54Y107_SLICE_X82Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996996699669966)
  ) CLBLL_L_X54Y107_SLICE_X82Y107_BLUT (
.I0(CLBLL_L_X54Y108_SLICE_X83Y108_AO5),
.I1(CLBLL_L_X54Y107_SLICE_X83Y107_DO6),
.I2(CLBLL_R_X57Y101_SLICE_X87Y101_AQ),
.I3(CLBLL_L_X52Y107_SLICE_X78Y107_BO6),
.I4(CLBLL_R_X57Y99_SLICE_X86Y99_BQ),
.I5(CLBLM_R_X53Y108_SLICE_X81Y108_A_XOR),
.O5(CLBLL_L_X54Y107_SLICE_X82Y107_BO5),
.O6(CLBLL_L_X54Y107_SLICE_X82Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h9966669955aaaa55)
  ) CLBLL_L_X54Y107_SLICE_X82Y107_ALUT (
.I0(CLBLL_L_X54Y106_SLICE_X83Y106_DO6),
.I1(CLBLM_L_X56Y101_SLICE_X85Y101_BQ),
.I2(1'b1),
.I3(CLBLL_L_X54Y107_SLICE_X83Y107_AO5),
.I4(CLBLM_R_X53Y107_SLICE_X80Y107_BO6),
.I5(CLBLL_R_X57Y101_SLICE_X87Y101_DQ),
.O5(CLBLL_L_X54Y107_SLICE_X82Y107_AO5),
.O6(CLBLL_L_X54Y107_SLICE_X82Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h20b380eca0ff00a0)
  ) CLBLL_L_X54Y107_SLICE_X83Y107_DLUT (
.I0(CLBLL_R_X57Y101_SLICE_X87Y101_DQ),
.I1(CLBLL_R_X57Y101_SLICE_X87Y101_AQ),
.I2(CLBLM_L_X56Y101_SLICE_X85Y101_BQ),
.I3(CLBLM_R_X53Y107_SLICE_X80Y107_BO6),
.I4(CLBLM_R_X53Y108_SLICE_X81Y108_A_XOR),
.I5(CLBLL_R_X57Y99_SLICE_X86Y99_BQ),
.O5(CLBLL_L_X54Y107_SLICE_X83Y107_DO5),
.O6(CLBLL_L_X54Y107_SLICE_X83Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdeaa5aaa48000000)
  ) CLBLL_L_X54Y107_SLICE_X83Y107_CLUT (
.I0(CLBLM_R_X53Y108_SLICE_X81Y108_B_XOR),
.I1(CLBLL_R_X57Y101_SLICE_X87Y101_AQ),
.I2(CLBLM_L_X56Y101_SLICE_X85Y101_BQ),
.I3(CLBLL_R_X57Y99_SLICE_X86Y99_BQ),
.I4(CLBLM_R_X53Y108_SLICE_X81Y108_A_XOR),
.I5(CLBLL_L_X52Y107_SLICE_X78Y107_BO6),
.O5(CLBLL_L_X54Y107_SLICE_X83Y107_CO5),
.O6(CLBLL_L_X54Y107_SLICE_X83Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb2c030c0e8c0c0c0)
  ) CLBLL_L_X54Y107_SLICE_X83Y107_BLUT (
.I0(CLBLM_R_X53Y108_SLICE_X81Y108_B_XOR),
.I1(CLBLM_R_X53Y108_SLICE_X81Y108_C_CY),
.I2(CLBLL_L_X52Y106_SLICE_X78Y106_AO6),
.I3(CLBLL_R_X57Y99_SLICE_X86Y99_BQ),
.I4(CLBLM_L_X56Y101_SLICE_X85Y101_BQ),
.I5(CLBLL_R_X57Y100_SLICE_X87Y100_BQ),
.O5(CLBLL_L_X54Y107_SLICE_X83Y107_BO5),
.O6(CLBLL_L_X54Y107_SLICE_X83Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf00000006a6a6a6a)
  ) CLBLL_L_X54Y107_SLICE_X83Y107_ALUT (
.I0(CLBLM_R_X53Y108_SLICE_X81Y108_A_XOR),
.I1(CLBLL_R_X57Y101_SLICE_X87Y101_AQ),
.I2(CLBLL_R_X57Y99_SLICE_X86Y99_BQ),
.I3(CLBLM_L_X56Y101_SLICE_X85Y101_BQ),
.I4(CLBLM_R_X53Y108_SLICE_X81Y108_B_XOR),
.I5(1'b1),
.O5(CLBLL_L_X54Y107_SLICE_X83Y107_AO5),
.O6(CLBLL_L_X54Y107_SLICE_X83Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_L_X54Y108_SLICE_X82Y108_CARRY4 (
.CI(CLBLL_L_X54Y107_SLICE_X82Y107_COUT),
.CO({CLBLL_L_X54Y108_SLICE_X82Y108_D_CY, CLBLL_L_X54Y108_SLICE_X82Y108_C_CY, CLBLL_L_X54Y108_SLICE_X82Y108_B_CY, CLBLL_L_X54Y108_SLICE_X82Y108_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLL_L_X54Y108_SLICE_X82Y108_D_XOR, CLBLL_L_X54Y108_SLICE_X82Y108_C_XOR, CLBLL_L_X54Y108_SLICE_X82Y108_B_XOR, CLBLL_L_X54Y108_SLICE_X82Y108_A_XOR}),
.S({CLBLL_L_X54Y108_SLICE_X82Y108_DO6, CLBLL_L_X54Y108_SLICE_X82Y108_CO6, CLBLL_L_X54Y108_SLICE_X82Y108_BO6, CLBLL_L_X54Y108_SLICE_X82Y108_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y108_SLICE_X82Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y108_SLICE_X82Y108_DO5),
.O6(CLBLL_L_X54Y108_SLICE_X82Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y108_SLICE_X82Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y108_SLICE_X82Y108_CO5),
.O6(CLBLL_L_X54Y108_SLICE_X82Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y108_SLICE_X82Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y108_SLICE_X82Y108_BO5),
.O6(CLBLL_L_X54Y108_SLICE_X82Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000000000000000)
  ) CLBLL_L_X54Y108_SLICE_X82Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_R_X57Y99_SLICE_X86Y99_AQ),
.I3(CLBLM_R_X53Y108_SLICE_X81Y108_C_CY),
.I4(CLBLL_R_X57Y99_SLICE_X86Y99_BQ),
.I5(CLBLL_R_X57Y100_SLICE_X87Y100_BQ),
.O5(CLBLL_L_X54Y108_SLICE_X82Y108_AO5),
.O6(CLBLL_L_X54Y108_SLICE_X82Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y108_SLICE_X83Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y108_SLICE_X83Y108_DO5),
.O6(CLBLL_L_X54Y108_SLICE_X83Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y108_SLICE_X83Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y108_SLICE_X83Y108_CO5),
.O6(CLBLL_L_X54Y108_SLICE_X83Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y108_SLICE_X83Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y108_SLICE_X83Y108_BO5),
.O6(CLBLL_L_X54Y108_SLICE_X83Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6666cccc5af05af0)
  ) CLBLL_L_X54Y108_SLICE_X83Y108_ALUT (
.I0(CLBLL_R_X57Y99_SLICE_X86Y99_BQ),
.I1(CLBLM_R_X53Y108_SLICE_X81Y108_C_CY),
.I2(CLBLM_R_X53Y108_SLICE_X81Y108_B_XOR),
.I3(CLBLM_L_X56Y101_SLICE_X85Y101_BQ),
.I4(CLBLL_R_X57Y100_SLICE_X87Y100_BQ),
.I5(1'b1),
.O5(CLBLL_L_X54Y108_SLICE_X83Y108_AO5),
.O6(CLBLL_L_X54Y108_SLICE_X83Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLL_L_X54Y109_SLICE_X82Y109_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(CLBLM_R_X15Y122_SLICE_X20Y122_AO6),
.D(CLBLL_L_X54Y103_SLICE_X82Y103_AQ),
.Q(CLBLL_L_X54Y109_SLICE_X82Y109_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y109_SLICE_X82Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y109_SLICE_X82Y109_DO5),
.O6(CLBLL_L_X54Y109_SLICE_X82Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y109_SLICE_X82Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y109_SLICE_X82Y109_CO5),
.O6(CLBLL_L_X54Y109_SLICE_X82Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y109_SLICE_X82Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y109_SLICE_X82Y109_BO5),
.O6(CLBLL_L_X54Y109_SLICE_X82Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0f0f0f)
  ) CLBLL_L_X54Y109_SLICE_X82Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X54Y109_SLICE_X82Y109_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y109_SLICE_X82Y109_AO5),
.O6(CLBLL_L_X54Y109_SLICE_X82Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y109_SLICE_X83Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y109_SLICE_X83Y109_DO5),
.O6(CLBLL_L_X54Y109_SLICE_X83Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y109_SLICE_X83Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y109_SLICE_X83Y109_CO5),
.O6(CLBLL_L_X54Y109_SLICE_X83Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y109_SLICE_X83Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y109_SLICE_X83Y109_BO5),
.O6(CLBLL_L_X54Y109_SLICE_X83Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X54Y109_SLICE_X83Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X54Y109_SLICE_X83Y109_AO5),
.O6(CLBLL_L_X54Y109_SLICE_X83Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X57Y97_SLICE_X86Y97_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_R_X57Y97_SLICE_X86Y97_AO6),
.Q(CLBLL_R_X57Y97_SLICE_X86Y97_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y97_SLICE_X86Y97_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y97_SLICE_X86Y97_DO5),
.O6(CLBLL_R_X57Y97_SLICE_X86Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00000000)
  ) CLBLL_R_X57Y97_SLICE_X86Y97_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X56Y98_SLICE_X85Y98_CQ),
.I4(1'b1),
.I5(CLBLM_L_X56Y98_SLICE_X85Y98_BQ),
.O5(CLBLL_R_X57Y97_SLICE_X86Y97_CO5),
.O6(CLBLL_R_X57Y97_SLICE_X86Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00fd007500a80020)
  ) CLBLL_R_X57Y97_SLICE_X86Y97_BLUT (
.I0(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I1(CLBLL_R_X57Y97_SLICE_X86Y97_CO6),
.I2(CLBLL_R_X57Y97_SLICE_X86Y97_AQ),
.I3(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I4(CLBLL_R_X57Y97_SLICE_X87Y97_AQ),
.I5(CLBLM_L_X50Y105_SLICE_X76Y105_AQ),
.O5(CLBLL_R_X57Y97_SLICE_X86Y97_BO5),
.O6(CLBLL_R_X57Y97_SLICE_X86Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeaabaaaf0f0f0f0)
  ) CLBLL_R_X57Y97_SLICE_X86Y97_ALUT (
.I0(CLBLL_R_X57Y97_SLICE_X86Y97_BO6),
.I1(CLBLM_L_X60Y99_SLICE_X91Y99_DO6),
.I2(CLBLL_R_X57Y97_SLICE_X86Y97_AQ),
.I3(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I4(CLBLM_L_X50Y104_SLICE_X76Y104_AQ),
.I5(CLBLL_R_X57Y98_SLICE_X86Y98_AO6),
.O5(CLBLL_R_X57Y97_SLICE_X86Y97_AO5),
.O6(CLBLL_R_X57Y97_SLICE_X86Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X57Y97_SLICE_X87Y97_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_R_X57Y97_SLICE_X87Y97_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_R_X57Y97_SLICE_X86Y97_AQ),
.Q(CLBLL_R_X57Y97_SLICE_X87Y97_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y97_SLICE_X87Y97_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y97_SLICE_X87Y97_DO5),
.O6(CLBLL_R_X57Y97_SLICE_X87Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y97_SLICE_X87Y97_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y97_SLICE_X87Y97_CO5),
.O6(CLBLL_R_X57Y97_SLICE_X87Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y97_SLICE_X87Y97_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y97_SLICE_X87Y97_BO5),
.O6(CLBLL_R_X57Y97_SLICE_X87Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0088008800000000)
  ) CLBLL_R_X57Y97_SLICE_X87Y97_ALUT (
.I0(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.I1(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I2(1'b1),
.I3(CLBLM_L_X56Y98_SLICE_X85Y98_BQ),
.I4(1'b1),
.I5(CLBLM_L_X56Y98_SLICE_X85Y98_CQ),
.O5(CLBLL_R_X57Y97_SLICE_X87Y97_AO5),
.O6(CLBLL_R_X57Y97_SLICE_X87Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffbf200000000)
  ) CLBLL_R_X57Y98_SLICE_X86Y98_DLUT (
.I0(CLBLM_R_X53Y99_SLICE_X81Y99_AQ),
.I1(CLBLM_L_X56Y99_SLICE_X85Y99_A5Q),
.I2(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I3(CLBLL_L_X54Y99_SLICE_X83Y99_A5Q),
.I4(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I5(CLBLM_L_X62Y99_SLICE_X92Y99_AO6),
.O5(CLBLL_R_X57Y98_SLICE_X86Y98_DO5),
.O6(CLBLL_R_X57Y98_SLICE_X86Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff9f200000000)
  ) CLBLL_R_X57Y98_SLICE_X86Y98_CLUT (
.I0(CLBLM_R_X53Y99_SLICE_X81Y99_AQ),
.I1(CLBLM_L_X56Y99_SLICE_X85Y99_A5Q),
.I2(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I3(CLBLL_L_X54Y99_SLICE_X83Y99_A5Q),
.I4(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I5(CLBLM_L_X62Y99_SLICE_X92Y99_AO6),
.O5(CLBLL_R_X57Y98_SLICE_X86Y98_CO5),
.O6(CLBLL_R_X57Y98_SLICE_X86Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ec00ff00cc00)
  ) CLBLL_R_X57Y98_SLICE_X86Y98_BLUT (
.I0(CLBLL_L_X54Y99_SLICE_X83Y99_A5Q),
.I1(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I2(CLBLM_R_X53Y99_SLICE_X81Y99_AQ),
.I3(CLBLM_L_X62Y99_SLICE_X92Y99_AO6),
.I4(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I5(CLBLM_L_X56Y99_SLICE_X85Y99_A5Q),
.O5(CLBLL_R_X57Y98_SLICE_X86Y98_BO5),
.O6(CLBLL_R_X57Y98_SLICE_X86Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ed00ff00dc00)
  ) CLBLL_R_X57Y98_SLICE_X86Y98_ALUT (
.I0(CLBLL_L_X54Y99_SLICE_X83Y99_A5Q),
.I1(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I2(CLBLM_R_X53Y99_SLICE_X81Y99_AQ),
.I3(CLBLM_L_X62Y99_SLICE_X92Y99_AO6),
.I4(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I5(CLBLM_L_X56Y99_SLICE_X85Y99_A5Q),
.O5(CLBLL_R_X57Y98_SLICE_X86Y98_AO5),
.O6(CLBLL_R_X57Y98_SLICE_X86Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X57Y98_SLICE_X87Y98_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_R_X57Y97_SLICE_X87Y97_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y98_SLICE_X89Y98_AQ),
.Q(CLBLL_R_X57Y98_SLICE_X87Y98_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X57Y98_SLICE_X87Y98_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_R_X57Y97_SLICE_X87Y97_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y98_SLICE_X89Y98_A5Q),
.Q(CLBLL_R_X57Y98_SLICE_X87Y98_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X57Y98_SLICE_X87Y98_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_R_X57Y97_SLICE_X87Y97_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y98_SLICE_X89Y98_CQ),
.Q(CLBLL_R_X57Y98_SLICE_X87Y98_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X57Y98_SLICE_X87Y98_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_R_X57Y97_SLICE_X87Y97_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y98_SLICE_X89Y98_C5Q),
.Q(CLBLL_R_X57Y98_SLICE_X87Y98_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y98_SLICE_X87Y98_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y98_SLICE_X87Y98_DO5),
.O6(CLBLL_R_X57Y98_SLICE_X87Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y98_SLICE_X87Y98_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y98_SLICE_X87Y98_CO5),
.O6(CLBLL_R_X57Y98_SLICE_X87Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y98_SLICE_X87Y98_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y98_SLICE_X87Y98_BO5),
.O6(CLBLL_R_X57Y98_SLICE_X87Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y98_SLICE_X87Y98_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y98_SLICE_X87Y98_AO5),
.O6(CLBLL_R_X57Y98_SLICE_X87Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLL_R_X57Y99_SLICE_X86Y99_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_R_X57Y100_SLICE_X87Y100_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_R_X57Y99_SLICE_X86Y99_AO6),
.Q(CLBLL_R_X57Y99_SLICE_X86Y99_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLL_R_X57Y99_SLICE_X86Y99_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_R_X57Y100_SLICE_X87Y100_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_R_X57Y99_SLICE_X86Y99_BO6),
.Q(CLBLL_R_X57Y99_SLICE_X86Y99_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y99_SLICE_X86Y99_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y99_SLICE_X86Y99_DO5),
.O6(CLBLL_R_X57Y99_SLICE_X86Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y99_SLICE_X86Y99_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y99_SLICE_X86Y99_CO5),
.O6(CLBLL_R_X57Y99_SLICE_X86Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa3ffa300a3f0a30)
  ) CLBLL_R_X57Y99_SLICE_X86Y99_BLUT (
.I0(CLBLL_R_X57Y101_SLICE_X87Y101_BO5),
.I1(CLBLM_L_X56Y98_SLICE_X84Y98_BQ),
.I2(CLBLM_L_X56Y99_SLICE_X85Y99_BQ),
.I3(CLBLL_L_X54Y99_SLICE_X82Y99_CQ),
.I4(CLBLM_R_X59Y96_SLICE_X89Y96_A5Q),
.I5(CLBLM_L_X62Y101_SLICE_X93Y101_CQ),
.O5(CLBLL_R_X57Y99_SLICE_X86Y99_BO5),
.O6(CLBLL_R_X57Y99_SLICE_X86Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaccf0ffaaccf0)
  ) CLBLL_R_X57Y99_SLICE_X86Y99_ALUT (
.I0(CLBLL_R_X57Y101_SLICE_X87Y101_BO5),
.I1(CLBLM_L_X56Y98_SLICE_X84Y98_BQ),
.I2(CLBLM_R_X59Y96_SLICE_X89Y96_A5Q),
.I3(CLBLL_L_X54Y99_SLICE_X82Y99_AQ),
.I4(CLBLL_L_X54Y98_SLICE_X83Y98_BQ),
.I5(1'b1),
.O5(CLBLL_R_X57Y99_SLICE_X86Y99_AO5),
.O6(CLBLL_R_X57Y99_SLICE_X86Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLL_R_X57Y99_SLICE_X87Y99_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_R_X57Y99_SLICE_X87Y99_AO6),
.Q(CLBLL_R_X57Y99_SLICE_X87Y99_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y99_SLICE_X87Y99_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y99_SLICE_X87Y99_DO5),
.O6(CLBLL_R_X57Y99_SLICE_X87Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3030303030303030)
  ) CLBLL_R_X57Y99_SLICE_X87Y99_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X56Y99_SLICE_X85Y99_BQ),
.I2(CLBLL_L_X54Y99_SLICE_X82Y99_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y99_SLICE_X87Y99_CO5),
.O6(CLBLL_R_X57Y99_SLICE_X87Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he0e0e0e0e0e0e0e0)
  ) CLBLL_R_X57Y99_SLICE_X87Y99_BLUT (
.I0(CLBLM_L_X56Y99_SLICE_X84Y99_BQ),
.I1(CLBLM_L_X56Y99_SLICE_X84Y99_AQ),
.I2(CLBLM_L_X60Y98_SLICE_X91Y98_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y99_SLICE_X87Y99_BO5),
.O6(CLBLL_R_X57Y99_SLICE_X87Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaf0aaffaac0aa)
  ) CLBLL_R_X57Y99_SLICE_X87Y99_ALUT (
.I0(CLBLL_R_X57Y99_SLICE_X87Y99_AQ),
.I1(CLBLL_R_X57Y100_SLICE_X86Y100_AO6),
.I2(CLBLM_R_X59Y100_SLICE_X88Y100_AO6),
.I3(CLBLM_L_X62Y99_SLICE_X92Y99_AO6),
.I4(CLBLM_L_X60Y98_SLICE_X90Y98_CO5),
.I5(CLBLL_R_X57Y99_SLICE_X87Y99_CO6),
.O5(CLBLL_R_X57Y99_SLICE_X87Y99_AO5),
.O6(CLBLL_R_X57Y99_SLICE_X87Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLL_R_X57Y100_SLICE_X86Y100_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLL_R_X57Y100_SLICE_X87Y100_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_R_X57Y100_SLICE_X86Y100_AO5),
.Q(CLBLL_R_X57Y100_SLICE_X86Y100_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLL_R_X57Y100_SLICE_X86Y100_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLL_R_X57Y100_SLICE_X87Y100_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_R_X57Y100_SLICE_X86Y100_BO6),
.Q(CLBLL_R_X57Y100_SLICE_X86Y100_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLL_R_X57Y100_SLICE_X86Y100_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLL_R_X57Y100_SLICE_X87Y100_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_R_X57Y100_SLICE_X86Y100_CO6),
.Q(CLBLL_R_X57Y100_SLICE_X86Y100_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLL_R_X57Y100_SLICE_X86Y100_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLL_R_X57Y100_SLICE_X87Y100_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_R_X57Y100_SLICE_X86Y100_DO6),
.Q(CLBLL_R_X57Y100_SLICE_X86Y100_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00aaaa0f0fcccc)
  ) CLBLL_R_X57Y100_SLICE_X86Y100_DLUT (
.I0(CLBLM_L_X60Y100_SLICE_X90Y100_AO6),
.I1(CLBLM_R_X59Y98_SLICE_X89Y98_AQ),
.I2(CLBLM_L_X56Y98_SLICE_X84Y98_AQ),
.I3(CLBLM_L_X62Y100_SLICE_X92Y100_AQ),
.I4(CLBLM_L_X56Y99_SLICE_X85Y99_BQ),
.I5(CLBLL_L_X54Y99_SLICE_X82Y99_CQ),
.O5(CLBLL_R_X57Y100_SLICE_X86Y100_DO5),
.O6(CLBLL_R_X57Y100_SLICE_X86Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e45500e4e4ffaa)
  ) CLBLL_R_X57Y100_SLICE_X86Y100_CLUT (
.I0(CLBLM_L_X56Y99_SLICE_X85Y99_BQ),
.I1(CLBLM_L_X60Y100_SLICE_X90Y100_AO5),
.I2(CLBLM_L_X62Y100_SLICE_X92Y100_BQ),
.I3(CLBLM_R_X59Y98_SLICE_X89Y98_A5Q),
.I4(CLBLL_L_X54Y99_SLICE_X82Y99_CQ),
.I5(CLBLM_L_X56Y100_SLICE_X85Y100_AQ),
.O5(CLBLL_R_X57Y100_SLICE_X86Y100_CO5),
.O6(CLBLL_R_X57Y100_SLICE_X86Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffaafaaf5f0a5a0)
  ) CLBLL_R_X57Y100_SLICE_X86Y100_BLUT (
.I0(CLBLL_L_X54Y99_SLICE_X82Y99_AQ),
.I1(1'b1),
.I2(CLBLL_L_X54Y98_SLICE_X83Y98_BQ),
.I3(CLBLM_R_X59Y98_SLICE_X89Y98_A5Q),
.I4(CLBLM_L_X60Y100_SLICE_X90Y100_AO5),
.I5(CLBLM_L_X56Y100_SLICE_X85Y100_AQ),
.O5(CLBLL_R_X57Y100_SLICE_X86Y100_BO5),
.O6(CLBLL_R_X57Y100_SLICE_X86Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55550000fafaee44)
  ) CLBLL_R_X57Y100_SLICE_X86Y100_ALUT (
.I0(CLBLL_L_X54Y99_SLICE_X82Y99_AQ),
.I1(CLBLM_R_X59Y98_SLICE_X89Y98_AQ),
.I2(CLBLM_L_X60Y100_SLICE_X90Y100_AO6),
.I3(CLBLM_L_X56Y98_SLICE_X84Y98_AQ),
.I4(CLBLL_L_X54Y98_SLICE_X83Y98_BQ),
.I5(1'b1),
.O5(CLBLL_R_X57Y100_SLICE_X86Y100_AO5),
.O6(CLBLL_R_X57Y100_SLICE_X86Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLL_R_X57Y100_SLICE_X87Y100_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLL_R_X57Y100_SLICE_X87Y100_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_R_X57Y100_SLICE_X87Y100_AO6),
.Q(CLBLL_R_X57Y100_SLICE_X87Y100_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLL_R_X57Y100_SLICE_X87Y100_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLL_R_X57Y100_SLICE_X87Y100_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_R_X57Y100_SLICE_X87Y100_BO6),
.Q(CLBLL_R_X57Y100_SLICE_X87Y100_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLL_R_X57Y100_SLICE_X87Y100_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLL_R_X57Y100_SLICE_X87Y100_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_R_X57Y100_SLICE_X87Y100_CO6),
.Q(CLBLL_R_X57Y100_SLICE_X87Y100_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00cc00cc00)
  ) CLBLL_R_X57Y100_SLICE_X87Y100_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X60Y98_SLICE_X91Y98_BQ),
.I2(1'b1),
.I3(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y100_SLICE_X87Y100_DO5),
.O6(CLBLL_R_X57Y100_SLICE_X87Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00ff33e2e2e2e2)
  ) CLBLL_R_X57Y100_SLICE_X87Y100_CLUT (
.I0(CLBLM_R_X59Y98_SLICE_X89Y98_B5Q),
.I1(CLBLL_L_X54Y99_SLICE_X82Y99_CQ),
.I2(CLBLM_L_X60Y101_SLICE_X91Y101_CO5),
.I3(CLBLM_L_X62Y100_SLICE_X92Y100_CQ),
.I4(CLBLM_L_X56Y100_SLICE_X85Y100_BQ),
.I5(CLBLM_L_X56Y99_SLICE_X85Y99_BQ),
.O5(CLBLL_R_X57Y100_SLICE_X87Y100_CO5),
.O6(CLBLL_R_X57Y100_SLICE_X87Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff0f0cacacaca)
  ) CLBLL_R_X57Y100_SLICE_X87Y100_BLUT (
.I0(CLBLM_R_X59Y96_SLICE_X89Y96_AQ),
.I1(CLBLL_R_X57Y101_SLICE_X87Y101_BO6),
.I2(CLBLL_L_X54Y98_SLICE_X83Y98_BQ),
.I3(1'b1),
.I4(CLBLM_L_X56Y100_SLICE_X85Y100_DQ),
.I5(CLBLL_L_X54Y99_SLICE_X82Y99_AQ),
.O5(CLBLL_R_X57Y100_SLICE_X87Y100_BO5),
.O6(CLBLL_R_X57Y100_SLICE_X87Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff0f0fc0cfc0c)
  ) CLBLL_R_X57Y100_SLICE_X87Y100_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X59Y98_SLICE_X89Y98_B5Q),
.I2(CLBLL_L_X54Y98_SLICE_X83Y98_BQ),
.I3(CLBLM_L_X60Y101_SLICE_X91Y101_CO5),
.I4(CLBLM_L_X56Y100_SLICE_X85Y100_BQ),
.I5(CLBLL_L_X54Y99_SLICE_X82Y99_AQ),
.O5(CLBLL_R_X57Y100_SLICE_X87Y100_AO5),
.O6(CLBLL_R_X57Y100_SLICE_X87Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X57Y101_SLICE_X86Y101_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y100_SLICE_X90Y100_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_R_X57Y101_SLICE_X86Y101_AO6),
.Q(CLBLL_R_X57Y101_SLICE_X86Y101_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y101_SLICE_X86Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y101_SLICE_X86Y101_DO5),
.O6(CLBLL_R_X57Y101_SLICE_X86Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y101_SLICE_X86Y101_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y101_SLICE_X86Y101_CO5),
.O6(CLBLL_R_X57Y101_SLICE_X86Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccc0ccc088880000)
  ) CLBLL_R_X57Y101_SLICE_X86Y101_BLUT (
.I0(CLBLL_L_X54Y101_SLICE_X83Y101_CO6),
.I1(CLBLM_L_X62Y99_SLICE_X92Y99_AO6),
.I2(CLBLM_L_X60Y99_SLICE_X91Y99_AO5),
.I3(CLBLL_R_X57Y97_SLICE_X86Y97_CO6),
.I4(CLBLL_L_X52Y105_SLICE_X78Y105_AO5),
.I5(CLBLL_R_X57Y101_SLICE_X86Y101_AO5),
.O5(CLBLL_R_X57Y101_SLICE_X86Y101_BO5),
.O6(CLBLL_R_X57Y101_SLICE_X86Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0fcc0fff000000)
  ) CLBLL_R_X57Y101_SLICE_X86Y101_ALUT (
.I0(CLBLM_L_X50Y104_SLICE_X76Y104_AQ),
.I1(CLBLM_R_X49Y104_SLICE_X74Y104_AQ),
.I2(CLBLL_R_X57Y101_SLICE_X86Y101_AQ),
.I3(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I4(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I5(1'b1),
.O5(CLBLL_R_X57Y101_SLICE_X86Y101_AO5),
.O6(CLBLL_R_X57Y101_SLICE_X86Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLL_R_X57Y101_SLICE_X87Y101_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLL_R_X57Y100_SLICE_X87Y100_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_R_X57Y101_SLICE_X87Y101_AO6),
.Q(CLBLL_R_X57Y101_SLICE_X87Y101_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLL_R_X57Y101_SLICE_X87Y101_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLL_R_X57Y100_SLICE_X87Y100_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_R_X57Y101_SLICE_X87Y101_CO6),
.Q(CLBLL_R_X57Y101_SLICE_X87Y101_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLL_R_X57Y101_SLICE_X87Y101_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLL_R_X57Y100_SLICE_X87Y100_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_R_X57Y101_SLICE_X87Y101_DO6),
.Q(CLBLL_R_X57Y101_SLICE_X87Y101_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf377f344c077c044)
  ) CLBLL_R_X57Y101_SLICE_X87Y101_DLUT (
.I0(CLBLM_L_X56Y100_SLICE_X85Y100_DQ),
.I1(CLBLM_L_X56Y99_SLICE_X85Y99_BQ),
.I2(CLBLM_L_X62Y101_SLICE_X93Y101_BQ),
.I3(CLBLL_L_X54Y99_SLICE_X82Y99_CQ),
.I4(CLBLM_R_X59Y96_SLICE_X89Y96_AQ),
.I5(CLBLL_R_X57Y101_SLICE_X87Y101_BO6),
.O5(CLBLL_R_X57Y101_SLICE_X87Y101_DO5),
.O6(CLBLL_R_X57Y101_SLICE_X87Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5fc05fcf50c050c)
  ) CLBLL_R_X57Y101_SLICE_X87Y101_CLUT (
.I0(CLBLL_L_X54Y101_SLICE_X82Y101_BQ),
.I1(CLBLM_R_X59Y98_SLICE_X89Y98_CQ),
.I2(CLBLL_L_X54Y99_SLICE_X82Y99_CQ),
.I3(CLBLM_L_X56Y99_SLICE_X85Y99_BQ),
.I4(CLBLM_L_X64Y100_SLICE_X97Y100_AQ),
.I5(CLBLM_L_X62Y101_SLICE_X92Y101_DO6),
.O5(CLBLL_R_X57Y101_SLICE_X87Y101_CO5),
.O6(CLBLL_R_X57Y101_SLICE_X87Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc3030bb88bb88)
  ) CLBLL_R_X57Y101_SLICE_X87Y101_BLUT (
.I0(CLBLM_L_X62Y101_SLICE_X92Y101_CQ),
.I1(CLBLM_L_X62Y99_SLICE_X92Y99_BQ),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLM_L_X60Y101_SLICE_X91Y101_BQ),
.I5(1'b1),
.O5(CLBLL_R_X57Y101_SLICE_X87Y101_BO5),
.O6(CLBLL_R_X57Y101_SLICE_X87Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcff0cfffc0f0c0)
  ) CLBLL_R_X57Y101_SLICE_X87Y101_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X62Y101_SLICE_X92Y101_DO6),
.I2(CLBLL_L_X54Y98_SLICE_X83Y98_BQ),
.I3(CLBLL_L_X54Y99_SLICE_X82Y99_AQ),
.I4(CLBLL_L_X54Y101_SLICE_X82Y101_BQ),
.I5(CLBLM_R_X59Y98_SLICE_X89Y98_CQ),
.O5(CLBLL_R_X57Y101_SLICE_X87Y101_AO5),
.O6(CLBLL_R_X57Y101_SLICE_X87Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLL_R_X57Y102_SLICE_X86Y102_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_R_X57Y102_SLICE_X86Y102_DO6),
.Q(CLBLL_R_X57Y102_SLICE_X86Y102_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLL_R_X57Y102_SLICE_X86Y102_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_R_X57Y102_SLICE_X86Y102_BO6),
.Q(CLBLL_R_X57Y102_SLICE_X86Y102_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010000000000)
  ) CLBLL_R_X57Y102_SLICE_X86Y102_DLUT (
.I0(CLBLM_R_X49Y106_SLICE_X75Y106_CQ),
.I1(CLBLM_R_X49Y106_SLICE_X75Y106_DQ),
.I2(CLBLM_R_X49Y104_SLICE_X75Y104_DQ),
.I3(CLBLM_R_X49Y104_SLICE_X75Y104_CQ),
.I4(CLBLM_R_X49Y107_SLICE_X75Y107_CQ),
.I5(CLBLM_L_X56Y100_SLICE_X85Y100_BO6),
.O5(CLBLL_R_X57Y102_SLICE_X86Y102_DO5),
.O6(CLBLL_R_X57Y102_SLICE_X86Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffeff)
  ) CLBLL_R_X57Y102_SLICE_X86Y102_CLUT (
.I0(CLBLM_R_X49Y106_SLICE_X75Y106_CQ),
.I1(CLBLM_R_X49Y106_SLICE_X75Y106_DQ),
.I2(CLBLM_R_X49Y104_SLICE_X75Y104_CQ),
.I3(CLBLM_R_X49Y104_SLICE_X75Y104_BQ),
.I4(CLBLM_R_X49Y104_SLICE_X75Y104_DQ),
.I5(CLBLM_R_X49Y107_SLICE_X75Y107_CQ),
.O5(CLBLL_R_X57Y102_SLICE_X86Y102_CO5),
.O6(CLBLL_R_X57Y102_SLICE_X86Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00000000)
  ) CLBLL_R_X57Y102_SLICE_X86Y102_BLUT (
.I0(CLBLL_R_X57Y102_SLICE_X86Y102_DO6),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X49Y104_SLICE_X75Y104_BQ),
.O5(CLBLL_R_X57Y102_SLICE_X86Y102_BO5),
.O6(CLBLL_R_X57Y102_SLICE_X86Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000a0a088888888)
  ) CLBLL_R_X57Y102_SLICE_X86Y102_ALUT (
.I0(CLBLM_R_X49Y104_SLICE_X75Y104_AQ),
.I1(CLBLL_R_X57Y102_SLICE_X86Y102_DO6),
.I2(CLBLM_L_X56Y102_SLICE_X85Y102_BO6),
.I3(1'b1),
.I4(CLBLL_R_X57Y102_SLICE_X86Y102_CO6),
.I5(1'b1),
.O5(CLBLL_R_X57Y102_SLICE_X86Y102_AO5),
.O6(CLBLL_R_X57Y102_SLICE_X86Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y102_SLICE_X87Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y102_SLICE_X87Y102_DO5),
.O6(CLBLL_R_X57Y102_SLICE_X87Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y102_SLICE_X87Y102_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y102_SLICE_X87Y102_CO5),
.O6(CLBLL_R_X57Y102_SLICE_X87Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y102_SLICE_X87Y102_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y102_SLICE_X87Y102_BO5),
.O6(CLBLL_R_X57Y102_SLICE_X87Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y102_SLICE_X87Y102_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y102_SLICE_X87Y102_AO5),
.O6(CLBLL_R_X57Y102_SLICE_X87Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLL_R_X57Y103_SLICE_X86Y103_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(CLBLM_R_X15Y122_SLICE_X20Y122_AO6),
.D(CLBLL_R_X57Y103_SLICE_X86Y103_AO5),
.Q(CLBLL_R_X57Y103_SLICE_X86Y103_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLL_R_X57Y103_SLICE_X86Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(CLBLM_R_X15Y122_SLICE_X20Y122_AO6),
.D(CLBLL_R_X57Y103_SLICE_X86Y103_AO6),
.Q(CLBLL_R_X57Y103_SLICE_X86Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y103_SLICE_X86Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y103_SLICE_X86Y103_DO5),
.O6(CLBLL_R_X57Y103_SLICE_X86Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y103_SLICE_X86Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y103_SLICE_X86Y103_CO5),
.O6(CLBLL_R_X57Y103_SLICE_X86Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y103_SLICE_X86Y103_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y103_SLICE_X86Y103_BO5),
.O6(CLBLL_R_X57Y103_SLICE_X86Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00f0555500cc)
  ) CLBLL_R_X57Y103_SLICE_X86Y103_ALUT (
.I0(CLBLM_R_X49Y119_SLICE_X74Y119_BQ),
.I1(CLBLL_R_X57Y103_SLICE_X86Y103_A5Q),
.I2(CLBLL_R_X57Y103_SLICE_X86Y103_AQ),
.I3(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.I4(CLBLM_R_X49Y119_SLICE_X74Y119_AQ),
.I5(1'b1),
.O5(CLBLL_R_X57Y103_SLICE_X86Y103_AO5),
.O6(CLBLL_R_X57Y103_SLICE_X86Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X57Y103_SLICE_X87Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y100_SLICE_X90Y100_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_R_X57Y103_SLICE_X87Y103_AO6),
.Q(CLBLL_R_X57Y103_SLICE_X87Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y103_SLICE_X87Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y103_SLICE_X87Y103_DO5),
.O6(CLBLL_R_X57Y103_SLICE_X87Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y103_SLICE_X87Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y103_SLICE_X87Y103_CO5),
.O6(CLBLL_R_X57Y103_SLICE_X87Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y103_SLICE_X87Y103_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y103_SLICE_X87Y103_BO5),
.O6(CLBLL_R_X57Y103_SLICE_X87Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ffffdf80)
  ) CLBLL_R_X57Y103_SLICE_X87Y103_ALUT (
.I0(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I1(CLBLL_R_X57Y105_SLICE_X87Y105_D_XOR),
.I2(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I3(CLBLL_R_X57Y106_SLICE_X86Y106_D_XOR),
.I4(CLBLM_L_X62Y102_SLICE_X92Y102_AO5),
.I5(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.O5(CLBLL_R_X57Y103_SLICE_X87Y103_AO5),
.O6(CLBLL_R_X57Y103_SLICE_X87Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X57Y104_SLICE_X86Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X56Y103_SLICE_X85Y103_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_R_X57Y104_SLICE_X86Y104_AO6),
.Q(CLBLL_R_X57Y104_SLICE_X86Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X57Y104_SLICE_X86Y104_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X56Y103_SLICE_X85Y103_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_R_X57Y104_SLICE_X86Y104_BO6),
.Q(CLBLL_R_X57Y104_SLICE_X86Y104_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X57Y104_SLICE_X86Y104_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X56Y103_SLICE_X85Y103_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_R_X57Y104_SLICE_X86Y104_CO6),
.Q(CLBLL_R_X57Y104_SLICE_X86Y104_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f555500ff3333)
  ) CLBLL_R_X57Y104_SLICE_X86Y104_DLUT (
.I0(CLBLL_R_X57Y104_SLICE_X86Y104_BQ),
.I1(CLBLL_R_X57Y104_SLICE_X86Y104_AQ),
.I2(CLBLL_R_X57Y101_SLICE_X86Y101_AQ),
.I3(CLBLM_L_X60Y108_SLICE_X91Y108_AQ),
.I4(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I5(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.O5(CLBLL_R_X57Y104_SLICE_X86Y104_DO5),
.O6(CLBLL_R_X57Y104_SLICE_X86Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000d8d8d8d8)
  ) CLBLL_R_X57Y104_SLICE_X86Y104_CLUT (
.I0(CLBLL_L_X54Y101_SLICE_X83Y101_BO6),
.I1(CLBLL_R_X57Y104_SLICE_X86Y104_CQ),
.I2(CLBLM_R_X53Y103_SLICE_X81Y103_B_XOR),
.I3(1'b1),
.I4(CLBLM_L_X50Y105_SLICE_X77Y105_AQ),
.I5(CLBLM_L_X62Y100_SLICE_X92Y100_AO5),
.O5(CLBLL_R_X57Y104_SLICE_X86Y104_CO5),
.O6(CLBLL_R_X57Y104_SLICE_X86Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cff0ffc0cf000)
  ) CLBLL_R_X57Y104_SLICE_X86Y104_BLUT (
.I0(1'b1),
.I1(CLBLL_R_X57Y104_SLICE_X86Y104_BQ),
.I2(CLBLM_L_X62Y100_SLICE_X92Y100_AO5),
.I3(CLBLM_L_X50Y104_SLICE_X76Y104_AQ),
.I4(CLBLL_L_X54Y101_SLICE_X83Y101_BO6),
.I5(CLBLM_R_X53Y103_SLICE_X81Y103_A_XOR),
.O5(CLBLL_R_X57Y104_SLICE_X86Y104_BO5),
.O6(CLBLL_R_X57Y104_SLICE_X86Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00f0f0aaaa)
  ) CLBLL_R_X57Y104_SLICE_X86Y104_ALUT (
.I0(CLBLL_L_X54Y106_SLICE_X82Y106_B_XOR),
.I1(1'b1),
.I2(CLBLL_R_X57Y104_SLICE_X86Y104_AQ),
.I3(CLBLM_L_X50Y104_SLICE_X76Y104_AQ),
.I4(CLBLL_L_X54Y101_SLICE_X83Y101_BO6),
.I5(CLBLM_L_X60Y99_SLICE_X90Y99_AO5),
.O5(CLBLL_R_X57Y104_SLICE_X86Y104_AO5),
.O6(CLBLL_R_X57Y104_SLICE_X86Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X57Y104_SLICE_X87Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X56Y103_SLICE_X85Y103_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_R_X57Y104_SLICE_X87Y104_AO6),
.Q(CLBLL_R_X57Y104_SLICE_X87Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X57Y104_SLICE_X87Y104_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X56Y103_SLICE_X85Y103_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_R_X57Y104_SLICE_X87Y104_BO6),
.Q(CLBLL_R_X57Y104_SLICE_X87Y104_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X57Y104_SLICE_X87Y104_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X56Y103_SLICE_X85Y103_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_R_X57Y104_SLICE_X87Y104_CO6),
.Q(CLBLL_R_X57Y104_SLICE_X87Y104_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5300530f53f053ff)
  ) CLBLL_R_X57Y104_SLICE_X87Y104_DLUT (
.I0(CLBLL_R_X57Y105_SLICE_X86Y105_AQ),
.I1(CLBLL_R_X57Y104_SLICE_X87Y104_CQ),
.I2(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I3(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I4(CLBLL_R_X57Y104_SLICE_X87Y104_AQ),
.I5(CLBLL_R_X57Y109_SLICE_X86Y109_BQ),
.O5(CLBLL_R_X57Y104_SLICE_X87Y104_DO5),
.O6(CLBLL_R_X57Y104_SLICE_X87Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00d8d8d8d8)
  ) CLBLL_R_X57Y104_SLICE_X87Y104_CLUT (
.I0(CLBLL_L_X54Y101_SLICE_X83Y101_BO6),
.I1(CLBLL_R_X57Y104_SLICE_X87Y104_CQ),
.I2(CLBLM_R_X53Y103_SLICE_X81Y103_C_XOR),
.I3(CLBLM_R_X49Y105_SLICE_X75Y105_CQ),
.I4(1'b1),
.I5(CLBLM_L_X62Y100_SLICE_X92Y100_AO5),
.O5(CLBLL_R_X57Y104_SLICE_X87Y104_CO5),
.O6(CLBLL_R_X57Y104_SLICE_X87Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hefefeaea45454040)
  ) CLBLL_R_X57Y104_SLICE_X87Y104_BLUT (
.I0(CLBLM_L_X60Y99_SLICE_X90Y99_AO5),
.I1(CLBLL_R_X57Y104_SLICE_X87Y104_BQ),
.I2(CLBLL_L_X54Y101_SLICE_X83Y101_BO6),
.I3(1'b1),
.I4(CLBLL_L_X54Y108_SLICE_X82Y108_A_XOR),
.I5(CLBLM_L_X50Y107_SLICE_X77Y107_AQ),
.O5(CLBLL_R_X57Y104_SLICE_X87Y104_BO5),
.O6(CLBLL_R_X57Y104_SLICE_X87Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcffcc30303300)
  ) CLBLL_R_X57Y104_SLICE_X87Y104_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X60Y99_SLICE_X90Y99_AO5),
.I2(CLBLL_R_X57Y104_SLICE_X87Y104_AQ),
.I3(CLBLL_L_X54Y106_SLICE_X82Y106_D_XOR),
.I4(CLBLL_L_X54Y101_SLICE_X83Y101_BO6),
.I5(CLBLM_R_X49Y105_SLICE_X75Y105_CQ),
.O5(CLBLL_R_X57Y104_SLICE_X87Y104_AO5),
.O6(CLBLL_R_X57Y104_SLICE_X87Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X57Y105_SLICE_X86Y105_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y100_SLICE_X90Y100_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_R_X57Y105_SLICE_X86Y105_AO6),
.Q(CLBLL_R_X57Y105_SLICE_X86Y105_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X57Y105_SLICE_X86Y105_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y100_SLICE_X90Y100_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_R_X57Y105_SLICE_X86Y105_BO6),
.Q(CLBLL_R_X57Y105_SLICE_X86Y105_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h407043734c7c4f7f)
  ) CLBLL_R_X57Y105_SLICE_X86Y105_DLUT (
.I0(CLBLL_R_X57Y105_SLICE_X86Y105_BQ),
.I1(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I2(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I3(CLBLL_R_X57Y109_SLICE_X86Y109_CQ),
.I4(CLBLM_L_X56Y105_SLICE_X84Y105_AQ),
.I5(CLBLM_L_X56Y105_SLICE_X85Y105_DQ),
.O5(CLBLL_R_X57Y105_SLICE_X86Y105_DO5),
.O6(CLBLL_R_X57Y105_SLICE_X86Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfece3e0ef2c23202)
  ) CLBLL_R_X57Y105_SLICE_X86Y105_CLUT (
.I0(CLBLM_L_X56Y105_SLICE_X85Y105_AQ),
.I1(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I2(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I3(CLBLL_R_X57Y104_SLICE_X86Y104_CQ),
.I4(CLBLM_R_X59Y106_SLICE_X88Y106_BQ),
.I5(CLBLL_R_X57Y109_SLICE_X86Y109_AQ),
.O5(CLBLL_R_X57Y105_SLICE_X86Y105_CO5),
.O6(CLBLL_R_X57Y105_SLICE_X86Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000fffff780)
  ) CLBLL_R_X57Y105_SLICE_X86Y105_BLUT (
.I0(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I1(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I2(CLBLL_R_X57Y105_SLICE_X87Y105_C_XOR),
.I3(CLBLL_R_X57Y106_SLICE_X86Y106_C_XOR),
.I4(CLBLM_L_X62Y98_SLICE_X92Y98_AO6),
.I5(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.O5(CLBLL_R_X57Y105_SLICE_X86Y105_BO5),
.O6(CLBLL_R_X57Y105_SLICE_X86Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccfdffeccc)
  ) CLBLL_R_X57Y105_SLICE_X86Y105_ALUT (
.I0(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I1(CLBLM_L_X62Y105_SLICE_X92Y105_AO6),
.I2(CLBLL_R_X57Y105_SLICE_X87Y105_B_XOR),
.I3(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I4(CLBLL_R_X57Y106_SLICE_X86Y106_B_XOR),
.I5(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.O5(CLBLL_R_X57Y105_SLICE_X86Y105_AO5),
.O6(CLBLL_R_X57Y105_SLICE_X86Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_R_X57Y105_SLICE_X87Y105_CARRY4 (
.CI(1'b0),
.CO({CLBLL_R_X57Y105_SLICE_X87Y105_D_CY, CLBLL_R_X57Y105_SLICE_X87Y105_C_CY, CLBLL_R_X57Y105_SLICE_X87Y105_B_CY, CLBLL_R_X57Y105_SLICE_X87Y105_A_CY}),
.CYINIT(CLBLL_R_X57Y101_SLICE_X86Y101_AQ),
.DI({CLBLL_R_X57Y103_SLICE_X87Y103_AQ, CLBLL_R_X57Y105_SLICE_X86Y105_BQ, CLBLL_R_X57Y105_SLICE_X86Y105_AQ, CLBLL_R_X57Y105_SLICE_X87Y105_AO5}),
.O({CLBLL_R_X57Y105_SLICE_X87Y105_D_XOR, CLBLL_R_X57Y105_SLICE_X87Y105_C_XOR, CLBLL_R_X57Y105_SLICE_X87Y105_B_XOR, CLBLL_R_X57Y105_SLICE_X87Y105_A_XOR}),
.S({CLBLL_R_X57Y105_SLICE_X87Y105_DO6, CLBLL_R_X57Y105_SLICE_X87Y105_CO6, CLBLL_R_X57Y105_SLICE_X87Y105_BO6, CLBLL_R_X57Y105_SLICE_X87Y105_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555555)
  ) CLBLL_R_X57Y105_SLICE_X87Y105_DLUT (
.I0(CLBLL_R_X57Y103_SLICE_X87Y103_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y105_SLICE_X87Y105_DO5),
.O6(CLBLL_R_X57Y105_SLICE_X87Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffffffff)
  ) CLBLL_R_X57Y105_SLICE_X87Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_R_X57Y105_SLICE_X86Y105_BQ),
.O5(CLBLL_R_X57Y105_SLICE_X87Y105_CO5),
.O6(CLBLL_R_X57Y105_SLICE_X87Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffff0000ffff)
  ) CLBLL_R_X57Y105_SLICE_X87Y105_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_R_X57Y105_SLICE_X86Y105_AQ),
.I5(1'b1),
.O5(CLBLL_R_X57Y105_SLICE_X87Y105_BO5),
.O6(CLBLL_R_X57Y105_SLICE_X87Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ffff00ff00)
  ) CLBLL_R_X57Y105_SLICE_X87Y105_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X59Y106_SLICE_X88Y106_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y105_SLICE_X87Y105_AO5),
.O6(CLBLL_R_X57Y105_SLICE_X87Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_R_X57Y106_SLICE_X86Y106_CARRY4 (
.CI(1'b0),
.CO({CLBLL_R_X57Y106_SLICE_X86Y106_D_CY, CLBLL_R_X57Y106_SLICE_X86Y106_C_CY, CLBLL_R_X57Y106_SLICE_X86Y106_B_CY, CLBLL_R_X57Y106_SLICE_X86Y106_A_CY}),
.CYINIT(CLBLL_R_X57Y101_SLICE_X86Y101_AQ),
.DI({1'b0, 1'b0, 1'b0, CLBLL_R_X57Y106_SLICE_X86Y106_AO5}),
.O({CLBLL_R_X57Y106_SLICE_X86Y106_D_XOR, CLBLL_R_X57Y106_SLICE_X86Y106_C_XOR, CLBLL_R_X57Y106_SLICE_X86Y106_B_XOR, CLBLL_R_X57Y106_SLICE_X86Y106_A_XOR}),
.S({CLBLL_R_X57Y106_SLICE_X86Y106_DO6, CLBLL_R_X57Y106_SLICE_X86Y106_CO6, CLBLL_R_X57Y106_SLICE_X86Y106_BO6, CLBLL_R_X57Y106_SLICE_X86Y106_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLL_R_X57Y106_SLICE_X86Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_R_X57Y103_SLICE_X87Y103_AQ),
.O5(CLBLL_R_X57Y106_SLICE_X86Y106_DO5),
.O6(CLBLL_R_X57Y106_SLICE_X86Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLL_R_X57Y106_SLICE_X86Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_R_X57Y105_SLICE_X86Y105_BQ),
.O5(CLBLL_R_X57Y106_SLICE_X86Y106_CO5),
.O6(CLBLL_R_X57Y106_SLICE_X86Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLL_R_X57Y106_SLICE_X86Y106_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_R_X57Y105_SLICE_X86Y105_AQ),
.O5(CLBLL_R_X57Y106_SLICE_X86Y106_BO5),
.O6(CLBLL_R_X57Y106_SLICE_X86Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0000000000)
  ) CLBLL_R_X57Y106_SLICE_X86Y106_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X59Y106_SLICE_X88Y106_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y106_SLICE_X86Y106_AO5),
.O6(CLBLL_R_X57Y106_SLICE_X86Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLL_R_X57Y106_SLICE_X87Y106_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLL_R_X57Y99_SLICE_X87Y99_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_R_X57Y106_SLICE_X87Y106_AO5),
.Q(CLBLL_R_X57Y106_SLICE_X87Y106_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_R_X57Y106_SLICE_X87Y106_CARRY4 (
.CI(CLBLL_R_X57Y105_SLICE_X87Y105_COUT),
.CO({CLBLL_R_X57Y106_SLICE_X87Y106_D_CY, CLBLL_R_X57Y106_SLICE_X87Y106_C_CY, CLBLL_R_X57Y106_SLICE_X87Y106_B_CY, CLBLL_R_X57Y106_SLICE_X87Y106_A_CY}),
.CYINIT(1'b0),
.DI({CLBLM_L_X60Y108_SLICE_X91Y108_AQ, CLBLM_R_X59Y106_SLICE_X88Y106_AQ, CLBLL_R_X57Y108_SLICE_X87Y108_BQ, CLBLL_R_X57Y108_SLICE_X87Y108_AQ}),
.O({CLBLL_R_X57Y106_SLICE_X87Y106_D_XOR, CLBLL_R_X57Y106_SLICE_X87Y106_C_XOR, CLBLL_R_X57Y106_SLICE_X87Y106_B_XOR, CLBLL_R_X57Y106_SLICE_X87Y106_A_XOR}),
.S({CLBLL_R_X57Y106_SLICE_X87Y106_DO6, CLBLL_R_X57Y106_SLICE_X87Y106_CO6, CLBLL_R_X57Y106_SLICE_X87Y106_BO6, CLBLL_R_X57Y106_SLICE_X87Y106_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333333333333)
  ) CLBLL_R_X57Y106_SLICE_X87Y106_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X60Y108_SLICE_X91Y108_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y106_SLICE_X87Y106_DO5),
.O6(CLBLL_R_X57Y106_SLICE_X87Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555555)
  ) CLBLL_R_X57Y106_SLICE_X87Y106_CLUT (
.I0(CLBLM_R_X59Y106_SLICE_X88Y106_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y106_SLICE_X87Y106_CO5),
.O6(CLBLL_R_X57Y106_SLICE_X87Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333333333333)
  ) CLBLL_R_X57Y106_SLICE_X87Y106_BLUT (
.I0(1'b1),
.I1(CLBLL_R_X57Y108_SLICE_X87Y108_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y106_SLICE_X87Y106_BO5),
.O6(CLBLL_R_X57Y106_SLICE_X87Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffffff00ff00)
  ) CLBLL_R_X57Y106_SLICE_X87Y106_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X49Y106_SLICE_X75Y106_DQ),
.I4(CLBLL_R_X57Y108_SLICE_X87Y108_AQ),
.I5(1'b1),
.O5(CLBLL_R_X57Y106_SLICE_X87Y106_AO5),
.O6(CLBLL_R_X57Y106_SLICE_X87Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_R_X57Y107_SLICE_X86Y107_CARRY4 (
.CI(CLBLL_R_X57Y106_SLICE_X86Y106_COUT),
.CO({CLBLL_R_X57Y107_SLICE_X86Y107_D_CY, CLBLL_R_X57Y107_SLICE_X86Y107_C_CY, CLBLL_R_X57Y107_SLICE_X86Y107_B_CY, CLBLL_R_X57Y107_SLICE_X86Y107_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLL_R_X57Y107_SLICE_X86Y107_D_XOR, CLBLL_R_X57Y107_SLICE_X86Y107_C_XOR, CLBLL_R_X57Y107_SLICE_X86Y107_B_XOR, CLBLL_R_X57Y107_SLICE_X86Y107_A_XOR}),
.S({CLBLL_R_X57Y107_SLICE_X86Y107_DO6, CLBLL_R_X57Y107_SLICE_X86Y107_CO6, CLBLL_R_X57Y107_SLICE_X86Y107_BO6, CLBLL_R_X57Y107_SLICE_X86Y107_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLL_R_X57Y107_SLICE_X86Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X60Y108_SLICE_X91Y108_AQ),
.O5(CLBLL_R_X57Y107_SLICE_X86Y107_DO5),
.O6(CLBLL_R_X57Y107_SLICE_X86Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLL_R_X57Y107_SLICE_X86Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X59Y106_SLICE_X88Y106_AQ),
.O5(CLBLL_R_X57Y107_SLICE_X86Y107_CO5),
.O6(CLBLL_R_X57Y107_SLICE_X86Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLL_R_X57Y107_SLICE_X86Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_R_X57Y108_SLICE_X87Y108_BQ),
.O5(CLBLL_R_X57Y107_SLICE_X86Y107_BO5),
.O6(CLBLL_R_X57Y107_SLICE_X86Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLL_R_X57Y107_SLICE_X86Y107_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_R_X57Y108_SLICE_X87Y108_AQ),
.O5(CLBLL_R_X57Y107_SLICE_X86Y107_AO5),
.O6(CLBLL_R_X57Y107_SLICE_X86Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_R_X57Y107_SLICE_X87Y107_CARRY4 (
.CI(CLBLL_R_X57Y106_SLICE_X87Y106_COUT),
.CO({CLBLL_R_X57Y107_SLICE_X87Y107_D_CY, CLBLL_R_X57Y107_SLICE_X87Y107_C_CY, CLBLL_R_X57Y107_SLICE_X87Y107_B_CY, CLBLL_R_X57Y107_SLICE_X87Y107_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, CLBLL_R_X57Y109_SLICE_X86Y109_BQ, CLBLL_R_X57Y109_SLICE_X86Y109_AQ}),
.O({CLBLL_R_X57Y107_SLICE_X87Y107_D_XOR, CLBLL_R_X57Y107_SLICE_X87Y107_C_XOR, CLBLL_R_X57Y107_SLICE_X87Y107_B_XOR, CLBLL_R_X57Y107_SLICE_X87Y107_A_XOR}),
.S({CLBLL_R_X57Y107_SLICE_X87Y107_DO6, CLBLL_R_X57Y107_SLICE_X87Y107_CO6, CLBLL_R_X57Y107_SLICE_X87Y107_BO6, CLBLL_R_X57Y107_SLICE_X87Y107_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y107_SLICE_X87Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y107_SLICE_X87Y107_DO5),
.O6(CLBLL_R_X57Y107_SLICE_X87Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00ff00ff)
  ) CLBLL_R_X57Y107_SLICE_X87Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_R_X57Y109_SLICE_X86Y109_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y107_SLICE_X87Y107_CO5),
.O6(CLBLL_R_X57Y107_SLICE_X87Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555555)
  ) CLBLL_R_X57Y107_SLICE_X87Y107_BLUT (
.I0(CLBLL_R_X57Y109_SLICE_X86Y109_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y107_SLICE_X87Y107_BO5),
.O6(CLBLL_R_X57Y107_SLICE_X87Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00ff00ff)
  ) CLBLL_R_X57Y107_SLICE_X87Y107_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_R_X57Y109_SLICE_X86Y109_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y107_SLICE_X87Y107_AO5),
.O6(CLBLL_R_X57Y107_SLICE_X87Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_R_X57Y108_SLICE_X86Y108_CARRY4 (
.CI(CLBLL_R_X57Y107_SLICE_X86Y107_COUT),
.CO({CLBLL_R_X57Y108_SLICE_X86Y108_D_CY, CLBLL_R_X57Y108_SLICE_X86Y108_C_CY, CLBLL_R_X57Y108_SLICE_X86Y108_B_CY, CLBLL_R_X57Y108_SLICE_X86Y108_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLL_R_X57Y108_SLICE_X86Y108_D_XOR, CLBLL_R_X57Y108_SLICE_X86Y108_C_XOR, CLBLL_R_X57Y108_SLICE_X86Y108_B_XOR, CLBLL_R_X57Y108_SLICE_X86Y108_A_XOR}),
.S({CLBLL_R_X57Y108_SLICE_X86Y108_DO6, CLBLL_R_X57Y108_SLICE_X86Y108_CO6, CLBLL_R_X57Y108_SLICE_X86Y108_BO6, CLBLL_R_X57Y108_SLICE_X86Y108_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y108_SLICE_X86Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y108_SLICE_X86Y108_DO5),
.O6(CLBLL_R_X57Y108_SLICE_X86Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLL_R_X57Y108_SLICE_X86Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_R_X57Y109_SLICE_X86Y109_CQ),
.O5(CLBLL_R_X57Y108_SLICE_X86Y108_CO5),
.O6(CLBLL_R_X57Y108_SLICE_X86Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLL_R_X57Y108_SLICE_X86Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_R_X57Y109_SLICE_X86Y109_BQ),
.O5(CLBLL_R_X57Y108_SLICE_X86Y108_BO5),
.O6(CLBLL_R_X57Y108_SLICE_X86Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLL_R_X57Y108_SLICE_X86Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_R_X57Y109_SLICE_X86Y109_AQ),
.O5(CLBLL_R_X57Y108_SLICE_X86Y108_AO5),
.O6(CLBLL_R_X57Y108_SLICE_X86Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X57Y108_SLICE_X87Y108_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y100_SLICE_X90Y100_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_R_X57Y108_SLICE_X87Y108_AO6),
.Q(CLBLL_R_X57Y108_SLICE_X87Y108_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X57Y108_SLICE_X87Y108_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y100_SLICE_X90Y100_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_R_X57Y108_SLICE_X87Y108_BO6),
.Q(CLBLL_R_X57Y108_SLICE_X87Y108_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33cc00e2e2e2e2)
  ) CLBLL_R_X57Y108_SLICE_X87Y108_DLUT (
.I0(CLBLL_R_X57Y106_SLICE_X87Y106_AQ),
.I1(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I2(CLBLL_R_X57Y110_SLICE_X87Y110_C_XOR),
.I3(CLBLL_R_X57Y108_SLICE_X87Y108_BQ),
.I4(CLBLL_R_X57Y107_SLICE_X86Y107_B_XOR),
.I5(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.O5(CLBLL_R_X57Y108_SLICE_X87Y108_DO5),
.O6(CLBLL_R_X57Y108_SLICE_X87Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0f0aaaaff00)
  ) CLBLL_R_X57Y108_SLICE_X87Y108_CLUT (
.I0(CLBLL_R_X57Y109_SLICE_X87Y109_C_XOR),
.I1(CLBLL_R_X57Y105_SLICE_X86Y105_AQ),
.I2(CLBLL_R_X57Y106_SLICE_X86Y106_B_XOR),
.I3(CLBLM_R_X59Y103_SLICE_X88Y103_DQ),
.I4(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I5(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.O5(CLBLL_R_X57Y108_SLICE_X87Y108_CO5),
.O6(CLBLL_R_X57Y108_SLICE_X87Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3202ffff2222)
  ) CLBLL_R_X57Y108_SLICE_X87Y108_BLUT (
.I0(CLBLL_R_X57Y107_SLICE_X86Y107_B_XOR),
.I1(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I2(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I3(CLBLL_R_X57Y106_SLICE_X87Y106_B_XOR),
.I4(CLBLM_L_X62Y108_SLICE_X92Y108_BO5),
.I5(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.O5(CLBLL_R_X57Y108_SLICE_X87Y108_BO5),
.O6(CLBLL_R_X57Y108_SLICE_X87Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbabbbbbbaaaaaaa)
  ) CLBLL_R_X57Y108_SLICE_X87Y108_ALUT (
.I0(CLBLM_L_X62Y106_SLICE_X93Y106_BO5),
.I1(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I2(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I3(CLBLL_R_X57Y106_SLICE_X87Y106_A_XOR),
.I4(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I5(CLBLL_R_X57Y107_SLICE_X86Y107_A_XOR),
.O5(CLBLL_R_X57Y108_SLICE_X87Y108_AO5),
.O6(CLBLL_R_X57Y108_SLICE_X87Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X57Y109_SLICE_X86Y109_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y100_SLICE_X90Y100_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_R_X57Y109_SLICE_X86Y109_AO6),
.Q(CLBLL_R_X57Y109_SLICE_X86Y109_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X57Y109_SLICE_X86Y109_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y100_SLICE_X90Y100_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_R_X57Y109_SLICE_X86Y109_BO6),
.Q(CLBLL_R_X57Y109_SLICE_X86Y109_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X57Y109_SLICE_X86Y109_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y100_SLICE_X90Y100_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_R_X57Y109_SLICE_X86Y109_CO6),
.Q(CLBLL_R_X57Y109_SLICE_X86Y109_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2e2e2ff33cc00)
  ) CLBLL_R_X57Y109_SLICE_X86Y109_DLUT (
.I0(CLBLL_R_X57Y111_SLICE_X87Y111_C_XOR),
.I1(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I2(CLBLL_R_X57Y109_SLICE_X86Y109_BQ),
.I3(CLBLL_R_X57Y108_SLICE_X86Y108_B_XOR),
.I4(CLBLM_R_X59Y99_SLICE_X89Y99_BQ),
.I5(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.O5(CLBLL_R_X57Y109_SLICE_X86Y109_DO5),
.O6(CLBLL_R_X57Y109_SLICE_X86Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0aaccccaaaa)
  ) CLBLL_R_X57Y109_SLICE_X86Y109_CLUT (
.I0(CLBLL_R_X57Y108_SLICE_X86Y108_C_XOR),
.I1(CLBLM_L_X62Y100_SLICE_X93Y100_BO6),
.I2(CLBLL_R_X57Y107_SLICE_X87Y107_C_XOR),
.I3(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I4(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I5(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.O5(CLBLL_R_X57Y109_SLICE_X86Y109_CO5),
.O6(CLBLL_R_X57Y109_SLICE_X86Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafc0a0cfcfc0c0c)
  ) CLBLL_R_X57Y109_SLICE_X86Y109_BLUT (
.I0(CLBLL_R_X57Y107_SLICE_X87Y107_B_XOR),
.I1(CLBLL_R_X57Y108_SLICE_X86Y108_B_XOR),
.I2(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I3(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I4(CLBLM_L_X62Y100_SLICE_X93Y100_AO6),
.I5(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.O5(CLBLL_R_X57Y109_SLICE_X86Y109_BO5),
.O6(CLBLL_R_X57Y109_SLICE_X86Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefc0e0cf4fc040c)
  ) CLBLL_R_X57Y109_SLICE_X86Y109_ALUT (
.I0(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I1(CLBLL_R_X57Y108_SLICE_X86Y108_A_XOR),
.I2(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I3(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I4(CLBLM_L_X62Y97_SLICE_X92Y97_BO6),
.I5(CLBLL_R_X57Y107_SLICE_X87Y107_A_XOR),
.O5(CLBLL_R_X57Y109_SLICE_X86Y109_AO5),
.O6(CLBLL_R_X57Y109_SLICE_X86Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_R_X57Y109_SLICE_X87Y109_CARRY4 (
.CI(1'b0),
.CO({CLBLL_R_X57Y109_SLICE_X87Y109_D_CY, CLBLL_R_X57Y109_SLICE_X87Y109_C_CY, CLBLL_R_X57Y109_SLICE_X87Y109_B_CY, CLBLL_R_X57Y109_SLICE_X87Y109_A_CY}),
.CYINIT(1'b0),
.DI({CLBLL_R_X57Y105_SLICE_X86Y105_BQ, CLBLL_R_X57Y105_SLICE_X86Y105_AQ, CLBLM_R_X59Y106_SLICE_X88Y106_BQ, CLBLL_R_X57Y101_SLICE_X86Y101_AQ}),
.O({CLBLL_R_X57Y109_SLICE_X87Y109_D_XOR, CLBLL_R_X57Y109_SLICE_X87Y109_C_XOR, CLBLL_R_X57Y109_SLICE_X87Y109_B_XOR, CLBLL_R_X57Y109_SLICE_X87Y109_A_XOR}),
.S({CLBLL_R_X57Y109_SLICE_X87Y109_DO6, CLBLL_R_X57Y109_SLICE_X87Y109_CO6, CLBLL_R_X57Y109_SLICE_X87Y109_BO6, CLBLL_R_X57Y109_SLICE_X87Y109_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555555aaaaaaaa)
  ) CLBLL_R_X57Y109_SLICE_X87Y109_DLUT (
.I0(CLBLM_R_X59Y98_SLICE_X89Y98_B5Q),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_R_X57Y105_SLICE_X86Y105_BQ),
.O5(CLBLL_R_X57Y109_SLICE_X87Y109_DO5),
.O6(CLBLL_R_X57Y109_SLICE_X87Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555555aaaaaaaa)
  ) CLBLL_R_X57Y109_SLICE_X87Y109_CLUT (
.I0(CLBLM_R_X59Y98_SLICE_X89Y98_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_R_X57Y105_SLICE_X86Y105_AQ),
.O5(CLBLL_R_X57Y109_SLICE_X87Y109_CO5),
.O6(CLBLL_R_X57Y109_SLICE_X87Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3c3c3c3c3c)
  ) CLBLL_R_X57Y109_SLICE_X87Y109_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X59Y106_SLICE_X88Y106_BQ),
.I2(CLBLM_R_X59Y98_SLICE_X89Y98_A5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y109_SLICE_X87Y109_BO5),
.O6(CLBLL_R_X57Y109_SLICE_X87Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffffffff0000)
  ) CLBLL_R_X57Y109_SLICE_X87Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_R_X57Y101_SLICE_X86Y101_AQ),
.I5(CLBLM_R_X59Y98_SLICE_X89Y98_AQ),
.O5(CLBLL_R_X57Y109_SLICE_X87Y109_AO5),
.O6(CLBLL_R_X57Y109_SLICE_X87Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y110_SLICE_X86Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y110_SLICE_X86Y110_DO5),
.O6(CLBLL_R_X57Y110_SLICE_X86Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y110_SLICE_X86Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y110_SLICE_X86Y110_CO5),
.O6(CLBLL_R_X57Y110_SLICE_X86Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y110_SLICE_X86Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y110_SLICE_X86Y110_BO5),
.O6(CLBLL_R_X57Y110_SLICE_X86Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y110_SLICE_X86Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y110_SLICE_X86Y110_AO5),
.O6(CLBLL_R_X57Y110_SLICE_X86Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_R_X57Y110_SLICE_X87Y110_CARRY4 (
.CI(CLBLL_R_X57Y109_SLICE_X87Y109_COUT),
.CO({CLBLL_R_X57Y110_SLICE_X87Y110_D_CY, CLBLL_R_X57Y110_SLICE_X87Y110_C_CY, CLBLL_R_X57Y110_SLICE_X87Y110_B_CY, CLBLL_R_X57Y110_SLICE_X87Y110_A_CY}),
.CYINIT(1'b0),
.DI({CLBLM_R_X59Y106_SLICE_X88Y106_AQ, CLBLL_R_X57Y108_SLICE_X87Y108_BQ, CLBLL_R_X57Y108_SLICE_X87Y108_AQ, CLBLL_R_X57Y103_SLICE_X87Y103_AQ}),
.O({CLBLL_R_X57Y110_SLICE_X87Y110_D_XOR, CLBLL_R_X57Y110_SLICE_X87Y110_C_XOR, CLBLL_R_X57Y110_SLICE_X87Y110_B_XOR, CLBLL_R_X57Y110_SLICE_X87Y110_A_XOR}),
.S({CLBLL_R_X57Y110_SLICE_X87Y110_DO6, CLBLL_R_X57Y110_SLICE_X87Y110_CO6, CLBLL_R_X57Y110_SLICE_X87Y110_BO6, CLBLL_R_X57Y110_SLICE_X87Y110_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6666666666666666)
  ) CLBLL_R_X57Y110_SLICE_X87Y110_DLUT (
.I0(CLBLM_R_X59Y106_SLICE_X88Y106_AQ),
.I1(CLBLM_R_X59Y96_SLICE_X89Y96_A5Q),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y110_SLICE_X87Y110_DO5),
.O6(CLBLL_R_X57Y110_SLICE_X87Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6666666666666666)
  ) CLBLL_R_X57Y110_SLICE_X87Y110_CLUT (
.I0(CLBLL_R_X57Y108_SLICE_X87Y108_BQ),
.I1(CLBLM_R_X59Y96_SLICE_X89Y96_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y110_SLICE_X87Y110_CO5),
.O6(CLBLL_R_X57Y110_SLICE_X87Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3c3c3c3c3c)
  ) CLBLL_R_X57Y110_SLICE_X87Y110_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X59Y98_SLICE_X89Y98_C5Q),
.I2(CLBLL_R_X57Y108_SLICE_X87Y108_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y110_SLICE_X87Y110_BO5),
.O6(CLBLL_R_X57Y110_SLICE_X87Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0ff0f00f0ff0f0)
  ) CLBLL_R_X57Y110_SLICE_X87Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X59Y98_SLICE_X89Y98_CQ),
.I3(1'b1),
.I4(CLBLL_R_X57Y103_SLICE_X87Y103_AQ),
.I5(1'b1),
.O5(CLBLL_R_X57Y110_SLICE_X87Y110_AO5),
.O6(CLBLL_R_X57Y110_SLICE_X87Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y111_SLICE_X86Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y111_SLICE_X86Y111_DO5),
.O6(CLBLL_R_X57Y111_SLICE_X86Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y111_SLICE_X86Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y111_SLICE_X86Y111_CO5),
.O6(CLBLL_R_X57Y111_SLICE_X86Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y111_SLICE_X86Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y111_SLICE_X86Y111_BO5),
.O6(CLBLL_R_X57Y111_SLICE_X86Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y111_SLICE_X86Y111_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y111_SLICE_X86Y111_AO5),
.O6(CLBLL_R_X57Y111_SLICE_X86Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_R_X57Y111_SLICE_X87Y111_CARRY4 (
.CI(CLBLL_R_X57Y110_SLICE_X87Y110_COUT),
.CO({CLBLL_R_X57Y111_SLICE_X87Y111_D_CY, CLBLL_R_X57Y111_SLICE_X87Y111_C_CY, CLBLL_R_X57Y111_SLICE_X87Y111_B_CY, CLBLL_R_X57Y111_SLICE_X87Y111_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLL_R_X57Y111_SLICE_X87Y111_D_XOR, CLBLL_R_X57Y111_SLICE_X87Y111_C_XOR, CLBLL_R_X57Y111_SLICE_X87Y111_B_XOR, CLBLL_R_X57Y111_SLICE_X87Y111_A_XOR}),
.S({CLBLL_R_X57Y111_SLICE_X87Y111_DO6, CLBLL_R_X57Y111_SLICE_X87Y111_CO6, CLBLL_R_X57Y111_SLICE_X87Y111_BO6, CLBLL_R_X57Y111_SLICE_X87Y111_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLL_R_X57Y111_SLICE_X87Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_R_X57Y109_SLICE_X86Y109_CQ),
.O5(CLBLL_R_X57Y111_SLICE_X87Y111_DO5),
.O6(CLBLL_R_X57Y111_SLICE_X87Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLL_R_X57Y111_SLICE_X87Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_R_X57Y109_SLICE_X86Y109_BQ),
.O5(CLBLL_R_X57Y111_SLICE_X87Y111_CO5),
.O6(CLBLL_R_X57Y111_SLICE_X87Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLL_R_X57Y111_SLICE_X87Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_R_X57Y109_SLICE_X86Y109_AQ),
.O5(CLBLL_R_X57Y111_SLICE_X87Y111_BO5),
.O6(CLBLL_R_X57Y111_SLICE_X87Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLL_R_X57Y111_SLICE_X87Y111_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X60Y108_SLICE_X91Y108_AQ),
.O5(CLBLL_R_X57Y111_SLICE_X87Y111_AO5),
.O6(CLBLL_R_X57Y111_SLICE_X87Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X32Y119_SLICE_X46Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(CLBLM_R_X15Y122_SLICE_X20Y122_AO6),
.D(LIOB33_X0Y119_IOB_X0Y119_I),
.Q(CLBLM_L_X32Y119_SLICE_X46Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X32Y119_SLICE_X46Y119_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(CLBLM_R_X15Y122_SLICE_X20Y122_AO6),
.D(LIOB33_X0Y117_IOB_X0Y118_I),
.Q(CLBLM_L_X32Y119_SLICE_X46Y119_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X32Y119_SLICE_X46Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X32Y119_SLICE_X46Y119_DO5),
.O6(CLBLM_L_X32Y119_SLICE_X46Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X32Y119_SLICE_X46Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X32Y119_SLICE_X46Y119_CO5),
.O6(CLBLM_L_X32Y119_SLICE_X46Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X32Y119_SLICE_X46Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X32Y119_SLICE_X46Y119_BO5),
.O6(CLBLM_L_X32Y119_SLICE_X46Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X32Y119_SLICE_X46Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X32Y119_SLICE_X46Y119_AO5),
.O6(CLBLM_L_X32Y119_SLICE_X46Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X32Y119_SLICE_X47Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X32Y119_SLICE_X47Y119_DO5),
.O6(CLBLM_L_X32Y119_SLICE_X47Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X32Y119_SLICE_X47Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X32Y119_SLICE_X47Y119_CO5),
.O6(CLBLM_L_X32Y119_SLICE_X47Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X32Y119_SLICE_X47Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X32Y119_SLICE_X47Y119_BO5),
.O6(CLBLM_L_X32Y119_SLICE_X47Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X32Y119_SLICE_X47Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X32Y119_SLICE_X47Y119_AO5),
.O6(CLBLM_L_X32Y119_SLICE_X47Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X50Y104_SLICE_X76Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X56Y98_SLICE_X84Y98_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X50Y104_SLICE_X76Y104_AO6),
.Q(CLBLM_L_X50Y104_SLICE_X76Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555555333300ff)
  ) CLBLM_L_X50Y104_SLICE_X76Y104_DLUT (
.I0(CLBLL_R_X57Y100_SLICE_X86Y100_CQ),
.I1(CLBLL_R_X57Y97_SLICE_X86Y97_AQ),
.I2(1'b1),
.I3(CLBLL_R_X57Y99_SLICE_X86Y99_BQ),
.I4(CLBLM_R_X53Y101_SLICE_X80Y101_BQ),
.I5(CLBLL_L_X54Y100_SLICE_X82Y100_BQ),
.O5(CLBLM_L_X50Y104_SLICE_X76Y104_DO5),
.O6(CLBLM_L_X50Y104_SLICE_X76Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he6b3b380e6b3b380)
  ) CLBLM_L_X50Y104_SLICE_X76Y104_CLUT (
.I0(CLBLM_R_X53Y101_SLICE_X80Y101_BQ),
.I1(CLBLL_L_X54Y100_SLICE_X82Y100_BQ),
.I2(CLBLL_R_X57Y101_SLICE_X87Y101_CQ),
.I3(CLBLL_R_X57Y100_SLICE_X86Y100_DQ),
.I4(CLBLL_R_X57Y100_SLICE_X86Y100_AQ),
.I5(1'b1),
.O5(CLBLM_L_X50Y104_SLICE_X76Y104_CO5),
.O6(CLBLM_L_X50Y104_SLICE_X76Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55335f33aa33a033)
  ) CLBLM_L_X50Y104_SLICE_X76Y104_BLUT (
.I0(CLBLL_R_X57Y100_SLICE_X86Y100_AQ),
.I1(CLBLM_L_X50Y104_SLICE_X76Y104_DO6),
.I2(CLBLL_L_X54Y100_SLICE_X82Y100_BQ),
.I3(CLBLM_R_X53Y101_SLICE_X81Y101_AQ),
.I4(CLBLM_R_X53Y101_SLICE_X80Y101_BQ),
.I5(CLBLL_R_X57Y100_SLICE_X86Y100_DQ),
.O5(CLBLM_L_X50Y104_SLICE_X76Y104_BO5),
.O6(CLBLM_L_X50Y104_SLICE_X76Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hef23ef23ec20ec20)
  ) CLBLM_L_X50Y104_SLICE_X76Y104_ALUT (
.I0(CLBLM_L_X50Y107_SLICE_X76Y107_CO6),
.I1(CLBLM_R_X53Y100_SLICE_X81Y100_AQ),
.I2(CLBLM_R_X53Y101_SLICE_X81Y101_AQ),
.I3(CLBLM_L_X50Y104_SLICE_X76Y104_BO6),
.I4(1'b1),
.I5(CLBLM_L_X50Y104_SLICE_X76Y104_CO6),
.O5(CLBLM_L_X50Y104_SLICE_X76Y104_AO5),
.O6(CLBLM_L_X50Y104_SLICE_X76Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X50Y104_SLICE_X77Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X50Y104_SLICE_X77Y104_DO5),
.O6(CLBLM_L_X50Y104_SLICE_X77Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X50Y104_SLICE_X77Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X50Y104_SLICE_X77Y104_CO5),
.O6(CLBLM_L_X50Y104_SLICE_X77Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X50Y104_SLICE_X77Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X50Y104_SLICE_X77Y104_BO5),
.O6(CLBLM_L_X50Y104_SLICE_X77Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbbfebaebebbaba)
  ) CLBLM_L_X50Y104_SLICE_X77Y104_ALUT (
.I0(CLBLM_R_X53Y101_SLICE_X81Y101_AQ),
.I1(CLBLL_L_X54Y100_SLICE_X82Y100_BQ),
.I2(CLBLL_R_X57Y100_SLICE_X86Y100_BQ),
.I3(CLBLM_L_X56Y101_SLICE_X85Y101_DQ),
.I4(CLBLL_R_X57Y100_SLICE_X86Y100_CQ),
.I5(CLBLM_R_X53Y101_SLICE_X80Y101_BQ),
.O5(CLBLM_L_X50Y104_SLICE_X77Y104_AO5),
.O6(CLBLM_L_X50Y104_SLICE_X77Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X50Y105_SLICE_X76Y105_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X56Y98_SLICE_X84Y98_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X50Y105_SLICE_X76Y105_AO6),
.Q(CLBLM_L_X50Y105_SLICE_X76Y105_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X50Y105_SLICE_X76Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X50Y105_SLICE_X76Y105_DO5),
.O6(CLBLM_L_X50Y105_SLICE_X76Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff00000b03)
  ) CLBLM_L_X50Y105_SLICE_X76Y105_CLUT (
.I0(CLBLM_R_X53Y100_SLICE_X81Y100_AQ),
.I1(CLBLL_R_X57Y97_SLICE_X86Y97_AQ),
.I2(CLBLL_L_X52Y105_SLICE_X78Y105_AO6),
.I3(CLBLM_R_X53Y101_SLICE_X80Y101_BQ),
.I4(CLBLM_R_X53Y101_SLICE_X81Y101_AQ),
.I5(1'b1),
.O5(CLBLM_L_X50Y105_SLICE_X76Y105_CO5),
.O6(CLBLM_L_X50Y105_SLICE_X76Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55550f0f00cccccc)
  ) CLBLM_L_X50Y105_SLICE_X76Y105_BLUT (
.I0(CLBLL_R_X57Y99_SLICE_X86Y99_BQ),
.I1(CLBLM_R_X53Y100_SLICE_X81Y100_AQ),
.I2(CLBLM_L_X56Y101_SLICE_X85Y101_DQ),
.I3(CLBLL_R_X57Y97_SLICE_X86Y97_AQ),
.I4(CLBLL_L_X54Y100_SLICE_X82Y100_BQ),
.I5(1'b1),
.O5(CLBLM_L_X50Y105_SLICE_X76Y105_BO5),
.O6(CLBLM_L_X50Y105_SLICE_X76Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000dddc0000dddc)
  ) CLBLM_L_X50Y105_SLICE_X76Y105_ALUT (
.I0(CLBLM_L_X50Y105_SLICE_X76Y105_BO5),
.I1(CLBLL_L_X52Y105_SLICE_X78Y105_CO6),
.I2(CLBLM_L_X50Y111_SLICE_X76Y111_AO6),
.I3(CLBLM_L_X50Y111_SLICE_X76Y111_BO6),
.I4(CLBLM_L_X50Y105_SLICE_X76Y105_CO5),
.I5(1'b1),
.O5(CLBLM_L_X50Y105_SLICE_X76Y105_AO5),
.O6(CLBLM_L_X50Y105_SLICE_X76Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X50Y105_SLICE_X77Y105_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X56Y98_SLICE_X84Y98_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X50Y105_SLICE_X77Y105_F7AMUX_O),
.Q(CLBLM_L_X50Y105_SLICE_X77Y105_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbff008888ff00)
  ) CLBLM_L_X50Y105_SLICE_X77Y105_DLUT (
.I0(CLBLL_R_X57Y97_SLICE_X86Y97_AQ),
.I1(CLBLM_R_X53Y101_SLICE_X80Y101_BQ),
.I2(1'b1),
.I3(CLBLL_R_X57Y101_SLICE_X87Y101_DQ),
.I4(CLBLL_L_X54Y100_SLICE_X82Y100_BQ),
.I5(CLBLL_R_X57Y100_SLICE_X86Y100_DQ),
.O5(CLBLM_L_X50Y105_SLICE_X77Y105_DO5),
.O6(CLBLM_L_X50Y105_SLICE_X77Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h569a569a7b7b4848)
  ) CLBLM_L_X50Y105_SLICE_X77Y105_CLUT (
.I0(CLBLL_R_X57Y99_SLICE_X86Y99_BQ),
.I1(CLBLM_L_X50Y106_SLICE_X77Y106_AO5),
.I2(CLBLL_R_X57Y99_SLICE_X86Y99_AQ),
.I3(CLBLL_L_X52Y106_SLICE_X78Y106_AO5),
.I4(CLBLM_L_X50Y105_SLICE_X77Y105_DO6),
.I5(CLBLM_R_X49Y106_SLICE_X74Y106_CO6),
.O5(CLBLM_L_X50Y105_SLICE_X77Y105_CO5),
.O6(CLBLM_L_X50Y105_SLICE_X77Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0e0e0d0d0)
  ) CLBLM_L_X50Y105_SLICE_X77Y105_BLUT (
.I0(CLBLM_R_X49Y108_SLICE_X75Y108_B_XOR),
.I1(CLBLM_L_X50Y106_SLICE_X77Y106_AO6),
.I2(CLBLM_L_X50Y104_SLICE_X77Y104_AO6),
.I3(1'b1),
.I4(CLBLM_L_X50Y107_SLICE_X76Y107_AO6),
.I5(CLBLL_L_X54Y100_SLICE_X82Y100_BQ),
.O5(CLBLM_L_X50Y105_SLICE_X77Y105_BO5),
.O6(CLBLM_L_X50Y105_SLICE_X77Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fa55af01b1bb1b1)
  ) CLBLM_L_X50Y105_SLICE_X77Y105_ALUT (
.I0(CLBLM_R_X49Y106_SLICE_X74Y106_CO6),
.I1(CLBLL_L_X52Y105_SLICE_X78Y105_BO5),
.I2(CLBLL_R_X57Y100_SLICE_X86Y100_CQ),
.I3(CLBLL_R_X57Y100_SLICE_X86Y100_DQ),
.I4(CLBLL_R_X57Y100_SLICE_X86Y100_BQ),
.I5(CLBLM_L_X50Y106_SLICE_X77Y106_AO5),
.O5(CLBLM_L_X50Y105_SLICE_X77Y105_AO5),
.O6(CLBLM_L_X50Y105_SLICE_X77Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X50Y105_SLICE_X77Y105_MUXF7A (
.I0(CLBLM_L_X50Y105_SLICE_X77Y105_BO6),
.I1(CLBLM_L_X50Y105_SLICE_X77Y105_AO6),
.O(CLBLM_L_X50Y105_SLICE_X77Y105_F7AMUX_O),
.S(CLBLM_R_X53Y100_SLICE_X81Y100_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X50Y106_SLICE_X76Y106_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X56Y98_SLICE_X84Y98_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X50Y106_SLICE_X76Y106_AO6),
.Q(CLBLM_L_X50Y106_SLICE_X76Y106_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X50Y106_SLICE_X76Y106_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X56Y98_SLICE_X84Y98_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X50Y106_SLICE_X76Y106_CO6),
.Q(CLBLM_L_X50Y106_SLICE_X76Y106_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h03fc1dd1cf301dd1)
  ) CLBLM_L_X50Y106_SLICE_X76Y106_DLUT (
.I0(CLBLM_L_X50Y106_SLICE_X77Y106_BO6),
.I1(CLBLM_L_X50Y106_SLICE_X77Y106_AO5),
.I2(CLBLL_R_X57Y101_SLICE_X87Y101_AQ),
.I3(CLBLL_R_X57Y101_SLICE_X87Y101_CQ),
.I4(CLBLM_R_X49Y106_SLICE_X74Y106_CO6),
.I5(CLBLM_L_X50Y106_SLICE_X76Y106_BO6),
.O5(CLBLM_L_X50Y106_SLICE_X76Y106_DO5),
.O6(CLBLM_L_X50Y106_SLICE_X76Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0ffccccf000)
  ) CLBLM_L_X50Y106_SLICE_X76Y106_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X50Y106_SLICE_X77Y106_CO6),
.I2(CLBLM_R_X49Y108_SLICE_X74Y108_DO6),
.I3(CLBLM_R_X53Y101_SLICE_X81Y101_AQ),
.I4(CLBLM_R_X53Y100_SLICE_X81Y100_AQ),
.I5(CLBLL_L_X52Y107_SLICE_X78Y107_AO5),
.O5(CLBLM_L_X50Y106_SLICE_X76Y106_CO5),
.O6(CLBLM_L_X50Y106_SLICE_X76Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffcfffffffe)
  ) CLBLM_L_X50Y106_SLICE_X76Y106_BLUT (
.I0(CLBLL_R_X57Y101_SLICE_X87Y101_CQ),
.I1(CLBLL_R_X57Y100_SLICE_X86Y100_CQ),
.I2(CLBLL_R_X57Y100_SLICE_X86Y100_DQ),
.I3(CLBLL_R_X57Y100_SLICE_X87Y100_CQ),
.I4(CLBLM_L_X56Y101_SLICE_X85Y101_CQ),
.I5(1'b1),
.O5(CLBLM_L_X50Y106_SLICE_X76Y106_BO5),
.O6(CLBLM_L_X50Y106_SLICE_X76Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaccccaaaaff00)
  ) CLBLM_L_X50Y106_SLICE_X76Y106_ALUT (
.I0(CLBLM_L_X50Y106_SLICE_X76Y106_DO6),
.I1(CLBLM_R_X49Y107_SLICE_X74Y107_BO6),
.I2(1'b1),
.I3(CLBLL_L_X52Y106_SLICE_X79Y106_AO5),
.I4(CLBLM_R_X53Y100_SLICE_X81Y100_AQ),
.I5(CLBLM_R_X53Y101_SLICE_X81Y101_AQ),
.O5(CLBLM_L_X50Y106_SLICE_X76Y106_AO5),
.O6(CLBLM_L_X50Y106_SLICE_X76Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X50Y106_SLICE_X77Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X50Y106_SLICE_X77Y106_DO5),
.O6(CLBLM_L_X50Y106_SLICE_X77Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1d771d44e2bbe288)
  ) CLBLM_L_X50Y106_SLICE_X77Y106_CLUT (
.I0(CLBLM_L_X56Y101_SLICE_X85Y101_BQ),
.I1(CLBLM_R_X49Y106_SLICE_X74Y106_CO6),
.I2(CLBLM_L_X50Y106_SLICE_X76Y106_BO5),
.I3(CLBLM_L_X50Y106_SLICE_X77Y106_AO5),
.I4(CLBLM_L_X50Y106_SLICE_X77Y106_BO5),
.I5(CLBLM_L_X56Y101_SLICE_X85Y101_DQ),
.O5(CLBLM_L_X50Y106_SLICE_X77Y106_CO5),
.O6(CLBLM_L_X50Y106_SLICE_X77Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000ff0ffcacacaca)
  ) CLBLM_L_X50Y106_SLICE_X77Y106_BLUT (
.I0(CLBLL_R_X57Y101_SLICE_X87Y101_CQ),
.I1(CLBLL_R_X57Y101_SLICE_X87Y101_DQ),
.I2(CLBLL_L_X54Y100_SLICE_X82Y100_BQ),
.I3(CLBLL_R_X57Y100_SLICE_X87Y100_CQ),
.I4(CLBLM_L_X56Y101_SLICE_X85Y101_DQ),
.I5(1'b1),
.O5(CLBLM_L_X50Y106_SLICE_X77Y106_BO5),
.O6(CLBLM_L_X50Y106_SLICE_X77Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hef0f4f0ff050f050)
  ) CLBLM_L_X50Y106_SLICE_X77Y106_ALUT (
.I0(CLBLM_R_X53Y101_SLICE_X80Y101_BQ),
.I1(CLBLM_L_X50Y108_SLICE_X76Y108_B_XOR),
.I2(CLBLM_R_X53Y101_SLICE_X81Y101_AQ),
.I3(CLBLL_L_X54Y100_SLICE_X82Y100_BQ),
.I4(CLBLM_L_X50Y108_SLICE_X77Y108_B_XOR),
.I5(1'b1),
.O5(CLBLM_L_X50Y106_SLICE_X77Y106_AO5),
.O6(CLBLM_L_X50Y106_SLICE_X77Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X50Y107_SLICE_X76Y107_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X56Y98_SLICE_X84Y98_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X50Y107_SLICE_X76Y107_BO6),
.Q(CLBLM_L_X50Y107_SLICE_X76Y107_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf606fc0cfc0cfc0c)
  ) CLBLM_L_X50Y107_SLICE_X76Y107_DLUT (
.I0(CLBLM_R_X49Y109_SLICE_X75Y109_C_XOR),
.I1(CLBLM_R_X49Y109_SLICE_X75Y109_D_XOR),
.I2(CLBLL_L_X54Y100_SLICE_X82Y100_BQ),
.I3(CLBLM_L_X50Y107_SLICE_X76Y107_AO5),
.I4(CLBLM_R_X49Y109_SLICE_X75Y109_B_XOR),
.I5(CLBLM_R_X49Y107_SLICE_X74Y107_DO6),
.O5(CLBLM_L_X50Y107_SLICE_X76Y107_DO5),
.O6(CLBLM_L_X50Y107_SLICE_X76Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haffa0550dd88dd88)
  ) CLBLM_L_X50Y107_SLICE_X76Y107_CLUT (
.I0(CLBLL_L_X54Y100_SLICE_X82Y100_BQ),
.I1(CLBLM_L_X50Y108_SLICE_X76Y108_A_XOR),
.I2(CLBLL_R_X57Y97_SLICE_X86Y97_AQ),
.I3(CLBLM_R_X49Y108_SLICE_X75Y108_A_XOR),
.I4(CLBLM_L_X50Y108_SLICE_X77Y108_A_XOR),
.I5(CLBLM_R_X53Y101_SLICE_X80Y101_BQ),
.O5(CLBLM_L_X50Y107_SLICE_X76Y107_CO5),
.O6(CLBLM_L_X50Y107_SLICE_X76Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff3c00000f3c0)
  ) CLBLM_L_X50Y107_SLICE_X76Y107_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X53Y101_SLICE_X81Y101_AQ),
.I2(CLBLM_L_X50Y111_SLICE_X76Y111_CO6),
.I3(CLBLL_L_X52Y107_SLICE_X78Y107_BO5),
.I4(CLBLM_R_X53Y100_SLICE_X81Y100_AQ),
.I5(CLBLM_R_X49Y106_SLICE_X75Y106_CO6),
.O5(CLBLM_L_X50Y107_SLICE_X76Y107_BO5),
.O6(CLBLM_L_X50Y107_SLICE_X76Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5fffffccccff00)
  ) CLBLM_L_X50Y107_SLICE_X76Y107_ALUT (
.I0(CLBLL_R_X57Y97_SLICE_X86Y97_AQ),
.I1(CLBLM_L_X50Y109_SLICE_X77Y109_D_XOR),
.I2(CLBLM_R_X49Y108_SLICE_X75Y108_A_XOR),
.I3(CLBLM_L_X50Y109_SLICE_X76Y109_D_XOR),
.I4(CLBLM_R_X53Y101_SLICE_X80Y101_BQ),
.I5(1'b1),
.O5(CLBLM_L_X50Y107_SLICE_X76Y107_AO5),
.O6(CLBLM_L_X50Y107_SLICE_X76Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X50Y107_SLICE_X77Y107_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X56Y98_SLICE_X84Y98_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X50Y107_SLICE_X77Y107_AO6),
.Q(CLBLM_L_X50Y107_SLICE_X77Y107_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X50Y107_SLICE_X77Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X50Y107_SLICE_X77Y107_DO5),
.O6(CLBLM_L_X50Y107_SLICE_X77Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X50Y107_SLICE_X77Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X50Y107_SLICE_X77Y107_CO5),
.O6(CLBLM_L_X50Y107_SLICE_X77Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fc3c3fc0c0c0c)
  ) CLBLM_L_X50Y107_SLICE_X77Y107_BLUT (
.I0(1'b1),
.I1(CLBLL_R_X57Y99_SLICE_X86Y99_AQ),
.I2(CLBLL_L_X54Y100_SLICE_X82Y100_BQ),
.I3(CLBLL_R_X57Y100_SLICE_X87Y100_CQ),
.I4(CLBLM_R_X53Y101_SLICE_X80Y101_BQ),
.I5(CLBLL_R_X57Y99_SLICE_X86Y99_BQ),
.O5(CLBLM_L_X50Y107_SLICE_X77Y107_BO5),
.O6(CLBLM_L_X50Y107_SLICE_X77Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0cfc0cfc0)
  ) CLBLM_L_X50Y107_SLICE_X77Y107_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X50Y105_SLICE_X77Y105_CO6),
.I2(CLBLM_R_X53Y100_SLICE_X81Y100_AQ),
.I3(CLBLM_L_X50Y107_SLICE_X77Y107_BO6),
.I4(CLBLM_L_X50Y107_SLICE_X76Y107_DO6),
.I5(CLBLM_R_X53Y101_SLICE_X81Y101_AQ),
.O5(CLBLM_L_X50Y107_SLICE_X77Y107_AO5),
.O6(CLBLM_L_X50Y107_SLICE_X77Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X50Y108_SLICE_X76Y108_CARRY4 (
.CI(1'b0),
.CO({CLBLM_L_X50Y108_SLICE_X76Y108_D_CY, CLBLM_L_X50Y108_SLICE_X76Y108_C_CY, CLBLM_L_X50Y108_SLICE_X76Y108_B_CY, CLBLM_L_X50Y108_SLICE_X76Y108_A_CY}),
.CYINIT(1'b1),
.DI({CLBLL_R_X57Y100_SLICE_X87Y100_CQ, CLBLM_L_X56Y101_SLICE_X85Y101_CQ, CLBLL_R_X57Y100_SLICE_X86Y100_CQ, CLBLL_R_X57Y100_SLICE_X86Y100_DQ}),
.O({CLBLM_L_X50Y108_SLICE_X76Y108_D_XOR, CLBLM_L_X50Y108_SLICE_X76Y108_C_XOR, CLBLM_L_X50Y108_SLICE_X76Y108_B_XOR, CLBLM_L_X50Y108_SLICE_X76Y108_A_XOR}),
.S({CLBLM_L_X50Y108_SLICE_X76Y108_DO6, CLBLM_L_X50Y108_SLICE_X76Y108_CO6, CLBLM_L_X50Y108_SLICE_X76Y108_BO6, CLBLM_L_X50Y108_SLICE_X76Y108_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a5a5a5a5a5a5a5)
  ) CLBLM_L_X50Y108_SLICE_X76Y108_DLUT (
.I0(CLBLL_R_X57Y100_SLICE_X87Y100_AQ),
.I1(1'b1),
.I2(CLBLL_R_X57Y100_SLICE_X87Y100_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X50Y108_SLICE_X76Y108_DO5),
.O6(CLBLM_L_X50Y108_SLICE_X76Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a5a5a5a5a5a5a5)
  ) CLBLM_L_X50Y108_SLICE_X76Y108_CLUT (
.I0(CLBLM_L_X56Y101_SLICE_X85Y101_AQ),
.I1(1'b1),
.I2(CLBLM_L_X56Y101_SLICE_X85Y101_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X50Y108_SLICE_X76Y108_CO5),
.O6(CLBLM_L_X50Y108_SLICE_X76Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc3333cccc3333)
  ) CLBLM_L_X50Y108_SLICE_X76Y108_BLUT (
.I0(1'b1),
.I1(CLBLL_R_X57Y100_SLICE_X86Y100_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_R_X57Y100_SLICE_X86Y100_BQ),
.I5(1'b1),
.O5(CLBLM_L_X50Y108_SLICE_X76Y108_BO5),
.O6(CLBLM_L_X50Y108_SLICE_X76Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf00ff00ff00ff00f)
  ) CLBLM_L_X50Y108_SLICE_X76Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_R_X57Y100_SLICE_X86Y100_DQ),
.I3(CLBLL_R_X57Y100_SLICE_X86Y100_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X50Y108_SLICE_X76Y108_AO5),
.O6(CLBLM_L_X50Y108_SLICE_X76Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X50Y108_SLICE_X77Y108_CARRY4 (
.CI(1'b0),
.CO({CLBLM_L_X50Y108_SLICE_X77Y108_D_CY, CLBLM_L_X50Y108_SLICE_X77Y108_C_CY, CLBLM_L_X50Y108_SLICE_X77Y108_B_CY, CLBLM_L_X50Y108_SLICE_X77Y108_A_CY}),
.CYINIT(1'b1),
.DI({CLBLM_L_X50Y108_SLICE_X77Y108_DO5, CLBLM_L_X50Y108_SLICE_X77Y108_CO5, CLBLM_L_X50Y108_SLICE_X77Y108_BO5, 1'b1}),
.O({CLBLM_L_X50Y108_SLICE_X77Y108_D_XOR, CLBLM_L_X50Y108_SLICE_X77Y108_C_XOR, CLBLM_L_X50Y108_SLICE_X77Y108_B_XOR, CLBLM_L_X50Y108_SLICE_X77Y108_A_XOR}),
.S({CLBLM_L_X50Y108_SLICE_X77Y108_DO6, CLBLM_L_X50Y108_SLICE_X77Y108_CO6, CLBLM_L_X50Y108_SLICE_X77Y108_BO6, CLBLM_L_X50Y108_SLICE_X77Y108_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5f05a0f55005500)
  ) CLBLM_L_X50Y108_SLICE_X77Y108_DLUT (
.I0(CLBLM_L_X56Y101_SLICE_X85Y101_AQ),
.I1(1'b1),
.I2(CLBLL_R_X57Y100_SLICE_X87Y100_AQ),
.I3(CLBLM_L_X56Y101_SLICE_X85Y101_CQ),
.I4(CLBLL_R_X57Y100_SLICE_X87Y100_CQ),
.I5(1'b1),
.O5(CLBLM_L_X50Y108_SLICE_X77Y108_DO5),
.O6(CLBLM_L_X50Y108_SLICE_X77Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a569690000cccc)
  ) CLBLM_L_X50Y108_SLICE_X77Y108_CLUT (
.I0(CLBLM_L_X56Y101_SLICE_X85Y101_AQ),
.I1(CLBLL_R_X57Y100_SLICE_X86Y100_CQ),
.I2(CLBLM_L_X56Y101_SLICE_X85Y101_CQ),
.I3(1'b1),
.I4(CLBLL_R_X57Y100_SLICE_X86Y100_BQ),
.I5(1'b1),
.O5(CLBLM_L_X50Y108_SLICE_X77Y108_CO5),
.O6(CLBLM_L_X50Y108_SLICE_X77Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4bb4d22dbbbb2222)
  ) CLBLM_L_X50Y108_SLICE_X77Y108_BLUT (
.I0(CLBLL_R_X57Y97_SLICE_X86Y97_AQ),
.I1(CLBLL_R_X57Y100_SLICE_X86Y100_AQ),
.I2(CLBLL_R_X57Y100_SLICE_X86Y100_BQ),
.I3(CLBLL_R_X57Y100_SLICE_X86Y100_CQ),
.I4(CLBLL_R_X57Y100_SLICE_X86Y100_DQ),
.I5(1'b1),
.O5(CLBLM_L_X50Y108_SLICE_X77Y108_BO5),
.O6(CLBLM_L_X50Y108_SLICE_X77Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf00f0ff0f00f0ff0)
  ) CLBLM_L_X50Y108_SLICE_X77Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_R_X57Y97_SLICE_X86Y97_AQ),
.I3(CLBLL_R_X57Y100_SLICE_X86Y100_AQ),
.I4(CLBLL_R_X57Y100_SLICE_X86Y100_DQ),
.I5(1'b1),
.O5(CLBLM_L_X50Y108_SLICE_X77Y108_AO5),
.O6(CLBLM_L_X50Y108_SLICE_X77Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X50Y109_SLICE_X76Y109_CARRY4 (
.CI(CLBLM_L_X50Y108_SLICE_X76Y108_COUT),
.CO({CLBLM_L_X50Y109_SLICE_X76Y109_D_CY, CLBLM_L_X50Y109_SLICE_X76Y109_C_CY, CLBLM_L_X50Y109_SLICE_X76Y109_B_CY, CLBLM_L_X50Y109_SLICE_X76Y109_A_CY}),
.CYINIT(1'b0),
.DI({CLBLL_R_X57Y99_SLICE_X86Y99_BQ, CLBLL_R_X57Y101_SLICE_X87Y101_DQ, CLBLM_L_X56Y101_SLICE_X85Y101_DQ, CLBLL_R_X57Y101_SLICE_X87Y101_CQ}),
.O({CLBLM_L_X50Y109_SLICE_X76Y109_D_XOR, CLBLM_L_X50Y109_SLICE_X76Y109_C_XOR, CLBLM_L_X50Y109_SLICE_X76Y109_B_XOR, CLBLM_L_X50Y109_SLICE_X76Y109_A_XOR}),
.S({CLBLM_L_X50Y109_SLICE_X76Y109_DO6, CLBLM_L_X50Y109_SLICE_X76Y109_CO6, CLBLM_L_X50Y109_SLICE_X76Y109_BO6, CLBLM_L_X50Y109_SLICE_X76Y109_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0000ff00ff)
  ) CLBLM_L_X50Y109_SLICE_X76Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_R_X57Y99_SLICE_X86Y99_BQ),
.I4(1'b1),
.I5(CLBLL_R_X57Y99_SLICE_X86Y99_AQ),
.O5(CLBLM_L_X50Y109_SLICE_X76Y109_DO5),
.O6(CLBLM_L_X50Y109_SLICE_X76Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a5a5a5a5a5a5a5)
  ) CLBLM_L_X50Y109_SLICE_X76Y109_CLUT (
.I0(CLBLL_R_X57Y100_SLICE_X87Y100_BQ),
.I1(1'b1),
.I2(CLBLL_R_X57Y101_SLICE_X87Y101_DQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X50Y109_SLICE_X76Y109_CO5),
.O6(CLBLM_L_X50Y109_SLICE_X76Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00f0ff0f00f0f)
  ) CLBLM_L_X50Y109_SLICE_X76Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X56Y101_SLICE_X85Y101_BQ),
.I3(1'b1),
.I4(CLBLM_L_X56Y101_SLICE_X85Y101_DQ),
.I5(1'b1),
.O5(CLBLM_L_X50Y109_SLICE_X76Y109_BO5),
.O6(CLBLM_L_X50Y109_SLICE_X76Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc33cc33cc33cc33)
  ) CLBLM_L_X50Y109_SLICE_X76Y109_ALUT (
.I0(1'b1),
.I1(CLBLL_R_X57Y101_SLICE_X87Y101_CQ),
.I2(1'b1),
.I3(CLBLL_R_X57Y101_SLICE_X87Y101_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X50Y109_SLICE_X76Y109_AO5),
.O6(CLBLM_L_X50Y109_SLICE_X76Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X50Y109_SLICE_X77Y109_CARRY4 (
.CI(CLBLM_L_X50Y108_SLICE_X77Y108_COUT),
.CO({CLBLM_L_X50Y109_SLICE_X77Y109_D_CY, CLBLM_L_X50Y109_SLICE_X77Y109_C_CY, CLBLM_L_X50Y109_SLICE_X77Y109_B_CY, CLBLM_L_X50Y109_SLICE_X77Y109_A_CY}),
.CYINIT(1'b0),
.DI({CLBLM_L_X50Y109_SLICE_X77Y109_DO5, CLBLM_L_X50Y109_SLICE_X77Y109_CO5, CLBLM_L_X50Y109_SLICE_X77Y109_BO5, CLBLM_L_X50Y109_SLICE_X77Y109_AO5}),
.O({CLBLM_L_X50Y109_SLICE_X77Y109_D_XOR, CLBLM_L_X50Y109_SLICE_X77Y109_C_XOR, CLBLM_L_X50Y109_SLICE_X77Y109_B_XOR, CLBLM_L_X50Y109_SLICE_X77Y109_A_XOR}),
.S({CLBLM_L_X50Y109_SLICE_X77Y109_DO6, CLBLM_L_X50Y109_SLICE_X77Y109_CO6, CLBLM_L_X50Y109_SLICE_X77Y109_BO6, CLBLM_L_X50Y109_SLICE_X77Y109_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9966cc3355550000)
  ) CLBLM_L_X50Y109_SLICE_X77Y109_DLUT (
.I0(CLBLL_R_X57Y100_SLICE_X87Y100_BQ),
.I1(CLBLL_R_X57Y99_SLICE_X86Y99_AQ),
.I2(1'b1),
.I3(CLBLL_R_X57Y99_SLICE_X86Y99_BQ),
.I4(CLBLL_R_X57Y101_SLICE_X87Y101_DQ),
.I5(1'b1),
.O5(CLBLM_L_X50Y109_SLICE_X77Y109_DO5),
.O6(CLBLM_L_X50Y109_SLICE_X77Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9696a5a533330000)
  ) CLBLM_L_X50Y109_SLICE_X77Y109_CLUT (
.I0(CLBLL_R_X57Y100_SLICE_X87Y100_BQ),
.I1(CLBLM_L_X56Y101_SLICE_X85Y101_BQ),
.I2(CLBLL_R_X57Y101_SLICE_X87Y101_DQ),
.I3(1'b1),
.I4(CLBLM_L_X56Y101_SLICE_X85Y101_DQ),
.I5(1'b1),
.O5(CLBLM_L_X50Y109_SLICE_X77Y109_CO5),
.O6(CLBLM_L_X50Y109_SLICE_X77Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc33cf00f33330000)
  ) CLBLM_L_X50Y109_SLICE_X77Y109_BLUT (
.I0(1'b1),
.I1(CLBLL_R_X57Y101_SLICE_X87Y101_AQ),
.I2(CLBLM_L_X56Y101_SLICE_X85Y101_BQ),
.I3(CLBLM_L_X56Y101_SLICE_X85Y101_DQ),
.I4(CLBLL_R_X57Y101_SLICE_X87Y101_CQ),
.I5(1'b1),
.O5(CLBLM_L_X50Y109_SLICE_X77Y109_BO5),
.O6(CLBLM_L_X50Y109_SLICE_X77Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc33ccc330f0f0000)
  ) CLBLM_L_X50Y109_SLICE_X77Y109_ALUT (
.I0(1'b1),
.I1(CLBLL_R_X57Y101_SLICE_X87Y101_AQ),
.I2(CLBLL_R_X57Y100_SLICE_X87Y100_AQ),
.I3(CLBLL_R_X57Y101_SLICE_X87Y101_CQ),
.I4(CLBLL_R_X57Y100_SLICE_X87Y100_CQ),
.I5(1'b1),
.O5(CLBLM_L_X50Y109_SLICE_X77Y109_AO5),
.O6(CLBLM_L_X50Y109_SLICE_X77Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X50Y110_SLICE_X76Y110_CARRY4 (
.CI(CLBLM_L_X50Y109_SLICE_X76Y109_COUT),
.CO({CLBLM_L_X50Y110_SLICE_X76Y110_D_CY, CLBLM_L_X50Y110_SLICE_X76Y110_C_CY, CLBLM_L_X50Y110_SLICE_X76Y110_B_CY, CLBLM_L_X50Y110_SLICE_X76Y110_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_L_X50Y110_SLICE_X76Y110_D_XOR, CLBLM_L_X50Y110_SLICE_X76Y110_C_XOR, CLBLM_L_X50Y110_SLICE_X76Y110_B_XOR, CLBLM_L_X50Y110_SLICE_X76Y110_A_XOR}),
.S({CLBLM_L_X50Y110_SLICE_X76Y110_DO6, CLBLM_L_X50Y110_SLICE_X76Y110_CO6, CLBLM_L_X50Y110_SLICE_X76Y110_BO6, CLBLM_L_X50Y110_SLICE_X76Y110_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X50Y110_SLICE_X76Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X50Y110_SLICE_X76Y110_DO5),
.O6(CLBLM_L_X50Y110_SLICE_X76Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X50Y110_SLICE_X76Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X50Y110_SLICE_X76Y110_CO5),
.O6(CLBLM_L_X50Y110_SLICE_X76Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X50Y110_SLICE_X76Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X50Y110_SLICE_X76Y110_BO5),
.O6(CLBLM_L_X50Y110_SLICE_X76Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffff)
  ) CLBLM_L_X50Y110_SLICE_X76Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X50Y110_SLICE_X76Y110_AO5),
.O6(CLBLM_L_X50Y110_SLICE_X76Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X50Y110_SLICE_X77Y110_CARRY4 (
.CI(CLBLM_L_X50Y109_SLICE_X77Y109_COUT),
.CO({CLBLM_L_X50Y110_SLICE_X77Y110_D_CY, CLBLM_L_X50Y110_SLICE_X77Y110_C_CY, CLBLM_L_X50Y110_SLICE_X77Y110_B_CY, CLBLM_L_X50Y110_SLICE_X77Y110_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_L_X50Y110_SLICE_X77Y110_D_XOR, CLBLM_L_X50Y110_SLICE_X77Y110_C_XOR, CLBLM_L_X50Y110_SLICE_X77Y110_B_XOR, CLBLM_L_X50Y110_SLICE_X77Y110_A_XOR}),
.S({CLBLM_L_X50Y110_SLICE_X77Y110_DO6, CLBLM_L_X50Y110_SLICE_X77Y110_CO6, CLBLM_L_X50Y110_SLICE_X77Y110_BO6, CLBLM_L_X50Y110_SLICE_X77Y110_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X50Y110_SLICE_X77Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X50Y110_SLICE_X77Y110_DO5),
.O6(CLBLM_L_X50Y110_SLICE_X77Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X50Y110_SLICE_X77Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X50Y110_SLICE_X77Y110_CO5),
.O6(CLBLM_L_X50Y110_SLICE_X77Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X50Y110_SLICE_X77Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X50Y110_SLICE_X77Y110_BO5),
.O6(CLBLM_L_X50Y110_SLICE_X77Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ffffff00ffff)
  ) CLBLM_L_X50Y110_SLICE_X77Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_R_X57Y99_SLICE_X86Y99_AQ),
.I4(CLBLL_R_X57Y99_SLICE_X86Y99_BQ),
.I5(1'b1),
.O5(CLBLM_L_X50Y110_SLICE_X77Y110_AO5),
.O6(CLBLM_L_X50Y110_SLICE_X77Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaacccccccc)
  ) CLBLM_L_X50Y111_SLICE_X76Y111_DLUT (
.I0(CLBLM_L_X50Y109_SLICE_X77Y109_C_XOR),
.I1(CLBLM_L_X50Y109_SLICE_X76Y109_C_XOR),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X53Y101_SLICE_X80Y101_BQ),
.O5(CLBLM_L_X50Y111_SLICE_X76Y111_DO5),
.O6(CLBLM_L_X50Y111_SLICE_X76Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff780078ff780078)
  ) CLBLM_L_X50Y111_SLICE_X76Y111_CLUT (
.I0(CLBLM_R_X49Y109_SLICE_X75Y109_B_XOR),
.I1(CLBLM_R_X49Y107_SLICE_X74Y107_DO6),
.I2(CLBLM_R_X49Y109_SLICE_X75Y109_C_XOR),
.I3(CLBLL_L_X54Y100_SLICE_X82Y100_BQ),
.I4(CLBLM_L_X50Y111_SLICE_X76Y111_DO6),
.I5(1'b1),
.O5(CLBLM_L_X50Y111_SLICE_X76Y111_CO5),
.O6(CLBLM_L_X50Y111_SLICE_X76Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff333f00ff330c00)
  ) CLBLM_L_X50Y111_SLICE_X76Y111_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X53Y101_SLICE_X80Y101_BQ),
.I2(CLBLM_L_X50Y110_SLICE_X77Y110_A_XOR),
.I3(CLBLL_L_X54Y100_SLICE_X82Y100_BQ),
.I4(CLBLM_R_X53Y100_SLICE_X81Y100_AQ),
.I5(CLBLM_L_X50Y110_SLICE_X76Y110_A_CY),
.O5(CLBLM_L_X50Y111_SLICE_X76Y111_BO5),
.O6(CLBLM_L_X50Y111_SLICE_X76Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000007fff8000)
  ) CLBLM_L_X50Y111_SLICE_X76Y111_ALUT (
.I0(CLBLM_R_X49Y107_SLICE_X74Y107_DO6),
.I1(CLBLM_R_X49Y109_SLICE_X75Y109_C_XOR),
.I2(CLBLM_R_X49Y109_SLICE_X75Y109_B_XOR),
.I3(CLBLM_R_X49Y109_SLICE_X75Y109_D_XOR),
.I4(CLBLM_R_X49Y110_SLICE_X75Y110_A_CY),
.I5(CLBLL_L_X54Y100_SLICE_X82Y100_BQ),
.O5(CLBLM_L_X50Y111_SLICE_X76Y111_AO5),
.O6(CLBLM_L_X50Y111_SLICE_X76Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X50Y111_SLICE_X77Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X50Y111_SLICE_X77Y111_DO5),
.O6(CLBLM_L_X50Y111_SLICE_X77Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X50Y111_SLICE_X77Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X50Y111_SLICE_X77Y111_CO5),
.O6(CLBLM_L_X50Y111_SLICE_X77Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X50Y111_SLICE_X77Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X50Y111_SLICE_X77Y111_BO5),
.O6(CLBLM_L_X50Y111_SLICE_X77Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X50Y111_SLICE_X77Y111_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X50Y111_SLICE_X77Y111_AO5),
.O6(CLBLM_L_X50Y111_SLICE_X77Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y97_SLICE_X84Y97_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y97_SLICE_X84Y97_BO6),
.Q(CLBLM_L_X56Y97_SLICE_X84Y97_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y97_SLICE_X84Y97_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y97_SLICE_X84Y97_DO6),
.Q(CLBLM_L_X56Y97_SLICE_X84Y97_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaffaaffeaffaa)
  ) CLBLM_L_X56Y97_SLICE_X84Y97_DLUT (
.I0(CLBLM_L_X56Y98_SLICE_X84Y98_CO6),
.I1(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.I2(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.I3(CLBLM_L_X56Y97_SLICE_X84Y97_AO5),
.I4(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I5(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.O5(CLBLM_L_X56Y97_SLICE_X84Y97_DO5),
.O6(CLBLM_L_X56Y97_SLICE_X84Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0008000000000101)
  ) CLBLM_L_X56Y97_SLICE_X84Y97_CLUT (
.I0(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.I1(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.I2(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.I3(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I4(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I5(1'b1),
.O5(CLBLM_L_X56Y97_SLICE_X84Y97_CO5),
.O6(CLBLM_L_X56Y97_SLICE_X84Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff80ccffffc0cc)
  ) CLBLM_L_X56Y97_SLICE_X84Y97_BLUT (
.I0(CLBLM_R_X49Y108_SLICE_X75Y108_DQ),
.I1(CLBLM_L_X56Y97_SLICE_X85Y97_BO5),
.I2(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.I3(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I4(CLBLM_L_X56Y98_SLICE_X84Y98_CO6),
.I5(CLBLM_R_X49Y107_SLICE_X75Y107_DQ),
.O5(CLBLM_L_X56Y97_SLICE_X84Y97_BO5),
.O6(CLBLM_L_X56Y97_SLICE_X84Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000f00080ccc0cc)
  ) CLBLM_L_X56Y97_SLICE_X84Y97_ALUT (
.I0(CLBLM_R_X49Y108_SLICE_X75Y108_DQ),
.I1(CLBLM_L_X56Y97_SLICE_X85Y97_BO5),
.I2(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.I3(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I4(CLBLM_R_X49Y107_SLICE_X75Y107_DQ),
.I5(1'b1),
.O5(CLBLM_L_X56Y97_SLICE_X84Y97_AO5),
.O6(CLBLM_L_X56Y97_SLICE_X84Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y97_SLICE_X85Y97_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y97_SLICE_X85Y97_AO6),
.Q(CLBLM_L_X56Y97_SLICE_X85Y97_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y97_SLICE_X85Y97_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y97_SLICE_X85Y97_CO6),
.Q(CLBLM_L_X56Y97_SLICE_X85Y97_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c088bb3333cc00)
  ) CLBLM_L_X56Y97_SLICE_X85Y97_DLUT (
.I0(CLBLM_L_X50Y105_SLICE_X76Y105_AQ),
.I1(CLBLM_L_X56Y97_SLICE_X85Y97_CQ),
.I2(CLBLM_L_X60Y98_SLICE_X90Y98_AQ),
.I3(CLBLM_L_X60Y97_SLICE_X90Y97_BO6),
.I4(CLBLM_L_X56Y97_SLICE_X84Y97_DQ),
.I5(CLBLL_L_X54Y98_SLICE_X83Y98_AQ),
.O5(CLBLM_L_X56Y97_SLICE_X85Y97_DO5),
.O6(CLBLM_L_X56Y97_SLICE_X85Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h020204040a0a0008)
  ) CLBLM_L_X56Y97_SLICE_X85Y97_CLUT (
.I0(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.I1(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.I2(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.I3(CLBLM_R_X49Y107_SLICE_X75Y107_DQ),
.I4(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I5(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.O5(CLBLM_L_X56Y97_SLICE_X85Y97_CO5),
.O6(CLBLM_L_X56Y97_SLICE_X85Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2200000044000000)
  ) CLBLM_L_X56Y97_SLICE_X85Y97_BLUT (
.I0(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.I1(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.I2(1'b1),
.I3(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.I4(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I5(1'b1),
.O5(CLBLM_L_X56Y97_SLICE_X85Y97_BO5),
.O6(CLBLM_L_X56Y97_SLICE_X85Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa2ff22ffa2ffa2)
  ) CLBLM_L_X56Y97_SLICE_X85Y97_ALUT (
.I0(CLBLM_L_X56Y97_SLICE_X85Y97_BO5),
.I1(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I2(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.I3(CLBLM_L_X56Y97_SLICE_X85Y97_BO6),
.I4(CLBLM_R_X49Y108_SLICE_X75Y108_DQ),
.I5(CLBLM_R_X49Y107_SLICE_X75Y107_DQ),
.O5(CLBLM_L_X56Y97_SLICE_X85Y97_AO5),
.O6(CLBLM_L_X56Y97_SLICE_X85Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y98_SLICE_X84Y98_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X56Y98_SLICE_X84Y98_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y98_SLICE_X84Y98_AO6),
.Q(CLBLM_L_X56Y98_SLICE_X84Y98_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y98_SLICE_X84Y98_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X56Y98_SLICE_X84Y98_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y98_SLICE_X84Y98_AO5),
.Q(CLBLM_L_X56Y98_SLICE_X84Y98_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00a0a0a0a0)
  ) CLBLM_L_X56Y98_SLICE_X84Y98_DLUT (
.I0(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.I1(CLBLM_L_X60Y98_SLICE_X91Y98_CQ),
.I2(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I3(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y98_SLICE_X84Y98_DO5),
.O6(CLBLM_L_X56Y98_SLICE_X84Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff04000000)
  ) CLBLM_L_X56Y98_SLICE_X84Y98_CLUT (
.I0(CLBLM_R_X49Y107_SLICE_X75Y107_DQ),
.I1(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.I2(CLBLM_R_X49Y108_SLICE_X75Y108_DQ),
.I3(CLBLM_L_X56Y97_SLICE_X84Y97_CO5),
.I4(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I5(CLBLL_L_X54Y102_SLICE_X82Y102_BO6),
.O5(CLBLM_L_X56Y98_SLICE_X84Y98_CO5),
.O6(CLBLM_L_X56Y98_SLICE_X84Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf2f0f2f0fcf0f0f0)
  ) CLBLM_L_X56Y98_SLICE_X84Y98_BLUT (
.I0(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I1(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.I2(CLBLM_L_X56Y98_SLICE_X85Y98_BO5),
.I3(CLBLM_L_X56Y98_SLICE_X84Y98_DO5),
.I4(CLBLM_L_X56Y97_SLICE_X84Y97_AO6),
.I5(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.O5(CLBLM_L_X56Y98_SLICE_X84Y98_BO5),
.O6(CLBLM_L_X56Y98_SLICE_X84Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00050005a000a000)
  ) CLBLM_L_X56Y98_SLICE_X84Y98_ALUT (
.I0(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I1(1'b1),
.I2(CLBLM_R_X49Y107_SLICE_X75Y107_DQ),
.I3(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y98_SLICE_X84Y98_AO5),
.O6(CLBLM_L_X56Y98_SLICE_X84Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y98_SLICE_X85Y98_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y98_SLICE_X85Y98_AO5),
.Q(CLBLM_L_X56Y98_SLICE_X85Y98_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y98_SLICE_X85Y98_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y98_SLICE_X85Y98_AO6),
.Q(CLBLM_L_X56Y98_SLICE_X85Y98_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y98_SLICE_X85Y98_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y98_SLICE_X85Y98_BO6),
.Q(CLBLM_L_X56Y98_SLICE_X85Y98_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y98_SLICE_X85Y98_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y98_SLICE_X85Y98_CO6),
.Q(CLBLM_L_X56Y98_SLICE_X85Y98_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y98_SLICE_X85Y98_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y98_SLICE_X85Y98_DO6),
.Q(CLBLM_L_X56Y98_SLICE_X85Y98_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3020313030303030)
  ) CLBLM_L_X56Y98_SLICE_X85Y98_DLUT (
.I0(CLBLL_R_X57Y102_SLICE_X86Y102_CO6),
.I1(CLBLM_L_X56Y98_SLICE_X84Y98_CO6),
.I2(CLBLM_L_X56Y98_SLICE_X84Y98_BO6),
.I3(CLBLM_R_X49Y104_SLICE_X74Y104_AQ),
.I4(CLBLM_R_X49Y104_SLICE_X75Y104_AQ),
.I5(CLBLM_L_X56Y100_SLICE_X85Y100_BO6),
.O5(CLBLM_L_X56Y98_SLICE_X85Y98_DO5),
.O6(CLBLM_L_X56Y98_SLICE_X85Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf606f606f606f606)
  ) CLBLM_L_X56Y98_SLICE_X85Y98_CLUT (
.I0(CLBLL_R_X57Y103_SLICE_X86Y103_AQ),
.I1(CLBLL_R_X57Y103_SLICE_X86Y103_A5Q),
.I2(CLBLL_L_X54Y98_SLICE_X83Y98_DO6),
.I3(CLBLM_R_X49Y108_SLICE_X75Y108_DQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y98_SLICE_X85Y98_CO5),
.O6(CLBLM_L_X56Y98_SLICE_X85Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h400004000f0ff0f0)
  ) CLBLM_L_X56Y98_SLICE_X85Y98_BLUT (
.I0(CLBLL_L_X54Y98_SLICE_X83Y98_DO6),
.I1(CLBLL_L_X54Y102_SLICE_X82Y102_BO6),
.I2(CLBLL_R_X57Y103_SLICE_X86Y103_AQ),
.I3(CLBLM_R_X49Y104_SLICE_X74Y104_AQ),
.I4(CLBLL_R_X57Y103_SLICE_X86Y103_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X56Y98_SLICE_X85Y98_BO5),
.O6(CLBLM_L_X56Y98_SLICE_X85Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000044f0f0f0f8)
  ) CLBLM_L_X56Y98_SLICE_X85Y98_ALUT (
.I0(CLBLM_R_X49Y104_SLICE_X75Y104_AQ),
.I1(CLBLM_L_X56Y100_SLICE_X85Y100_BO6),
.I2(CLBLM_L_X56Y98_SLICE_X84Y98_CO6),
.I3(CLBLM_R_X49Y104_SLICE_X74Y104_AQ),
.I4(CLBLL_R_X57Y102_SLICE_X86Y102_CO6),
.I5(1'b1),
.O5(CLBLM_L_X56Y98_SLICE_X85Y98_AO5),
.O6(CLBLM_L_X56Y98_SLICE_X85Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y99_SLICE_X84Y99_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_BQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y99_SLICE_X84Y99_AO6),
.Q(CLBLM_L_X56Y99_SLICE_X84Y99_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y99_SLICE_X84Y99_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_BQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y99_SLICE_X84Y99_BO6),
.Q(CLBLM_L_X56Y99_SLICE_X84Y99_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y99_SLICE_X84Y99_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y99_SLICE_X84Y99_DO5),
.O6(CLBLM_L_X56Y99_SLICE_X84Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00882200c0002200)
  ) CLBLM_L_X56Y99_SLICE_X84Y99_CLUT (
.I0(CLBLM_L_X56Y97_SLICE_X84Y97_CO5),
.I1(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.I2(CLBLM_L_X56Y97_SLICE_X85Y97_BO5),
.I3(CLBLM_R_X49Y107_SLICE_X75Y107_DQ),
.I4(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I5(CLBLM_R_X49Y108_SLICE_X75Y108_DQ),
.O5(CLBLM_L_X56Y99_SLICE_X84Y99_CO5),
.O6(CLBLM_L_X56Y99_SLICE_X84Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333333333333)
  ) CLBLM_L_X56Y99_SLICE_X84Y99_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X54Y98_SLICE_X82Y98_AO6),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y99_SLICE_X84Y99_BO5),
.O6(CLBLM_L_X56Y99_SLICE_X84Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff08ff00000808)
  ) CLBLM_L_X56Y99_SLICE_X84Y99_ALUT (
.I0(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I1(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.I2(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.I3(CLBLL_L_X54Y98_SLICE_X82Y98_AO6),
.I4(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.I5(CLBLM_R_X49Y108_SLICE_X75Y108_DQ),
.O5(CLBLM_L_X56Y99_SLICE_X84Y99_AO5),
.O6(CLBLM_L_X56Y99_SLICE_X84Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y99_SLICE_X85Y99_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y99_SLICE_X85Y99_AQ),
.Q(CLBLM_L_X56Y99_SLICE_X85Y99_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y99_SLICE_X85Y99_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y99_SLICE_X85Y99_AO6),
.Q(CLBLM_L_X56Y99_SLICE_X85Y99_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y99_SLICE_X85Y99_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y99_SLICE_X85Y99_BO6),
.Q(CLBLM_L_X56Y99_SLICE_X85Y99_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y99_SLICE_X85Y99_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y99_SLICE_X85Y99_CO6),
.Q(CLBLM_L_X56Y99_SLICE_X85Y99_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y99_SLICE_X85Y99_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y99_SLICE_X85Y99_DO5),
.O6(CLBLM_L_X56Y99_SLICE_X85Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0101000000000000)
  ) CLBLM_L_X56Y99_SLICE_X85Y99_CLUT (
.I0(CLBLM_R_X49Y106_SLICE_X75Y106_CQ),
.I1(CLBLL_L_X54Y102_SLICE_X82Y102_AO5),
.I2(CLBLM_R_X49Y104_SLICE_X75Y104_DQ),
.I3(1'b1),
.I4(CLBLM_R_X49Y104_SLICE_X75Y104_AQ),
.I5(CLBLM_L_X56Y102_SLICE_X85Y102_BO6),
.O5(CLBLM_L_X56Y99_SLICE_X85Y99_CO5),
.O6(CLBLM_L_X56Y99_SLICE_X85Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f800000088)
  ) CLBLM_L_X56Y99_SLICE_X85Y99_BLUT (
.I0(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I1(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.I2(CLBLM_L_X56Y97_SLICE_X84Y97_CO5),
.I3(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.I4(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.I5(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.O5(CLBLM_L_X56Y99_SLICE_X85Y99_BO5),
.O6(CLBLM_L_X56Y99_SLICE_X85Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff00ff00)
  ) CLBLM_L_X56Y99_SLICE_X85Y99_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_R_X57Y102_SLICE_X86Y102_AO6),
.I4(1'b1),
.I5(CLBLL_L_X52Y99_SLICE_X79Y99_AO6),
.O5(CLBLM_L_X56Y99_SLICE_X85Y99_AO5),
.O6(CLBLM_L_X56Y99_SLICE_X85Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y100_SLICE_X84Y100_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X56Y102_SLICE_X85Y102_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y100_SLICE_X84Y100_A_XOR),
.Q(CLBLM_L_X56Y100_SLICE_X84Y100_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y100_SLICE_X84Y100_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X56Y102_SLICE_X85Y102_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y100_SLICE_X84Y100_B_XOR),
.Q(CLBLM_L_X56Y100_SLICE_X84Y100_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y100_SLICE_X84Y100_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X56Y102_SLICE_X85Y102_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y100_SLICE_X84Y100_C_XOR),
.Q(CLBLM_L_X56Y100_SLICE_X84Y100_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y100_SLICE_X84Y100_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X56Y102_SLICE_X85Y102_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y100_SLICE_X84Y100_D_XOR),
.Q(CLBLM_L_X56Y100_SLICE_X84Y100_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X56Y100_SLICE_X84Y100_CARRY4 (
.CI(1'b0),
.CO({CLBLM_L_X56Y100_SLICE_X84Y100_D_CY, CLBLM_L_X56Y100_SLICE_X84Y100_C_CY, CLBLM_L_X56Y100_SLICE_X84Y100_B_CY, CLBLM_L_X56Y100_SLICE_X84Y100_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, CLBLM_L_X56Y100_SLICE_X84Y100_AO5}),
.O({CLBLM_L_X56Y100_SLICE_X84Y100_D_XOR, CLBLM_L_X56Y100_SLICE_X84Y100_C_XOR, CLBLM_L_X56Y100_SLICE_X84Y100_B_XOR, CLBLM_L_X56Y100_SLICE_X84Y100_A_XOR}),
.S({CLBLM_L_X56Y100_SLICE_X84Y100_DO6, CLBLM_L_X56Y100_SLICE_X84Y100_CO6, CLBLM_L_X56Y100_SLICE_X84Y100_BO6, CLBLM_L_X56Y100_SLICE_X84Y100_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000505000005050)
  ) CLBLM_L_X56Y100_SLICE_X84Y100_DLUT (
.I0(CLBLM_L_X56Y102_SLICE_X85Y102_AQ),
.I1(1'b1),
.I2(CLBLM_L_X56Y100_SLICE_X84Y100_DQ),
.I3(1'b1),
.I4(CLBLM_L_X56Y102_SLICE_X85Y102_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X56Y100_SLICE_X84Y100_DO5),
.O6(CLBLM_L_X56Y100_SLICE_X84Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0404040404040404)
  ) CLBLM_L_X56Y100_SLICE_X84Y100_CLUT (
.I0(CLBLM_L_X56Y102_SLICE_X85Y102_AQ),
.I1(CLBLM_L_X56Y100_SLICE_X84Y100_CQ),
.I2(CLBLM_L_X56Y102_SLICE_X85Y102_A5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y100_SLICE_X84Y100_CO5),
.O6(CLBLM_L_X56Y100_SLICE_X84Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0404040404040404)
  ) CLBLM_L_X56Y100_SLICE_X84Y100_BLUT (
.I0(CLBLM_L_X56Y102_SLICE_X85Y102_A5Q),
.I1(CLBLM_L_X56Y100_SLICE_X84Y100_BQ),
.I2(CLBLM_L_X56Y102_SLICE_X85Y102_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y100_SLICE_X84Y100_BO5),
.O6(CLBLM_L_X56Y100_SLICE_X84Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000050500005555)
  ) CLBLM_L_X56Y100_SLICE_X84Y100_ALUT (
.I0(CLBLM_L_X56Y102_SLICE_X85Y102_A5Q),
.I1(1'b1),
.I2(CLBLM_L_X56Y100_SLICE_X84Y100_AQ),
.I3(1'b1),
.I4(CLBLM_L_X56Y102_SLICE_X85Y102_AQ),
.I5(1'b1),
.O5(CLBLM_L_X56Y100_SLICE_X84Y100_AO5),
.O6(CLBLM_L_X56Y100_SLICE_X84Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y100_SLICE_X85Y100_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X56Y98_SLICE_X84Y98_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y100_SLICE_X85Y100_BO5),
.Q(CLBLM_L_X56Y100_SLICE_X85Y100_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y100_SLICE_X85Y100_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X56Y98_SLICE_X84Y98_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y100_SLICE_X85Y100_AO6),
.Q(CLBLM_L_X56Y100_SLICE_X85Y100_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y100_SLICE_X85Y100_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X56Y98_SLICE_X84Y98_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y100_SLICE_X85Y100_AO5),
.Q(CLBLM_L_X56Y100_SLICE_X85Y100_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y100_SLICE_X85Y100_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X56Y98_SLICE_X84Y98_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y97_SLICE_X84Y97_AO6),
.Q(CLBLM_L_X56Y100_SLICE_X85Y100_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y100_SLICE_X85Y100_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y100_SLICE_X85Y100_DO5),
.O6(CLBLM_L_X56Y100_SLICE_X85Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y100_SLICE_X85Y100_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y100_SLICE_X85Y100_CO5),
.O6(CLBLM_L_X56Y100_SLICE_X85Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010011110000)
  ) CLBLM_L_X56Y100_SLICE_X85Y100_BLUT (
.I0(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I1(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.I2(CLBLM_R_X49Y108_SLICE_X75Y108_DQ),
.I3(CLBLM_L_X56Y97_SLICE_X84Y97_CO5),
.I4(CLBLM_R_X49Y107_SLICE_X75Y107_DQ),
.I5(1'b1),
.O5(CLBLM_L_X56Y100_SLICE_X85Y100_BO5),
.O6(CLBLM_L_X56Y100_SLICE_X85Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5500000000aa0000)
  ) CLBLM_L_X56Y100_SLICE_X85Y100_ALUT (
.I0(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.I4(CLBLM_R_X49Y107_SLICE_X75Y107_DQ),
.I5(1'b1),
.O5(CLBLM_L_X56Y100_SLICE_X85Y100_AO5),
.O6(CLBLM_L_X56Y100_SLICE_X85Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y101_SLICE_X84Y101_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X56Y102_SLICE_X85Y102_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y101_SLICE_X84Y101_A_XOR),
.Q(CLBLM_L_X56Y101_SLICE_X84Y101_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y101_SLICE_X84Y101_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X56Y102_SLICE_X85Y102_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y101_SLICE_X84Y101_B_XOR),
.Q(CLBLM_L_X56Y101_SLICE_X84Y101_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y101_SLICE_X84Y101_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X56Y102_SLICE_X85Y102_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y101_SLICE_X84Y101_C_XOR),
.Q(CLBLM_L_X56Y101_SLICE_X84Y101_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y101_SLICE_X84Y101_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X56Y102_SLICE_X85Y102_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y101_SLICE_X84Y101_D_XOR),
.Q(CLBLM_L_X56Y101_SLICE_X84Y101_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X56Y101_SLICE_X84Y101_CARRY4 (
.CI(CLBLM_L_X56Y100_SLICE_X84Y100_COUT),
.CO({CLBLM_L_X56Y101_SLICE_X84Y101_D_CY, CLBLM_L_X56Y101_SLICE_X84Y101_C_CY, CLBLM_L_X56Y101_SLICE_X84Y101_B_CY, CLBLM_L_X56Y101_SLICE_X84Y101_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_L_X56Y101_SLICE_X84Y101_D_XOR, CLBLM_L_X56Y101_SLICE_X84Y101_C_XOR, CLBLM_L_X56Y101_SLICE_X84Y101_B_XOR, CLBLM_L_X56Y101_SLICE_X84Y101_A_XOR}),
.S({CLBLM_L_X56Y101_SLICE_X84Y101_DO6, CLBLM_L_X56Y101_SLICE_X84Y101_CO6, CLBLM_L_X56Y101_SLICE_X84Y101_BO6, CLBLM_L_X56Y101_SLICE_X84Y101_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000505000005050)
  ) CLBLM_L_X56Y101_SLICE_X84Y101_DLUT (
.I0(CLBLM_L_X56Y102_SLICE_X85Y102_AQ),
.I1(1'b1),
.I2(CLBLM_L_X56Y101_SLICE_X84Y101_DQ),
.I3(1'b1),
.I4(CLBLM_L_X56Y102_SLICE_X85Y102_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X56Y101_SLICE_X84Y101_DO5),
.O6(CLBLM_L_X56Y101_SLICE_X84Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000444400004444)
  ) CLBLM_L_X56Y101_SLICE_X84Y101_CLUT (
.I0(CLBLM_L_X56Y102_SLICE_X85Y102_AQ),
.I1(CLBLM_L_X56Y101_SLICE_X84Y101_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X56Y102_SLICE_X85Y102_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X56Y101_SLICE_X84Y101_CO5),
.O6(CLBLM_L_X56Y101_SLICE_X84Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0404040404040404)
  ) CLBLM_L_X56Y101_SLICE_X84Y101_BLUT (
.I0(CLBLM_L_X56Y102_SLICE_X85Y102_A5Q),
.I1(CLBLM_L_X56Y101_SLICE_X84Y101_BQ),
.I2(CLBLM_L_X56Y102_SLICE_X85Y102_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y101_SLICE_X84Y101_BO5),
.O6(CLBLM_L_X56Y101_SLICE_X84Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000505000005050)
  ) CLBLM_L_X56Y101_SLICE_X84Y101_ALUT (
.I0(CLBLM_L_X56Y102_SLICE_X85Y102_A5Q),
.I1(1'b1),
.I2(CLBLM_L_X56Y101_SLICE_X84Y101_AQ),
.I3(1'b1),
.I4(CLBLM_L_X56Y102_SLICE_X85Y102_AQ),
.I5(1'b1),
.O5(CLBLM_L_X56Y101_SLICE_X84Y101_AO5),
.O6(CLBLM_L_X56Y101_SLICE_X84Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y101_SLICE_X85Y101_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLL_R_X57Y100_SLICE_X87Y100_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y101_SLICE_X85Y101_AO6),
.Q(CLBLM_L_X56Y101_SLICE_X85Y101_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y101_SLICE_X85Y101_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLL_R_X57Y100_SLICE_X87Y100_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y101_SLICE_X85Y101_BO6),
.Q(CLBLM_L_X56Y101_SLICE_X85Y101_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y101_SLICE_X85Y101_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLL_R_X57Y100_SLICE_X87Y100_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y101_SLICE_X85Y101_CO6),
.Q(CLBLM_L_X56Y101_SLICE_X85Y101_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y101_SLICE_X85Y101_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLL_R_X57Y100_SLICE_X87Y100_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y101_SLICE_X85Y101_DO6),
.Q(CLBLM_L_X56Y101_SLICE_X85Y101_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcbfb0b3bc8f80838)
  ) CLBLM_L_X56Y101_SLICE_X85Y101_DLUT (
.I0(CLBLM_L_X62Y101_SLICE_X92Y101_DO5),
.I1(CLBLL_L_X54Y99_SLICE_X82Y99_CQ),
.I2(CLBLM_L_X56Y99_SLICE_X85Y99_BQ),
.I3(CLBLM_L_X56Y100_SLICE_X85Y100_CQ),
.I4(CLBLM_L_X64Y100_SLICE_X97Y100_BQ),
.I5(CLBLM_R_X59Y98_SLICE_X89Y98_C5Q),
.O5(CLBLM_L_X56Y101_SLICE_X85Y101_DO5),
.O6(CLBLM_L_X56Y101_SLICE_X85Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd1ffd133d1ccd100)
  ) CLBLM_L_X56Y101_SLICE_X85Y101_CLUT (
.I0(CLBLL_L_X54Y101_SLICE_X82Y101_AQ),
.I1(CLBLL_L_X54Y99_SLICE_X82Y99_CQ),
.I2(CLBLM_L_X62Y101_SLICE_X93Y101_AQ),
.I3(CLBLM_L_X56Y99_SLICE_X85Y99_BQ),
.I4(CLBLM_L_X60Y101_SLICE_X91Y101_CO6),
.I5(CLBLM_R_X59Y98_SLICE_X89Y98_BQ),
.O5(CLBLM_L_X56Y101_SLICE_X85Y101_CO5),
.O6(CLBLM_L_X56Y101_SLICE_X85Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0fff0fcfc0c0c)
  ) CLBLM_L_X56Y101_SLICE_X85Y101_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X59Y98_SLICE_X89Y98_C5Q),
.I2(CLBLL_L_X54Y98_SLICE_X83Y98_BQ),
.I3(CLBLM_L_X56Y100_SLICE_X85Y100_CQ),
.I4(CLBLM_L_X62Y101_SLICE_X92Y101_DO5),
.I5(CLBLL_L_X54Y99_SLICE_X82Y99_AQ),
.O5(CLBLM_L_X56Y101_SLICE_X85Y101_BO5),
.O6(CLBLM_L_X56Y101_SLICE_X85Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff0f0acacacac)
  ) CLBLM_L_X56Y101_SLICE_X85Y101_ALUT (
.I0(CLBLM_L_X60Y101_SLICE_X91Y101_CO6),
.I1(CLBLM_R_X59Y98_SLICE_X89Y98_BQ),
.I2(CLBLL_L_X54Y98_SLICE_X83Y98_BQ),
.I3(1'b1),
.I4(CLBLL_L_X54Y101_SLICE_X82Y101_AQ),
.I5(CLBLL_L_X54Y99_SLICE_X82Y99_AQ),
.O5(CLBLM_L_X56Y101_SLICE_X85Y101_AO5),
.O6(CLBLM_L_X56Y101_SLICE_X85Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y102_SLICE_X84Y102_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X56Y102_SLICE_X85Y102_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y102_SLICE_X84Y102_A_XOR),
.Q(CLBLM_L_X56Y102_SLICE_X84Y102_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y102_SLICE_X84Y102_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X56Y102_SLICE_X85Y102_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y102_SLICE_X84Y102_B_XOR),
.Q(CLBLM_L_X56Y102_SLICE_X84Y102_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y102_SLICE_X84Y102_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X56Y102_SLICE_X85Y102_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y102_SLICE_X84Y102_C_XOR),
.Q(CLBLM_L_X56Y102_SLICE_X84Y102_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y102_SLICE_X84Y102_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X56Y102_SLICE_X85Y102_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y102_SLICE_X84Y102_D_XOR),
.Q(CLBLM_L_X56Y102_SLICE_X84Y102_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X56Y102_SLICE_X84Y102_CARRY4 (
.CI(CLBLM_L_X56Y101_SLICE_X84Y101_COUT),
.CO({CLBLM_L_X56Y102_SLICE_X84Y102_D_CY, CLBLM_L_X56Y102_SLICE_X84Y102_C_CY, CLBLM_L_X56Y102_SLICE_X84Y102_B_CY, CLBLM_L_X56Y102_SLICE_X84Y102_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_L_X56Y102_SLICE_X84Y102_D_XOR, CLBLM_L_X56Y102_SLICE_X84Y102_C_XOR, CLBLM_L_X56Y102_SLICE_X84Y102_B_XOR, CLBLM_L_X56Y102_SLICE_X84Y102_A_XOR}),
.S({CLBLM_L_X56Y102_SLICE_X84Y102_DO6, CLBLM_L_X56Y102_SLICE_X84Y102_CO6, CLBLM_L_X56Y102_SLICE_X84Y102_BO6, CLBLM_L_X56Y102_SLICE_X84Y102_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1010101010101010)
  ) CLBLM_L_X56Y102_SLICE_X84Y102_DLUT (
.I0(CLBLM_L_X56Y102_SLICE_X85Y102_AQ),
.I1(CLBLM_L_X56Y102_SLICE_X85Y102_A5Q),
.I2(CLBLM_L_X56Y102_SLICE_X84Y102_DQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y102_SLICE_X84Y102_DO5),
.O6(CLBLM_L_X56Y102_SLICE_X84Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000044444444)
  ) CLBLM_L_X56Y102_SLICE_X84Y102_CLUT (
.I0(CLBLM_L_X56Y102_SLICE_X85Y102_AQ),
.I1(CLBLM_L_X56Y102_SLICE_X84Y102_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X56Y102_SLICE_X85Y102_A5Q),
.O5(CLBLM_L_X56Y102_SLICE_X84Y102_CO5),
.O6(CLBLM_L_X56Y102_SLICE_X84Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000c0c00000c0c)
  ) CLBLM_L_X56Y102_SLICE_X84Y102_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X56Y102_SLICE_X84Y102_BQ),
.I2(CLBLM_L_X56Y102_SLICE_X85Y102_A5Q),
.I3(1'b1),
.I4(CLBLM_L_X56Y102_SLICE_X85Y102_AQ),
.I5(1'b1),
.O5(CLBLM_L_X56Y102_SLICE_X84Y102_BO5),
.O6(CLBLM_L_X56Y102_SLICE_X84Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000f0000000f0)
  ) CLBLM_L_X56Y102_SLICE_X84Y102_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X56Y102_SLICE_X84Y102_AQ),
.I3(CLBLM_L_X56Y102_SLICE_X85Y102_A5Q),
.I4(CLBLM_L_X56Y102_SLICE_X85Y102_AQ),
.I5(1'b1),
.O5(CLBLM_L_X56Y102_SLICE_X84Y102_AO5),
.O6(CLBLM_L_X56Y102_SLICE_X84Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y102_SLICE_X85Y102_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y102_SLICE_X85Y102_AO5),
.Q(CLBLM_L_X56Y102_SLICE_X85Y102_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y102_SLICE_X85Y102_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y102_SLICE_X85Y102_AO6),
.Q(CLBLM_L_X56Y102_SLICE_X85Y102_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y102_SLICE_X85Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y102_SLICE_X85Y102_DO5),
.O6(CLBLM_L_X56Y102_SLICE_X85Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffafffafffafffa)
  ) CLBLM_L_X56Y102_SLICE_X85Y102_CLUT (
.I0(CLBLM_R_X63Y100_SLICE_X94Y100_AQ),
.I1(1'b1),
.I2(CLBLM_L_X56Y102_SLICE_X85Y102_AQ),
.I3(CLBLM_L_X56Y102_SLICE_X85Y102_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y102_SLICE_X85Y102_CO5),
.O6(CLBLM_L_X56Y102_SLICE_X85Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000400)
  ) CLBLM_L_X56Y102_SLICE_X85Y102_BLUT (
.I0(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I1(CLBLM_R_X49Y104_SLICE_X74Y104_AQ),
.I2(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.I3(CLBLM_L_X56Y97_SLICE_X84Y97_CO5),
.I4(CLBLM_R_X49Y107_SLICE_X75Y107_DQ),
.I5(CLBLM_R_X49Y108_SLICE_X75Y108_DQ),
.O5(CLBLM_L_X56Y102_SLICE_X85Y102_BO5),
.O6(CLBLM_L_X56Y102_SLICE_X85Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc000c000cc000000)
  ) CLBLM_L_X56Y102_SLICE_X85Y102_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I2(CLBLM_L_X56Y98_SLICE_X85Y98_AQ),
.I3(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.I4(CLBLM_L_X56Y99_SLICE_X85Y99_CQ),
.I5(1'b1),
.O5(CLBLM_L_X56Y102_SLICE_X85Y102_AO5),
.O6(CLBLM_L_X56Y102_SLICE_X85Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y103_SLICE_X84Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X56Y102_SLICE_X85Y102_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y103_SLICE_X84Y103_A_XOR),
.Q(CLBLM_L_X56Y103_SLICE_X84Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y103_SLICE_X84Y103_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X56Y102_SLICE_X85Y102_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y103_SLICE_X84Y103_B_XOR),
.Q(CLBLM_L_X56Y103_SLICE_X84Y103_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y103_SLICE_X84Y103_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X56Y102_SLICE_X85Y102_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y103_SLICE_X84Y103_C_XOR),
.Q(CLBLM_L_X56Y103_SLICE_X84Y103_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y103_SLICE_X84Y103_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X56Y102_SLICE_X85Y102_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y103_SLICE_X84Y103_D_XOR),
.Q(CLBLM_L_X56Y103_SLICE_X84Y103_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X56Y103_SLICE_X84Y103_CARRY4 (
.CI(CLBLM_L_X56Y102_SLICE_X84Y102_COUT),
.CO({CLBLM_L_X56Y103_SLICE_X84Y103_D_CY, CLBLM_L_X56Y103_SLICE_X84Y103_C_CY, CLBLM_L_X56Y103_SLICE_X84Y103_B_CY, CLBLM_L_X56Y103_SLICE_X84Y103_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_L_X56Y103_SLICE_X84Y103_D_XOR, CLBLM_L_X56Y103_SLICE_X84Y103_C_XOR, CLBLM_L_X56Y103_SLICE_X84Y103_B_XOR, CLBLM_L_X56Y103_SLICE_X84Y103_A_XOR}),
.S({CLBLM_L_X56Y103_SLICE_X84Y103_DO6, CLBLM_L_X56Y103_SLICE_X84Y103_CO6, CLBLM_L_X56Y103_SLICE_X84Y103_BO6, CLBLM_L_X56Y103_SLICE_X84Y103_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000505000005050)
  ) CLBLM_L_X56Y103_SLICE_X84Y103_DLUT (
.I0(CLBLM_L_X56Y102_SLICE_X85Y102_A5Q),
.I1(1'b1),
.I2(CLBLM_L_X56Y103_SLICE_X84Y103_DQ),
.I3(1'b1),
.I4(CLBLM_L_X56Y102_SLICE_X85Y102_AQ),
.I5(1'b1),
.O5(CLBLM_L_X56Y103_SLICE_X84Y103_DO5),
.O6(CLBLM_L_X56Y103_SLICE_X84Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000444400004444)
  ) CLBLM_L_X56Y103_SLICE_X84Y103_CLUT (
.I0(CLBLM_L_X56Y102_SLICE_X85Y102_A5Q),
.I1(CLBLM_L_X56Y103_SLICE_X84Y103_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X56Y102_SLICE_X85Y102_AQ),
.I5(1'b1),
.O5(CLBLM_L_X56Y103_SLICE_X84Y103_CO5),
.O6(CLBLM_L_X56Y103_SLICE_X84Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0404040404040404)
  ) CLBLM_L_X56Y103_SLICE_X84Y103_BLUT (
.I0(CLBLM_L_X56Y102_SLICE_X85Y102_AQ),
.I1(CLBLM_L_X56Y103_SLICE_X84Y103_BQ),
.I2(CLBLM_L_X56Y102_SLICE_X85Y102_A5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y103_SLICE_X84Y103_BO5),
.O6(CLBLM_L_X56Y103_SLICE_X84Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h1010101010101010)
  ) CLBLM_L_X56Y103_SLICE_X84Y103_ALUT (
.I0(CLBLM_L_X56Y102_SLICE_X85Y102_AQ),
.I1(CLBLM_L_X56Y102_SLICE_X85Y102_A5Q),
.I2(CLBLM_L_X56Y103_SLICE_X84Y103_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y103_SLICE_X84Y103_AO5),
.O6(CLBLM_L_X56Y103_SLICE_X84Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X56Y103_SLICE_X85Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X56Y103_SLICE_X85Y103_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y103_SLICE_X85Y103_AO6),
.Q(CLBLM_L_X56Y103_SLICE_X85Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X56Y103_SLICE_X85Y103_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X56Y103_SLICE_X85Y103_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y103_SLICE_X85Y103_BO6),
.Q(CLBLM_L_X56Y103_SLICE_X85Y103_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y103_SLICE_X85Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y103_SLICE_X85Y103_DO5),
.O6(CLBLM_L_X56Y103_SLICE_X85Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000000000)
  ) CLBLM_L_X56Y103_SLICE_X85Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.O5(CLBLM_L_X56Y103_SLICE_X85Y103_CO5),
.O6(CLBLM_L_X56Y103_SLICE_X85Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ccaaf0f0ccaa)
  ) CLBLM_L_X56Y103_SLICE_X85Y103_BLUT (
.I0(CLBLL_L_X54Y105_SLICE_X82Y105_B_XOR),
.I1(CLBLM_L_X56Y103_SLICE_X85Y103_BQ),
.I2(CLBLM_L_X50Y106_SLICE_X76Y106_AQ),
.I3(CLBLL_L_X54Y101_SLICE_X83Y101_BO6),
.I4(CLBLM_L_X62Y100_SLICE_X92Y100_AO5),
.I5(1'b1),
.O5(CLBLM_L_X56Y103_SLICE_X85Y103_BO5),
.O6(CLBLM_L_X56Y103_SLICE_X85Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8bbb888b8bbb888)
  ) CLBLM_L_X56Y103_SLICE_X85Y103_ALUT (
.I0(CLBLM_L_X50Y106_SLICE_X76Y106_AQ),
.I1(CLBLM_L_X60Y99_SLICE_X90Y99_AO5),
.I2(CLBLM_L_X56Y103_SLICE_X85Y103_AQ),
.I3(CLBLL_L_X54Y101_SLICE_X83Y101_BO6),
.I4(CLBLL_L_X54Y107_SLICE_X82Y107_B_XOR),
.I5(1'b1),
.O5(CLBLM_L_X56Y103_SLICE_X85Y103_AO5),
.O6(CLBLM_L_X56Y103_SLICE_X85Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y104_SLICE_X84Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X56Y102_SLICE_X85Y102_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y104_SLICE_X84Y104_A_XOR),
.Q(CLBLM_L_X56Y104_SLICE_X84Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X56Y104_SLICE_X84Y104_CARRY4 (
.CI(CLBLM_L_X56Y103_SLICE_X84Y103_COUT),
.CO({CLBLM_L_X56Y104_SLICE_X84Y104_D_CY, CLBLM_L_X56Y104_SLICE_X84Y104_C_CY, CLBLM_L_X56Y104_SLICE_X84Y104_B_CY, CLBLM_L_X56Y104_SLICE_X84Y104_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_L_X56Y104_SLICE_X84Y104_D_XOR, CLBLM_L_X56Y104_SLICE_X84Y104_C_XOR, CLBLM_L_X56Y104_SLICE_X84Y104_B_XOR, CLBLM_L_X56Y104_SLICE_X84Y104_A_XOR}),
.S({CLBLM_L_X56Y104_SLICE_X84Y104_DO6, CLBLM_L_X56Y104_SLICE_X84Y104_CO6, CLBLM_L_X56Y104_SLICE_X84Y104_BO6, CLBLM_L_X56Y104_SLICE_X84Y104_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y104_SLICE_X84Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y104_SLICE_X84Y104_DO5),
.O6(CLBLM_L_X56Y104_SLICE_X84Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y104_SLICE_X84Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y104_SLICE_X84Y104_CO5),
.O6(CLBLM_L_X56Y104_SLICE_X84Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y104_SLICE_X84Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y104_SLICE_X84Y104_BO5),
.O6(CLBLM_L_X56Y104_SLICE_X84Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000f0000000f0)
  ) CLBLM_L_X56Y104_SLICE_X84Y104_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X56Y104_SLICE_X84Y104_AQ),
.I3(CLBLM_L_X56Y102_SLICE_X85Y102_AQ),
.I4(CLBLM_L_X56Y102_SLICE_X85Y102_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X56Y104_SLICE_X84Y104_AO5),
.O6(CLBLM_L_X56Y104_SLICE_X84Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X56Y104_SLICE_X85Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X56Y103_SLICE_X85Y103_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y104_SLICE_X85Y104_AO6),
.Q(CLBLM_L_X56Y104_SLICE_X85Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y104_SLICE_X85Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y104_SLICE_X85Y104_DO5),
.O6(CLBLM_L_X56Y104_SLICE_X85Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y104_SLICE_X85Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y104_SLICE_X85Y104_CO5),
.O6(CLBLM_L_X56Y104_SLICE_X85Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y104_SLICE_X85Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y104_SLICE_X85Y104_BO5),
.O6(CLBLM_L_X56Y104_SLICE_X85Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcff3033fccc3000)
  ) CLBLM_L_X56Y104_SLICE_X85Y104_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X62Y100_SLICE_X92Y100_AO5),
.I2(CLBLM_L_X56Y104_SLICE_X85Y104_AQ),
.I3(CLBLL_L_X54Y101_SLICE_X83Y101_BO6),
.I4(CLBLM_L_X50Y107_SLICE_X77Y107_AQ),
.I5(CLBLL_L_X54Y106_SLICE_X82Y106_A_XOR),
.O5(CLBLM_L_X56Y104_SLICE_X85Y104_AO5),
.O6(CLBLM_L_X56Y104_SLICE_X85Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X56Y105_SLICE_X84Y105_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X56Y103_SLICE_X85Y103_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y105_SLICE_X84Y105_AO6),
.Q(CLBLM_L_X56Y105_SLICE_X84Y105_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X56Y105_SLICE_X84Y105_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X56Y103_SLICE_X85Y103_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y105_SLICE_X84Y105_BO6),
.Q(CLBLM_L_X56Y105_SLICE_X84Y105_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X56Y105_SLICE_X84Y105_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X56Y103_SLICE_X85Y103_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y105_SLICE_X84Y105_CO6),
.Q(CLBLM_L_X56Y105_SLICE_X84Y105_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y105_SLICE_X84Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y105_SLICE_X84Y105_DO5),
.O6(CLBLM_L_X56Y105_SLICE_X84Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ddf0ddf088f088)
  ) CLBLM_L_X56Y105_SLICE_X84Y105_CLUT (
.I0(CLBLL_L_X54Y101_SLICE_X83Y101_BO6),
.I1(CLBLM_L_X56Y105_SLICE_X84Y105_CQ),
.I2(CLBLM_L_X50Y107_SLICE_X76Y107_BQ),
.I3(CLBLM_L_X60Y99_SLICE_X90Y99_AO5),
.I4(1'b1),
.I5(CLBLL_L_X54Y107_SLICE_X82Y107_D_XOR),
.O5(CLBLM_L_X56Y105_SLICE_X84Y105_CO5),
.O6(CLBLM_L_X56Y105_SLICE_X84Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00ccccaaaa)
  ) CLBLM_L_X56Y105_SLICE_X84Y105_BLUT (
.I0(CLBLL_L_X54Y107_SLICE_X82Y107_C_XOR),
.I1(CLBLM_L_X56Y105_SLICE_X84Y105_BQ),
.I2(1'b1),
.I3(CLBLM_L_X50Y106_SLICE_X76Y106_CQ),
.I4(CLBLL_L_X54Y101_SLICE_X83Y101_BO6),
.I5(CLBLM_L_X60Y99_SLICE_X90Y99_AO5),
.O5(CLBLM_L_X56Y105_SLICE_X84Y105_BO5),
.O6(CLBLM_L_X56Y105_SLICE_X84Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaffaaf0aa00)
  ) CLBLM_L_X56Y105_SLICE_X84Y105_ALUT (
.I0(CLBLM_R_X49Y106_SLICE_X74Y106_AQ),
.I1(1'b1),
.I2(CLBLM_L_X56Y105_SLICE_X84Y105_AQ),
.I3(CLBLM_L_X60Y99_SLICE_X90Y99_AO5),
.I4(CLBLL_L_X54Y101_SLICE_X83Y101_BO6),
.I5(CLBLL_L_X54Y107_SLICE_X82Y107_A_XOR),
.O5(CLBLM_L_X56Y105_SLICE_X84Y105_AO5),
.O6(CLBLM_L_X56Y105_SLICE_X84Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X56Y105_SLICE_X85Y105_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X56Y103_SLICE_X85Y103_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y105_SLICE_X85Y105_AO6),
.Q(CLBLM_L_X56Y105_SLICE_X85Y105_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X56Y105_SLICE_X85Y105_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X56Y103_SLICE_X85Y103_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y105_SLICE_X85Y105_BO6),
.Q(CLBLM_L_X56Y105_SLICE_X85Y105_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X56Y105_SLICE_X85Y105_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X56Y103_SLICE_X85Y103_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y105_SLICE_X85Y105_CO6),
.Q(CLBLM_L_X56Y105_SLICE_X85Y105_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X56Y105_SLICE_X85Y105_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X56Y103_SLICE_X85Y103_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y105_SLICE_X85Y105_DO6),
.Q(CLBLM_L_X56Y105_SLICE_X85Y105_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00f0f06666)
  ) CLBLM_L_X56Y105_SLICE_X85Y105_DLUT (
.I0(CLBLM_R_X53Y103_SLICE_X81Y103_D_XOR),
.I1(CLBLM_R_X53Y106_SLICE_X81Y106_A_XOR),
.I2(CLBLM_L_X56Y105_SLICE_X85Y105_DQ),
.I3(CLBLM_R_X49Y106_SLICE_X74Y106_AQ),
.I4(CLBLL_L_X54Y101_SLICE_X83Y101_BO6),
.I5(CLBLM_L_X62Y100_SLICE_X92Y100_AO5),
.O5(CLBLM_L_X56Y105_SLICE_X85Y105_DO5),
.O6(CLBLM_L_X56Y105_SLICE_X85Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heeff4455eeaa4400)
  ) CLBLM_L_X56Y105_SLICE_X85Y105_CLUT (
.I0(CLBLM_L_X62Y100_SLICE_X92Y100_AO5),
.I1(CLBLM_L_X56Y105_SLICE_X85Y105_CQ),
.I2(1'b1),
.I3(CLBLL_L_X54Y101_SLICE_X83Y101_BO6),
.I4(CLBLM_L_X50Y107_SLICE_X76Y107_BQ),
.I5(CLBLL_L_X54Y105_SLICE_X82Y105_D_XOR),
.O5(CLBLM_L_X56Y105_SLICE_X85Y105_CO5),
.O6(CLBLM_L_X56Y105_SLICE_X85Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00cfcfff00c0c0)
  ) CLBLM_L_X56Y105_SLICE_X85Y105_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X56Y105_SLICE_X85Y105_BQ),
.I2(CLBLL_L_X54Y101_SLICE_X83Y101_BO6),
.I3(CLBLM_L_X50Y106_SLICE_X76Y106_CQ),
.I4(CLBLM_L_X62Y100_SLICE_X92Y100_AO5),
.I5(CLBLL_L_X54Y105_SLICE_X82Y105_C_XOR),
.O5(CLBLM_L_X56Y105_SLICE_X85Y105_BO5),
.O6(CLBLM_L_X56Y105_SLICE_X85Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd31fd31ec20ec20)
  ) CLBLM_L_X56Y105_SLICE_X85Y105_ALUT (
.I0(CLBLL_L_X54Y101_SLICE_X83Y101_BO6),
.I1(CLBLM_L_X60Y99_SLICE_X90Y99_AO5),
.I2(CLBLM_L_X56Y105_SLICE_X85Y105_AQ),
.I3(CLBLM_L_X50Y105_SLICE_X77Y105_AQ),
.I4(1'b1),
.I5(CLBLL_L_X54Y106_SLICE_X82Y106_C_XOR),
.O5(CLBLM_L_X56Y105_SLICE_X85Y105_AO5),
.O6(CLBLM_L_X56Y105_SLICE_X85Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X56Y111_SLICE_X84Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_R_X49Y111_SLICE_X75Y111_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y111_SLICE_X84Y111_AO6),
.Q(CLBLM_L_X56Y111_SLICE_X84Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y111_SLICE_X84Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y111_SLICE_X84Y111_DO5),
.O6(CLBLM_L_X56Y111_SLICE_X84Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y111_SLICE_X84Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y111_SLICE_X84Y111_CO5),
.O6(CLBLM_L_X56Y111_SLICE_X84Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y111_SLICE_X84Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y111_SLICE_X84Y111_BO5),
.O6(CLBLM_L_X56Y111_SLICE_X84Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0808000000000000)
  ) CLBLM_L_X56Y111_SLICE_X84Y111_ALUT (
.I0(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I1(CLBLL_R_X57Y102_SLICE_X86Y102_BQ),
.I2(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I3(1'b1),
.I4(CLBLL_R_X57Y102_SLICE_X86Y102_AQ),
.I5(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.O5(CLBLM_L_X56Y111_SLICE_X84Y111_AO5),
.O6(CLBLM_L_X56Y111_SLICE_X84Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y111_SLICE_X85Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y111_SLICE_X85Y111_DO5),
.O6(CLBLM_L_X56Y111_SLICE_X85Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y111_SLICE_X85Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y111_SLICE_X85Y111_CO5),
.O6(CLBLM_L_X56Y111_SLICE_X85Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y111_SLICE_X85Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y111_SLICE_X85Y111_BO5),
.O6(CLBLM_L_X56Y111_SLICE_X85Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y111_SLICE_X85Y111_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y111_SLICE_X85Y111_AO5),
.O6(CLBLM_L_X56Y111_SLICE_X85Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y96_SLICE_X90Y96_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_R_X57Y97_SLICE_X87Y97_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y96_SLICE_X89Y96_AQ),
.Q(CLBLM_L_X60Y96_SLICE_X90Y96_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y96_SLICE_X90Y96_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_R_X57Y97_SLICE_X87Y97_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y96_SLICE_X89Y96_A5Q),
.Q(CLBLM_L_X60Y96_SLICE_X90Y96_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y96_SLICE_X90Y96_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y96_SLICE_X90Y96_DO5),
.O6(CLBLM_L_X60Y96_SLICE_X90Y96_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y96_SLICE_X90Y96_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y96_SLICE_X90Y96_CO5),
.O6(CLBLM_L_X60Y96_SLICE_X90Y96_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y96_SLICE_X90Y96_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y96_SLICE_X90Y96_BO5),
.O6(CLBLM_L_X60Y96_SLICE_X90Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y96_SLICE_X90Y96_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y96_SLICE_X90Y96_AO5),
.O6(CLBLM_L_X60Y96_SLICE_X90Y96_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y96_SLICE_X91Y96_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y96_SLICE_X91Y96_DO5),
.O6(CLBLM_L_X60Y96_SLICE_X91Y96_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y96_SLICE_X91Y96_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y96_SLICE_X91Y96_CO5),
.O6(CLBLM_L_X60Y96_SLICE_X91Y96_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y96_SLICE_X91Y96_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y96_SLICE_X91Y96_BO5),
.O6(CLBLM_L_X60Y96_SLICE_X91Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y96_SLICE_X91Y96_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y96_SLICE_X91Y96_AO5),
.O6(CLBLM_L_X60Y96_SLICE_X91Y96_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X60Y97_SLICE_X90Y97_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y107_SLICE_X75Y107_DQ),
.Q(CLBLM_L_X60Y97_SLICE_X90Y97_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X60Y97_SLICE_X90Y97_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.D(CLBLM_L_X60Y97_SLICE_X90Y97_AO6),
.PRE(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.Q(CLBLM_L_X60Y97_SLICE_X90Y97_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X60Y97_SLICE_X90Y97_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.Q(CLBLM_L_X60Y97_SLICE_X90Y97_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X60Y97_SLICE_X90Y97_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X56Y97_SLICE_X84Y97_CO6),
.Q(CLBLM_L_X60Y97_SLICE_X90Y97_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33663366cc66cc66)
  ) CLBLM_L_X60Y97_SLICE_X90Y97_DLUT (
.I0(CLBLM_R_X59Y97_SLICE_X88Y97_BQ),
.I1(CLBLM_L_X60Y97_SLICE_X91Y97_AQ),
.I2(1'b1),
.I3(CLBLM_L_X60Y97_SLICE_X90Y97_A5Q),
.I4(1'b1),
.I5(CLBLL_R_X57Y97_SLICE_X86Y97_AQ),
.O5(CLBLM_L_X60Y97_SLICE_X90Y97_DO5),
.O6(CLBLM_L_X60Y97_SLICE_X90Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h665566aa665566aa)
  ) CLBLM_L_X60Y97_SLICE_X90Y97_CLUT (
.I0(CLBLM_L_X60Y97_SLICE_X91Y97_AQ),
.I1(CLBLM_R_X59Y96_SLICE_X88Y96_AQ),
.I2(1'b1),
.I3(CLBLM_L_X60Y97_SLICE_X90Y97_A5Q),
.I4(CLBLM_R_X59Y96_SLICE_X88Y96_BQ),
.I5(1'b1),
.O5(CLBLM_L_X60Y97_SLICE_X90Y97_CO5),
.O6(CLBLM_L_X60Y97_SLICE_X90Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffc)
  ) CLBLM_L_X60Y97_SLICE_X90Y97_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X50Y107_SLICE_X76Y107_BQ),
.I2(CLBLM_L_X60Y97_SLICE_X91Y97_AO6),
.I3(CLBLM_R_X49Y105_SLICE_X75Y105_CQ),
.I4(CLBLM_R_X49Y106_SLICE_X74Y106_AQ),
.I5(CLBLM_L_X50Y106_SLICE_X76Y106_CQ),
.O5(CLBLM_L_X60Y97_SLICE_X90Y97_BO5),
.O6(CLBLM_L_X60Y97_SLICE_X90Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h1313131313131313)
  ) CLBLM_L_X60Y97_SLICE_X90Y97_ALUT (
.I0(CLBLM_L_X56Y97_SLICE_X85Y97_DO6),
.I1(CLBLM_R_X63Y99_SLICE_X94Y99_DO5),
.I2(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y97_SLICE_X90Y97_AO5),
.O6(CLBLM_L_X60Y97_SLICE_X90Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X60Y97_SLICE_X91Y97_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y108_SLICE_X75Y108_DQ),
.Q(CLBLM_L_X60Y97_SLICE_X91Y97_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X60Y97_SLICE_X91Y97_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X60Y97_SLICE_X91Y97_BO6),
.Q(CLBLM_L_X60Y97_SLICE_X91Y97_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y97_SLICE_X91Y97_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y97_SLICE_X91Y97_DO5),
.O6(CLBLM_L_X60Y97_SLICE_X91Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y97_SLICE_X91Y97_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y97_SLICE_X91Y97_CO5),
.O6(CLBLM_L_X60Y97_SLICE_X91Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000000000)
  ) CLBLM_L_X60Y97_SLICE_X91Y97_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X63Y99_SLICE_X94Y99_DO5),
.I5(CLBLM_L_X62Y97_SLICE_X92Y97_CQ),
.O5(CLBLM_L_X60Y97_SLICE_X91Y97_BO5),
.O6(CLBLM_L_X60Y97_SLICE_X91Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefffeff000000)
  ) CLBLM_L_X60Y97_SLICE_X91Y97_ALUT (
.I0(CLBLM_L_X50Y106_SLICE_X76Y106_AQ),
.I1(CLBLM_L_X50Y104_SLICE_X76Y104_AQ),
.I2(CLBLM_L_X50Y105_SLICE_X77Y105_AQ),
.I3(CLBLM_L_X50Y107_SLICE_X77Y107_AQ),
.I4(CLBLM_L_X62Y100_SLICE_X92Y100_AO6),
.I5(1'b1),
.O5(CLBLM_L_X60Y97_SLICE_X91Y97_AO5),
.O6(CLBLM_L_X60Y97_SLICE_X91Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X60Y98_SLICE_X90Y98_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X60Y98_SLICE_X90Y98_AO6),
.Q(CLBLM_L_X60Y98_SLICE_X90Y98_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X60Y98_SLICE_X90Y98_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X60Y98_SLICE_X90Y98_BO6),
.Q(CLBLM_L_X60Y98_SLICE_X90Y98_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3733333305000000)
  ) CLBLM_L_X60Y98_SLICE_X90Y98_DLUT (
.I0(CLBLM_L_X60Y100_SLICE_X91Y100_CO5),
.I1(CLBLM_R_X53Y100_SLICE_X80Y100_AQ),
.I2(CLBLM_L_X62Y104_SLICE_X93Y104_AQ),
.I3(CLBLM_L_X60Y99_SLICE_X90Y99_AO6),
.I4(CLBLM_R_X59Y102_SLICE_X89Y102_AQ),
.I5(CLBLM_R_X53Y100_SLICE_X80Y100_A5Q),
.O5(CLBLM_L_X60Y98_SLICE_X90Y98_DO5),
.O6(CLBLM_L_X60Y98_SLICE_X90Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3c08000800)
  ) CLBLM_L_X60Y98_SLICE_X90Y98_CLUT (
.I0(CLBLM_R_X53Y100_SLICE_X80Y100_A5Q),
.I1(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I2(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I3(CLBLM_R_X53Y100_SLICE_X80Y100_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y98_SLICE_X90Y98_CO5),
.O6(CLBLM_L_X60Y98_SLICE_X90Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5c0c0c0c0c0c0c0c)
  ) CLBLM_L_X60Y98_SLICE_X90Y98_BLUT (
.I0(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I1(CLBLM_L_X60Y98_SLICE_X90Y98_BQ),
.I2(CLBLM_L_X62Y99_SLICE_X92Y99_AO6),
.I3(CLBLM_R_X53Y100_SLICE_X80Y100_A5Q),
.I4(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I5(CLBLM_R_X53Y100_SLICE_X80Y100_AQ),
.O5(CLBLM_L_X60Y98_SLICE_X90Y98_BO5),
.O6(CLBLM_L_X60Y98_SLICE_X90Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfff0f0cc00f0f0)
  ) CLBLM_L_X60Y98_SLICE_X90Y98_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X60Y97_SLICE_X90Y97_CO6),
.I2(CLBLM_L_X60Y98_SLICE_X90Y98_AQ),
.I3(CLBLM_L_X60Y97_SLICE_X90Y97_BQ),
.I4(CLBLM_L_X60Y98_SLICE_X91Y98_AQ),
.I5(CLBLM_L_X60Y97_SLICE_X90Y97_DO6),
.O5(CLBLM_L_X60Y98_SLICE_X90Y98_AO5),
.O6(CLBLM_L_X60Y98_SLICE_X90Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X60Y98_SLICE_X91Y98_A5_FDPE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y110_SLICE_X93Y110_BO6),
.D(CLBLM_L_X60Y98_SLICE_X90Y98_CO6),
.PRE(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.Q(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X60Y98_SLICE_X91Y98_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y110_SLICE_X93Y110_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X60Y98_SLICE_X91Y98_AO6),
.Q(CLBLM_L_X60Y98_SLICE_X91Y98_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X60Y98_SLICE_X91Y98_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y110_SLICE_X93Y110_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X60Y98_SLICE_X91Y98_AQ),
.Q(CLBLM_L_X60Y98_SLICE_X91Y98_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X60Y98_SLICE_X91Y98_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y110_SLICE_X93Y110_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X60Y98_SLICE_X91Y98_BQ),
.Q(CLBLM_L_X60Y98_SLICE_X91Y98_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X60Y98_SLICE_X91Y98_D_FDPE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y110_SLICE_X93Y110_BO6),
.D(CLBLM_L_X60Y98_SLICE_X91Y98_CQ),
.PRE(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.Q(CLBLM_L_X60Y98_SLICE_X91Y98_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y98_SLICE_X91Y98_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y98_SLICE_X91Y98_DO5),
.O6(CLBLM_L_X60Y98_SLICE_X91Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y98_SLICE_X91Y98_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y98_SLICE_X91Y98_CO5),
.O6(CLBLM_L_X60Y98_SLICE_X91Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y98_SLICE_X91Y98_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y98_SLICE_X91Y98_BO5),
.O6(CLBLM_L_X60Y98_SLICE_X91Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X60Y98_SLICE_X91Y98_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.O5(CLBLM_L_X60Y98_SLICE_X91Y98_AO5),
.O6(CLBLM_L_X60Y98_SLICE_X91Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y99_SLICE_X90Y99_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y99_SLICE_X92Y99_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X60Y99_SLICE_X90Y99_BO6),
.Q(CLBLM_L_X60Y99_SLICE_X90Y99_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y99_SLICE_X90Y99_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y99_SLICE_X92Y99_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X60Y99_SLICE_X90Y99_CO6),
.Q(CLBLM_L_X60Y99_SLICE_X90Y99_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f000f000f001f00)
  ) CLBLM_L_X60Y99_SLICE_X90Y99_DLUT (
.I0(CLBLM_L_X60Y100_SLICE_X91Y100_CO5),
.I1(CLBLM_L_X60Y100_SLICE_X91Y100_AO6),
.I2(CLBLM_R_X59Y100_SLICE_X88Y100_DO6),
.I3(CLBLM_L_X62Y99_SLICE_X92Y99_AO6),
.I4(CLBLM_R_X59Y102_SLICE_X89Y102_AQ),
.I5(CLBLM_L_X62Y104_SLICE_X93Y104_AQ),
.O5(CLBLM_L_X60Y99_SLICE_X90Y99_DO5),
.O6(CLBLM_L_X60Y99_SLICE_X90Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88ff00ff00ff00)
  ) CLBLM_L_X60Y99_SLICE_X90Y99_CLUT (
.I0(CLBLM_L_X62Y106_SLICE_X93Y106_AQ),
.I1(CLBLM_R_X63Y97_SLICE_X95Y97_F7AMUX_O),
.I2(1'b1),
.I3(CLBLM_R_X59Y102_SLICE_X88Y102_DO6),
.I4(CLBLM_R_X59Y102_SLICE_X89Y102_AQ),
.I5(CLBLM_L_X60Y110_SLICE_X91Y110_AQ),
.O5(CLBLM_L_X60Y99_SLICE_X90Y99_CO5),
.O6(CLBLM_L_X60Y99_SLICE_X90Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf780ff0088880000)
  ) CLBLM_L_X60Y99_SLICE_X90Y99_BLUT (
.I0(CLBLM_L_X60Y110_SLICE_X91Y110_AQ),
.I1(CLBLM_L_X62Y106_SLICE_X93Y106_AQ),
.I2(CLBLM_R_X63Y98_SLICE_X94Y98_F7AMUX_O),
.I3(CLBLM_R_X59Y103_SLICE_X88Y103_CO6),
.I4(CLBLM_R_X59Y102_SLICE_X89Y102_AQ),
.I5(1'b1),
.O5(CLBLM_L_X60Y99_SLICE_X90Y99_BO5),
.O6(CLBLM_L_X60Y99_SLICE_X90Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f000000010000)
  ) CLBLM_L_X60Y99_SLICE_X90Y99_ALUT (
.I0(CLBLM_R_X59Y102_SLICE_X89Y102_AQ),
.I1(CLBLM_L_X60Y99_SLICE_X91Y99_BO6),
.I2(CLBLM_R_X59Y102_SLICE_X88Y102_AQ),
.I3(CLBLM_L_X62Y104_SLICE_X93Y104_AQ),
.I4(CLBLM_L_X60Y98_SLICE_X90Y98_BQ),
.I5(1'b1),
.O5(CLBLM_L_X60Y99_SLICE_X90Y99_AO5),
.O6(CLBLM_L_X60Y99_SLICE_X90Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000001000)
  ) CLBLM_L_X60Y99_SLICE_X91Y99_DLUT (
.I0(CLBLM_R_X59Y102_SLICE_X88Y102_AQ),
.I1(CLBLM_L_X62Y111_SLICE_X92Y111_BO6),
.I2(CLBLM_R_X59Y102_SLICE_X89Y102_AQ),
.I3(CLBLM_L_X60Y98_SLICE_X90Y98_BQ),
.I4(CLBLM_L_X60Y99_SLICE_X91Y99_BO5),
.I5(CLBLM_L_X62Y104_SLICE_X93Y104_AQ),
.O5(CLBLM_L_X60Y99_SLICE_X91Y99_DO5),
.O6(CLBLM_L_X60Y99_SLICE_X91Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffd)
  ) CLBLM_L_X60Y99_SLICE_X91Y99_CLUT (
.I0(CLBLM_L_X62Y106_SLICE_X93Y106_AQ),
.I1(CLBLM_L_X62Y111_SLICE_X92Y111_BO6),
.I2(CLBLM_R_X59Y102_SLICE_X89Y102_AQ),
.I3(CLBLM_L_X62Y103_SLICE_X92Y103_AQ),
.I4(CLBLM_L_X60Y110_SLICE_X91Y110_AQ),
.I5(CLBLM_L_X62Y104_SLICE_X93Y104_AQ),
.O5(CLBLM_L_X60Y99_SLICE_X91Y99_CO5),
.O6(CLBLM_L_X60Y99_SLICE_X91Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7fff7ffffbbffbb)
  ) CLBLM_L_X60Y99_SLICE_X91Y99_BLUT (
.I0(CLBLM_L_X62Y103_SLICE_X92Y103_AQ),
.I1(CLBLM_L_X60Y110_SLICE_X91Y110_AQ),
.I2(CLBLM_L_X62Y110_SLICE_X92Y110_DO6),
.I3(CLBLM_L_X62Y106_SLICE_X93Y106_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y99_SLICE_X91Y99_BO5),
.O6(CLBLM_L_X60Y99_SLICE_X91Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff000000cc)
  ) CLBLM_L_X60Y99_SLICE_X91Y99_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X60Y98_SLICE_X90Y98_BQ),
.I2(1'b1),
.I3(CLBLM_R_X59Y102_SLICE_X88Y102_AQ),
.I4(CLBLM_L_X60Y99_SLICE_X91Y99_CO6),
.I5(1'b1),
.O5(CLBLM_L_X60Y99_SLICE_X91Y99_AO5),
.O6(CLBLM_L_X60Y99_SLICE_X91Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y100_SLICE_X90Y100_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y99_SLICE_X90Y99_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y100_SLICE_X88Y100_AO5),
.Q(CLBLM_L_X60Y100_SLICE_X90Y100_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h01000100ff00ff00)
  ) CLBLM_L_X60Y100_SLICE_X90Y100_DLUT (
.I0(CLBLM_R_X59Y102_SLICE_X89Y102_AQ),
.I1(CLBLM_L_X60Y100_SLICE_X91Y100_AO5),
.I2(CLBLM_L_X60Y100_SLICE_X91Y100_CO5),
.I3(CLBLM_L_X62Y99_SLICE_X92Y99_AO6),
.I4(1'b1),
.I5(CLBLM_R_X59Y100_SLICE_X88Y100_DO6),
.O5(CLBLM_L_X60Y100_SLICE_X90Y100_DO5),
.O6(CLBLM_L_X60Y100_SLICE_X90Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f000f002f002f00)
  ) CLBLM_L_X60Y100_SLICE_X90Y100_CLUT (
.I0(CLBLM_R_X59Y102_SLICE_X89Y102_AQ),
.I1(CLBLM_L_X60Y100_SLICE_X91Y100_AO5),
.I2(CLBLM_R_X59Y101_SLICE_X88Y101_AO6),
.I3(CLBLM_L_X62Y99_SLICE_X92Y99_AO6),
.I4(1'b1),
.I5(CLBLM_L_X60Y100_SLICE_X91Y100_CO5),
.O5(CLBLM_L_X60Y100_SLICE_X90Y100_CO5),
.O6(CLBLM_L_X60Y100_SLICE_X90Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h44444444444c4444)
  ) CLBLM_L_X60Y100_SLICE_X90Y100_BLUT (
.I0(CLBLM_R_X59Y101_SLICE_X88Y101_AO6),
.I1(CLBLM_L_X62Y99_SLICE_X92Y99_AO6),
.I2(CLBLM_L_X60Y100_SLICE_X91Y100_AO6),
.I3(CLBLM_L_X60Y100_SLICE_X91Y100_CO5),
.I4(CLBLM_R_X59Y102_SLICE_X89Y102_AQ),
.I5(CLBLM_L_X62Y104_SLICE_X93Y104_AQ),
.O5(CLBLM_L_X60Y100_SLICE_X90Y100_BO5),
.O6(CLBLM_L_X60Y100_SLICE_X90Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0ccaaffaa00)
  ) CLBLM_L_X60Y100_SLICE_X90Y100_ALUT (
.I0(CLBLM_L_X60Y99_SLICE_X90Y99_CQ),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(CLBLM_L_X60Y99_SLICE_X90Y99_AQ),
.I3(CLBLM_L_X62Y99_SLICE_X92Y99_BQ),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(1'b1),
.O5(CLBLM_L_X60Y100_SLICE_X90Y100_AO5),
.O6(CLBLM_L_X60Y100_SLICE_X90Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y100_SLICE_X91Y100_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y99_SLICE_X92Y99_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X60Y100_SLICE_X91Y100_BO6),
.Q(CLBLM_L_X60Y100_SLICE_X91Y100_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf053f053ff53ff53)
  ) CLBLM_L_X60Y100_SLICE_X91Y100_DLUT (
.I0(CLBLM_R_X59Y97_SLICE_X88Y97_BQ),
.I1(CLBLM_L_X62Y107_SLICE_X92Y107_AQ),
.I2(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I3(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I4(1'b1),
.I5(CLBLM_L_X62Y104_SLICE_X92Y104_AQ),
.O5(CLBLM_L_X60Y100_SLICE_X91Y100_DO5),
.O6(CLBLM_L_X60Y100_SLICE_X91Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefffefffffbfffb)
  ) CLBLM_L_X60Y100_SLICE_X91Y100_CLUT (
.I0(CLBLM_L_X62Y103_SLICE_X92Y103_AQ),
.I1(CLBLM_L_X62Y106_SLICE_X93Y106_AQ),
.I2(CLBLM_L_X62Y110_SLICE_X92Y110_DO6),
.I3(CLBLM_L_X60Y110_SLICE_X91Y110_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y100_SLICE_X91Y100_CO5),
.O6(CLBLM_L_X60Y100_SLICE_X91Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcaaacaaaaaaaaaaa)
  ) CLBLM_L_X60Y100_SLICE_X91Y100_BLUT (
.I0(CLBLM_L_X60Y101_SLICE_X91Y101_DO6),
.I1(CLBLM_R_X63Y99_SLICE_X94Y99_F7AMUX_O),
.I2(CLBLM_R_X59Y102_SLICE_X89Y102_AQ),
.I3(CLBLM_L_X60Y110_SLICE_X91Y110_AQ),
.I4(1'b1),
.I5(CLBLM_L_X62Y106_SLICE_X93Y106_AQ),
.O5(CLBLM_L_X60Y100_SLICE_X91Y100_BO5),
.O6(CLBLM_L_X60Y100_SLICE_X91Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff7fffdfffffff)
  ) CLBLM_L_X60Y100_SLICE_X91Y100_ALUT (
.I0(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I1(CLBLM_R_X59Y102_SLICE_X88Y102_AQ),
.I2(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I3(CLBLM_L_X60Y98_SLICE_X90Y98_BQ),
.I4(CLBLM_L_X62Y104_SLICE_X93Y104_AQ),
.I5(1'b1),
.O5(CLBLM_L_X60Y100_SLICE_X91Y100_AO5),
.O6(CLBLM_L_X60Y100_SLICE_X91Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y101_SLICE_X90Y101_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y102_SLICE_X92Y102_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X60Y101_SLICE_X90Y101_AO6),
.Q(CLBLM_L_X60Y101_SLICE_X90Y101_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaccaaaaaaaaaa)
  ) CLBLM_L_X60Y101_SLICE_X90Y101_DLUT (
.I0(CLBLM_R_X59Y104_SLICE_X89Y104_CQ),
.I1(CLBLM_L_X60Y105_SLICE_X90Y105_D_XOR),
.I2(1'b1),
.I3(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I4(1'b1),
.I5(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.O5(CLBLM_L_X60Y101_SLICE_X90Y101_DO5),
.O6(CLBLM_L_X60Y101_SLICE_X90Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00ffff0000)
  ) CLBLM_L_X60Y101_SLICE_X90Y101_CLUT (
.I0(CLBLM_L_X60Y105_SLICE_X90Y105_C_XOR),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I4(CLBLM_R_X59Y105_SLICE_X89Y105_CQ),
.I5(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.O5(CLBLM_L_X60Y101_SLICE_X90Y101_CO5),
.O6(CLBLM_L_X60Y101_SLICE_X90Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00bf00ff00)
  ) CLBLM_L_X60Y101_SLICE_X90Y101_BLUT (
.I0(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I1(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I2(CLBLL_L_X54Y101_SLICE_X83Y101_AO6),
.I3(CLBLM_R_X59Y101_SLICE_X89Y101_BO6),
.I4(CLBLM_L_X64Y100_SLICE_X97Y100_BQ),
.I5(CLBLM_L_X64Y100_SLICE_X97Y100_AQ),
.O5(CLBLM_L_X60Y101_SLICE_X90Y101_BO5),
.O6(CLBLM_L_X60Y101_SLICE_X90Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffec3320dfcc1300)
  ) CLBLM_L_X60Y101_SLICE_X90Y101_ALUT (
.I0(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I1(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I2(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I3(CLBLM_L_X60Y106_SLICE_X91Y106_D_XOR),
.I4(CLBLM_L_X62Y97_SLICE_X92Y97_AO6),
.I5(CLBLM_L_X60Y103_SLICE_X91Y103_D_XOR),
.O5(CLBLM_L_X60Y101_SLICE_X90Y101_AO5),
.O6(CLBLM_L_X60Y101_SLICE_X90Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y101_SLICE_X91Y101_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y99_SLICE_X92Y99_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X60Y101_SLICE_X91Y101_AO6),
.Q(CLBLM_L_X60Y101_SLICE_X91Y101_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y101_SLICE_X91Y101_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y99_SLICE_X92Y99_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X60Y101_SLICE_X91Y101_BO6),
.Q(CLBLM_L_X60Y101_SLICE_X91Y101_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h440c770c443f773f)
  ) CLBLM_L_X60Y101_SLICE_X91Y101_DLUT (
.I0(CLBLL_R_X57Y104_SLICE_X87Y104_DO6),
.I1(CLBLM_L_X62Y103_SLICE_X93Y103_BO6),
.I2(CLBLM_L_X64Y105_SLICE_X96Y105_DO6),
.I3(CLBLM_L_X62Y106_SLICE_X93Y106_CO6),
.I4(CLBLM_L_X60Y100_SLICE_X91Y100_DO6),
.I5(CLBLM_R_X59Y101_SLICE_X89Y101_CO6),
.O5(CLBLM_L_X60Y101_SLICE_X91Y101_DO5),
.O6(CLBLM_L_X60Y101_SLICE_X91Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88fafa5050)
  ) CLBLM_L_X60Y101_SLICE_X91Y101_CLUT (
.I0(CLBLM_L_X62Y99_SLICE_X92Y99_BQ),
.I1(CLBLM_L_X60Y100_SLICE_X91Y100_BQ),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(CLBLM_L_X60Y101_SLICE_X91Y101_AQ),
.I5(1'b1),
.O5(CLBLM_L_X60Y101_SLICE_X91Y101_CO5),
.O6(CLBLM_L_X60Y101_SLICE_X91Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeebbaa55441100)
  ) CLBLM_L_X60Y101_SLICE_X91Y101_BLUT (
.I0(CLBLM_L_X60Y99_SLICE_X90Y99_BO5),
.I1(CLBLM_L_X62Y103_SLICE_X93Y103_BO6),
.I2(1'b1),
.I3(CLBLM_L_X62Y105_SLICE_X92Y105_DO6),
.I4(CLBLM_R_X59Y105_SLICE_X89Y105_F7AMUX_O),
.I5(CLBLM_L_X62Y97_SLICE_X93Y97_F7AMUX_O),
.O5(CLBLM_L_X60Y101_SLICE_X91Y101_BO5),
.O6(CLBLM_L_X60Y101_SLICE_X91Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500ffaa7722)
  ) CLBLM_L_X60Y101_SLICE_X91Y101_ALUT (
.I0(CLBLM_L_X60Y99_SLICE_X90Y99_BO5),
.I1(CLBLM_R_X63Y96_SLICE_X95Y96_CO6),
.I2(1'b1),
.I3(CLBLM_R_X59Y102_SLICE_X89Y102_BO6),
.I4(CLBLM_R_X63Y101_SLICE_X95Y101_BO6),
.I5(CLBLM_L_X62Y106_SLICE_X93Y106_CO6),
.O5(CLBLM_L_X60Y101_SLICE_X91Y101_AO5),
.O6(CLBLM_L_X60Y101_SLICE_X91Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y102_SLICE_X90Y102_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y102_SLICE_X92Y102_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X60Y102_SLICE_X90Y102_AO6),
.Q(CLBLM_L_X60Y102_SLICE_X90Y102_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y102_SLICE_X90Y102_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y102_SLICE_X92Y102_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X60Y102_SLICE_X90Y102_BO6),
.Q(CLBLM_L_X60Y102_SLICE_X90Y102_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y102_SLICE_X90Y102_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y102_SLICE_X92Y102_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X60Y102_SLICE_X90Y102_CO6),
.Q(CLBLM_L_X60Y102_SLICE_X90Y102_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe02fffffe020000)
  ) CLBLM_L_X60Y102_SLICE_X90Y102_DLUT (
.I0(CLBLM_L_X60Y105_SLICE_X91Y105_C_XOR),
.I1(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I2(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I3(CLBLM_L_X60Y102_SLICE_X90Y102_AQ),
.I4(CLBLM_R_X59Y103_SLICE_X89Y103_CQ),
.I5(CLBLM_L_X60Y101_SLICE_X90Y101_DO6),
.O5(CLBLM_L_X60Y102_SLICE_X90Y102_DO5),
.O6(CLBLM_L_X60Y102_SLICE_X90Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ffffdf80)
  ) CLBLM_L_X60Y102_SLICE_X90Y102_CLUT (
.I0(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I1(CLBLM_L_X60Y102_SLICE_X91Y102_A_XOR),
.I2(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I3(CLBLM_L_X60Y105_SLICE_X91Y105_A_XOR),
.I4(CLBLM_L_X62Y103_SLICE_X93Y103_AO6),
.I5(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.O5(CLBLM_L_X60Y102_SLICE_X90Y102_CO5),
.O6(CLBLM_L_X60Y102_SLICE_X90Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0fdf8fff0)
  ) CLBLM_L_X60Y102_SLICE_X90Y102_BLUT (
.I0(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I1(CLBLM_L_X60Y102_SLICE_X91Y102_D_XOR),
.I2(CLBLM_L_X62Y102_SLICE_X92Y102_AO5),
.I3(CLBLM_L_X60Y105_SLICE_X91Y105_D_XOR),
.I4(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I5(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.O5(CLBLM_L_X60Y102_SLICE_X90Y102_BO5),
.O6(CLBLM_L_X60Y102_SLICE_X90Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00e400cc)
  ) CLBLM_L_X60Y102_SLICE_X90Y102_ALUT (
.I0(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I1(CLBLM_L_X60Y105_SLICE_X91Y105_C_XOR),
.I2(CLBLM_L_X60Y102_SLICE_X91Y102_C_XOR),
.I3(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I4(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I5(CLBLM_L_X62Y98_SLICE_X92Y98_AO6),
.O5(CLBLM_L_X60Y102_SLICE_X90Y102_AO5),
.O6(CLBLM_L_X60Y102_SLICE_X90Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y102_SLICE_X91Y102_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y102_SLICE_X92Y102_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X60Y102_SLICE_X91Y102_BO5),
.Q(CLBLM_L_X60Y102_SLICE_X91Y102_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X60Y102_SLICE_X91Y102_CARRY4 (
.CI(1'b0),
.CO({CLBLM_L_X60Y102_SLICE_X91Y102_D_CY, CLBLM_L_X60Y102_SLICE_X91Y102_C_CY, CLBLM_L_X60Y102_SLICE_X91Y102_B_CY, CLBLM_L_X60Y102_SLICE_X91Y102_A_CY}),
.CYINIT(CLBLM_L_X62Y102_SLICE_X92Y102_BQ),
.DI({CLBLM_L_X60Y102_SLICE_X90Y102_BQ, CLBLM_L_X60Y102_SLICE_X90Y102_AQ, CLBLM_L_X62Y104_SLICE_X92Y104_AQ, CLBLM_L_X60Y102_SLICE_X91Y102_AO5}),
.O({CLBLM_L_X60Y102_SLICE_X91Y102_D_XOR, CLBLM_L_X60Y102_SLICE_X91Y102_C_XOR, CLBLM_L_X60Y102_SLICE_X91Y102_B_XOR, CLBLM_L_X60Y102_SLICE_X91Y102_A_XOR}),
.S({CLBLM_L_X60Y102_SLICE_X91Y102_DO6, CLBLM_L_X60Y102_SLICE_X91Y102_CO6, CLBLM_L_X60Y102_SLICE_X91Y102_BO6, CLBLM_L_X60Y102_SLICE_X91Y102_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffffffff)
  ) CLBLM_L_X60Y102_SLICE_X91Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X60Y102_SLICE_X90Y102_BQ),
.O5(CLBLM_L_X60Y102_SLICE_X91Y102_DO5),
.O6(CLBLM_L_X60Y102_SLICE_X91Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555555)
  ) CLBLM_L_X60Y102_SLICE_X91Y102_CLUT (
.I0(CLBLM_L_X60Y102_SLICE_X90Y102_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y102_SLICE_X91Y102_CO5),
.O6(CLBLM_L_X60Y102_SLICE_X91Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333333ff00ff00)
  ) CLBLM_L_X60Y102_SLICE_X91Y102_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X62Y104_SLICE_X92Y104_AQ),
.I2(1'b1),
.I3(CLBLM_L_X62Y102_SLICE_X92Y102_AO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y102_SLICE_X91Y102_BO5),
.O6(CLBLM_L_X60Y102_SLICE_X91Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333333cccccccc)
  ) CLBLM_L_X60Y102_SLICE_X91Y102_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X60Y102_SLICE_X90Y102_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y102_SLICE_X91Y102_AO5),
.O6(CLBLM_L_X60Y102_SLICE_X91Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacaff0fcacaf000)
  ) CLBLM_L_X60Y103_SLICE_X90Y103_DLUT (
.I0(CLBLM_L_X60Y103_SLICE_X91Y103_AQ),
.I1(CLBLM_R_X59Y98_SLICE_X88Y98_CQ),
.I2(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I3(CLBLM_L_X60Y104_SLICE_X90Y104_AQ),
.I4(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I5(CLBLM_R_X59Y98_SLICE_X89Y98_CQ),
.O5(CLBLM_L_X60Y103_SLICE_X90Y103_DO5),
.O6(CLBLM_L_X60Y103_SLICE_X90Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fafa00000afa0)
  ) CLBLM_L_X60Y103_SLICE_X90Y103_CLUT (
.I0(CLBLM_R_X59Y96_SLICE_X88Y96_AQ),
.I1(1'b1),
.I2(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I3(CLBLM_L_X60Y102_SLICE_X91Y102_BQ),
.I4(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I5(CLBLM_L_X60Y102_SLICE_X90Y102_BQ),
.O5(CLBLM_L_X60Y103_SLICE_X90Y103_CO5),
.O6(CLBLM_L_X60Y103_SLICE_X90Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55e455e400e400e4)
  ) CLBLM_L_X60Y103_SLICE_X90Y103_BLUT (
.I0(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I1(CLBLM_L_X64Y108_SLICE_X96Y108_AQ),
.I2(CLBLM_R_X49Y109_SLICE_X74Y109_AQ),
.I3(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I4(1'b1),
.I5(CLBLM_R_X63Y104_SLICE_X94Y104_BQ),
.O5(CLBLM_L_X60Y103_SLICE_X90Y103_BO5),
.O6(CLBLM_L_X60Y103_SLICE_X90Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heef5eea044f544a0)
  ) CLBLM_L_X60Y103_SLICE_X90Y103_ALUT (
.I0(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I1(CLBLM_L_X56Y103_SLICE_X85Y103_BQ),
.I2(CLBLM_L_X60Y104_SLICE_X91Y104_AQ),
.I3(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I4(CLBLM_L_X56Y103_SLICE_X85Y103_AQ),
.I5(CLBLL_R_X57Y103_SLICE_X87Y103_AQ),
.O5(CLBLM_L_X60Y103_SLICE_X90Y103_AO5),
.O6(CLBLM_L_X60Y103_SLICE_X90Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X60Y103_SLICE_X90Y103_MUXF7A (
.I0(CLBLM_L_X60Y103_SLICE_X90Y103_BO6),
.I1(CLBLM_L_X60Y103_SLICE_X90Y103_AO6),
.O(CLBLM_L_X60Y103_SLICE_X90Y103_F7AMUX_O),
.S(CLBLM_L_X62Y106_SLICE_X93Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X60Y103_SLICE_X90Y103_MUXF7B (
.I0(CLBLM_L_X60Y103_SLICE_X90Y103_DO6),
.I1(CLBLM_L_X60Y103_SLICE_X90Y103_CO6),
.O(CLBLM_L_X60Y103_SLICE_X90Y103_F7BMUX_O),
.S(CLBLM_L_X62Y106_SLICE_X93Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLM_L_X60Y103_SLICE_X90Y103_MUXF8 (
.I0(CLBLM_L_X60Y103_SLICE_X90Y103_F7BMUX_O),
.I1(CLBLM_L_X60Y103_SLICE_X90Y103_F7AMUX_O),
.O(CLBLM_L_X60Y103_SLICE_X90Y103_F8MUX_O),
.S(CLBLM_L_X62Y103_SLICE_X93Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y103_SLICE_X91Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y100_SLICE_X90Y100_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X60Y103_SLICE_X91Y103_AO5),
.Q(CLBLM_L_X60Y103_SLICE_X91Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X60Y103_SLICE_X91Y103_CARRY4 (
.CI(CLBLM_L_X60Y102_SLICE_X91Y102_COUT),
.CO({CLBLM_L_X60Y103_SLICE_X91Y103_D_CY, CLBLM_L_X60Y103_SLICE_X91Y103_C_CY, CLBLM_L_X60Y103_SLICE_X91Y103_B_CY, CLBLM_L_X60Y103_SLICE_X91Y103_A_CY}),
.CYINIT(1'b0),
.DI({CLBLM_L_X60Y101_SLICE_X90Y101_AQ, CLBLM_L_X62Y106_SLICE_X92Y106_CQ, CLBLM_L_X62Y106_SLICE_X92Y106_BQ, CLBLM_L_X62Y104_SLICE_X92Y104_BQ}),
.O({CLBLM_L_X60Y103_SLICE_X91Y103_D_XOR, CLBLM_L_X60Y103_SLICE_X91Y103_C_XOR, CLBLM_L_X60Y103_SLICE_X91Y103_B_XOR, CLBLM_L_X60Y103_SLICE_X91Y103_A_XOR}),
.S({CLBLM_L_X60Y103_SLICE_X91Y103_DO6, CLBLM_L_X60Y103_SLICE_X91Y103_CO6, CLBLM_L_X60Y103_SLICE_X91Y103_BO6, CLBLM_L_X60Y103_SLICE_X91Y103_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffff0000ffff)
  ) CLBLM_L_X60Y103_SLICE_X91Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X60Y101_SLICE_X90Y101_AQ),
.I5(1'b1),
.O5(CLBLM_L_X60Y103_SLICE_X91Y103_DO5),
.O6(CLBLM_L_X60Y103_SLICE_X91Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0f0f0f)
  ) CLBLM_L_X60Y103_SLICE_X91Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X62Y106_SLICE_X92Y106_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y103_SLICE_X91Y103_CO5),
.O6(CLBLM_L_X60Y103_SLICE_X91Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffffffff)
  ) CLBLM_L_X60Y103_SLICE_X91Y103_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X62Y106_SLICE_X92Y106_BQ),
.O5(CLBLM_L_X60Y103_SLICE_X91Y103_BO5),
.O6(CLBLM_L_X60Y103_SLICE_X91Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333333f0f0f0f0)
  ) CLBLM_L_X60Y103_SLICE_X91Y103_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X62Y104_SLICE_X92Y104_BQ),
.I2(CLBLM_L_X62Y102_SLICE_X92Y102_AO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y103_SLICE_X91Y103_AO5),
.O6(CLBLM_L_X60Y103_SLICE_X91Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y104_SLICE_X90Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y99_SLICE_X90Y99_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X60Y104_SLICE_X90Y104_AO6),
.Q(CLBLM_L_X60Y104_SLICE_X90Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5ffa000f5ffa000)
  ) CLBLM_L_X60Y104_SLICE_X90Y104_DLUT (
.I0(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I1(1'b1),
.I2(CLBLM_L_X60Y105_SLICE_X90Y105_B_XOR),
.I3(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I4(CLBLM_R_X59Y106_SLICE_X89Y106_CQ),
.I5(1'b1),
.O5(CLBLM_L_X60Y104_SLICE_X90Y104_DO5),
.O6(CLBLM_L_X60Y104_SLICE_X90Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h11dd030311ddcfcf)
  ) CLBLM_L_X60Y104_SLICE_X90Y104_CLUT (
.I0(CLBLM_L_X60Y106_SLICE_X90Y106_AQ),
.I1(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I2(CLBLM_R_X59Y98_SLICE_X89Y98_C5Q),
.I3(CLBLM_R_X59Y100_SLICE_X89Y100_BQ),
.I4(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I5(CLBLM_R_X59Y112_SLICE_X89Y112_AQ),
.O5(CLBLM_L_X60Y104_SLICE_X90Y104_CO5),
.O6(CLBLM_L_X60Y104_SLICE_X90Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff03aaaafc00aaaa)
  ) CLBLM_L_X60Y104_SLICE_X90Y104_BLUT (
.I0(CLBLM_L_X60Y104_SLICE_X90Y104_DO6),
.I1(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I2(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I3(CLBLM_L_X60Y102_SLICE_X90Y102_CQ),
.I4(CLBLM_R_X59Y103_SLICE_X89Y103_CQ),
.I5(CLBLM_L_X60Y105_SLICE_X91Y105_A_XOR),
.O5(CLBLM_L_X60Y104_SLICE_X90Y104_BO5),
.O6(CLBLM_L_X60Y104_SLICE_X90Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff54ff55ff04ff00)
  ) CLBLM_L_X60Y104_SLICE_X90Y104_ALUT (
.I0(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I1(CLBLM_R_X59Y107_SLICE_X89Y107_D_XOR),
.I2(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I3(CLBLM_L_X62Y102_SLICE_X92Y102_AO5),
.I4(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I5(CLBLM_L_X60Y108_SLICE_X90Y108_D_XOR),
.O5(CLBLM_L_X60Y104_SLICE_X90Y104_AO5),
.O6(CLBLM_L_X60Y104_SLICE_X90Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y104_SLICE_X91Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y100_SLICE_X90Y100_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X60Y104_SLICE_X91Y104_AO5),
.Q(CLBLM_L_X60Y104_SLICE_X91Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X60Y104_SLICE_X91Y104_CARRY4 (
.CI(CLBLM_L_X60Y103_SLICE_X91Y103_COUT),
.CO({CLBLM_L_X60Y104_SLICE_X91Y104_D_CY, CLBLM_L_X60Y104_SLICE_X91Y104_C_CY, CLBLM_L_X60Y104_SLICE_X91Y104_B_CY, CLBLM_L_X60Y104_SLICE_X91Y104_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, CLBLM_L_X62Y107_SLICE_X92Y107_AQ, CLBLM_L_X60Y109_SLICE_X91Y109_AQ}),
.O({CLBLM_L_X60Y104_SLICE_X91Y104_D_XOR, CLBLM_L_X60Y104_SLICE_X91Y104_C_XOR, CLBLM_L_X60Y104_SLICE_X91Y104_B_XOR, CLBLM_L_X60Y104_SLICE_X91Y104_A_XOR}),
.S({CLBLM_L_X60Y104_SLICE_X91Y104_DO6, CLBLM_L_X60Y104_SLICE_X91Y104_CO6, CLBLM_L_X60Y104_SLICE_X91Y104_BO6, CLBLM_L_X60Y104_SLICE_X91Y104_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y104_SLICE_X91Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y104_SLICE_X91Y104_DO5),
.O6(CLBLM_L_X60Y104_SLICE_X91Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00ff00ff)
  ) CLBLM_L_X60Y104_SLICE_X91Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X60Y109_SLICE_X91Y109_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y104_SLICE_X91Y104_CO5),
.O6(CLBLM_L_X60Y104_SLICE_X91Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffff0000ffff)
  ) CLBLM_L_X60Y104_SLICE_X91Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X62Y107_SLICE_X92Y107_AQ),
.I5(1'b1),
.O5(CLBLM_L_X60Y104_SLICE_X91Y104_BO5),
.O6(CLBLM_L_X60Y104_SLICE_X91Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00fff0f0f0f0)
  ) CLBLM_L_X60Y104_SLICE_X91Y104_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X62Y102_SLICE_X92Y102_AO6),
.I3(CLBLM_L_X60Y109_SLICE_X91Y109_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y104_SLICE_X91Y104_AO5),
.O6(CLBLM_L_X60Y104_SLICE_X91Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X60Y105_SLICE_X90Y105_CARRY4 (
.CI(1'b0),
.CO({CLBLM_L_X60Y105_SLICE_X90Y105_D_CY, CLBLM_L_X60Y105_SLICE_X90Y105_C_CY, CLBLM_L_X60Y105_SLICE_X90Y105_B_CY, CLBLM_L_X60Y105_SLICE_X90Y105_A_CY}),
.CYINIT(1'b0),
.DI({CLBLM_L_X60Y102_SLICE_X90Y102_AQ, CLBLM_L_X62Y104_SLICE_X92Y104_AQ, CLBLM_L_X60Y102_SLICE_X90Y102_CQ, CLBLM_L_X62Y102_SLICE_X92Y102_BQ}),
.O({CLBLM_L_X60Y105_SLICE_X90Y105_D_XOR, CLBLM_L_X60Y105_SLICE_X90Y105_C_XOR, CLBLM_L_X60Y105_SLICE_X90Y105_B_XOR, CLBLM_L_X60Y105_SLICE_X90Y105_A_XOR}),
.S({CLBLM_L_X60Y105_SLICE_X90Y105_DO6, CLBLM_L_X60Y105_SLICE_X90Y105_CO6, CLBLM_L_X60Y105_SLICE_X90Y105_BO6, CLBLM_L_X60Y105_SLICE_X90Y105_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ffff00ff00)
  ) CLBLM_L_X60Y105_SLICE_X90Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X59Y98_SLICE_X89Y98_B5Q),
.I4(1'b1),
.I5(CLBLM_L_X60Y102_SLICE_X90Y102_AQ),
.O5(CLBLM_L_X60Y105_SLICE_X90Y105_DO5),
.O6(CLBLM_L_X60Y105_SLICE_X90Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6666666666666666)
  ) CLBLM_L_X60Y105_SLICE_X90Y105_CLUT (
.I0(CLBLM_R_X59Y98_SLICE_X89Y98_BQ),
.I1(CLBLM_L_X62Y104_SLICE_X92Y104_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y105_SLICE_X90Y105_CO5),
.O6(CLBLM_L_X60Y105_SLICE_X90Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0ff0f0f0f0)
  ) CLBLM_L_X60Y105_SLICE_X90Y105_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X60Y102_SLICE_X90Y102_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X59Y98_SLICE_X89Y98_A5Q),
.O5(CLBLM_L_X60Y105_SLICE_X90Y105_BO5),
.O6(CLBLM_L_X60Y105_SLICE_X90Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff00ff00ff00ff0)
  ) CLBLM_L_X60Y105_SLICE_X90Y105_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X62Y102_SLICE_X92Y102_BQ),
.I3(CLBLM_R_X59Y98_SLICE_X89Y98_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y105_SLICE_X90Y105_AO5),
.O6(CLBLM_L_X60Y105_SLICE_X90Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X60Y105_SLICE_X91Y105_CARRY4 (
.CI(1'b0),
.CO({CLBLM_L_X60Y105_SLICE_X91Y105_D_CY, CLBLM_L_X60Y105_SLICE_X91Y105_C_CY, CLBLM_L_X60Y105_SLICE_X91Y105_B_CY, CLBLM_L_X60Y105_SLICE_X91Y105_A_CY}),
.CYINIT(CLBLM_L_X62Y102_SLICE_X92Y102_BQ),
.DI({1'b0, 1'b0, 1'b0, CLBLM_L_X60Y105_SLICE_X91Y105_AO5}),
.O({CLBLM_L_X60Y105_SLICE_X91Y105_D_XOR, CLBLM_L_X60Y105_SLICE_X91Y105_C_XOR, CLBLM_L_X60Y105_SLICE_X91Y105_B_XOR, CLBLM_L_X60Y105_SLICE_X91Y105_A_XOR}),
.S({CLBLM_L_X60Y105_SLICE_X91Y105_DO6, CLBLM_L_X60Y105_SLICE_X91Y105_CO6, CLBLM_L_X60Y105_SLICE_X91Y105_BO6, CLBLM_L_X60Y105_SLICE_X91Y105_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X60Y105_SLICE_X91Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X60Y102_SLICE_X90Y102_BQ),
.O5(CLBLM_L_X60Y105_SLICE_X91Y105_DO5),
.O6(CLBLM_L_X60Y105_SLICE_X91Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X60Y105_SLICE_X91Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X60Y102_SLICE_X90Y102_AQ),
.O5(CLBLM_L_X60Y105_SLICE_X91Y105_CO5),
.O6(CLBLM_L_X60Y105_SLICE_X91Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X60Y105_SLICE_X91Y105_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X62Y104_SLICE_X92Y104_AQ),
.O5(CLBLM_L_X60Y105_SLICE_X91Y105_BO5),
.O6(CLBLM_L_X60Y105_SLICE_X91Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0000000000)
  ) CLBLM_L_X60Y105_SLICE_X91Y105_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X60Y102_SLICE_X90Y102_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y105_SLICE_X91Y105_AO5),
.O6(CLBLM_L_X60Y105_SLICE_X91Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y106_SLICE_X90Y106_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y100_SLICE_X90Y100_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X60Y106_SLICE_X90Y106_AO5),
.Q(CLBLM_L_X60Y106_SLICE_X90Y106_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X60Y106_SLICE_X90Y106_CARRY4 (
.CI(CLBLM_L_X60Y105_SLICE_X90Y105_COUT),
.CO({CLBLM_L_X60Y106_SLICE_X90Y106_D_CY, CLBLM_L_X60Y106_SLICE_X90Y106_C_CY, CLBLM_L_X60Y106_SLICE_X90Y106_B_CY, CLBLM_L_X60Y106_SLICE_X90Y106_A_CY}),
.CYINIT(1'b0),
.DI({CLBLM_L_X62Y106_SLICE_X92Y106_CQ, CLBLM_L_X62Y106_SLICE_X92Y106_BQ, CLBLM_L_X62Y104_SLICE_X92Y104_BQ, CLBLM_L_X60Y102_SLICE_X90Y102_BQ}),
.O({CLBLM_L_X60Y106_SLICE_X90Y106_D_XOR, CLBLM_L_X60Y106_SLICE_X90Y106_C_XOR, CLBLM_L_X60Y106_SLICE_X90Y106_B_XOR, CLBLM_L_X60Y106_SLICE_X90Y106_A_XOR}),
.S({CLBLM_L_X60Y106_SLICE_X90Y106_DO6, CLBLM_L_X60Y106_SLICE_X90Y106_CO6, CLBLM_L_X60Y106_SLICE_X90Y106_BO6, CLBLM_L_X60Y106_SLICE_X90Y106_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0ff0f0f0f0)
  ) CLBLM_L_X60Y106_SLICE_X90Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X62Y106_SLICE_X92Y106_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X59Y96_SLICE_X89Y96_A5Q),
.O5(CLBLM_L_X60Y106_SLICE_X90Y106_DO5),
.O6(CLBLM_L_X60Y106_SLICE_X90Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff00ff00ff00ff0)
  ) CLBLM_L_X60Y106_SLICE_X90Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X59Y96_SLICE_X89Y96_AQ),
.I3(CLBLM_L_X62Y106_SLICE_X92Y106_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y106_SLICE_X90Y106_CO5),
.O6(CLBLM_L_X60Y106_SLICE_X90Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5a5a5a5a5a)
  ) CLBLM_L_X60Y106_SLICE_X90Y106_BLUT (
.I0(CLBLM_L_X62Y104_SLICE_X92Y104_BQ),
.I1(1'b1),
.I2(CLBLM_R_X59Y98_SLICE_X89Y98_C5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y106_SLICE_X90Y106_BO5),
.O6(CLBLM_L_X60Y106_SLICE_X90Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ccccff00ff00)
  ) CLBLM_L_X60Y106_SLICE_X90Y106_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X59Y98_SLICE_X89Y98_CQ),
.I2(1'b1),
.I3(CLBLM_L_X62Y106_SLICE_X93Y106_BO6),
.I4(CLBLM_L_X60Y102_SLICE_X90Y102_BQ),
.I5(1'b1),
.O5(CLBLM_L_X60Y106_SLICE_X90Y106_AO5),
.O6(CLBLM_L_X60Y106_SLICE_X90Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X60Y106_SLICE_X91Y106_CARRY4 (
.CI(CLBLM_L_X60Y105_SLICE_X91Y105_COUT),
.CO({CLBLM_L_X60Y106_SLICE_X91Y106_D_CY, CLBLM_L_X60Y106_SLICE_X91Y106_C_CY, CLBLM_L_X60Y106_SLICE_X91Y106_B_CY, CLBLM_L_X60Y106_SLICE_X91Y106_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_L_X60Y106_SLICE_X91Y106_D_XOR, CLBLM_L_X60Y106_SLICE_X91Y106_C_XOR, CLBLM_L_X60Y106_SLICE_X91Y106_B_XOR, CLBLM_L_X60Y106_SLICE_X91Y106_A_XOR}),
.S({CLBLM_L_X60Y106_SLICE_X91Y106_DO6, CLBLM_L_X60Y106_SLICE_X91Y106_CO6, CLBLM_L_X60Y106_SLICE_X91Y106_BO6, CLBLM_L_X60Y106_SLICE_X91Y106_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X60Y106_SLICE_X91Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X60Y101_SLICE_X90Y101_AQ),
.O5(CLBLM_L_X60Y106_SLICE_X91Y106_DO5),
.O6(CLBLM_L_X60Y106_SLICE_X91Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X60Y106_SLICE_X91Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X62Y106_SLICE_X92Y106_CQ),
.O5(CLBLM_L_X60Y106_SLICE_X91Y106_CO5),
.O6(CLBLM_L_X60Y106_SLICE_X91Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X60Y106_SLICE_X91Y106_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X62Y106_SLICE_X92Y106_BQ),
.O5(CLBLM_L_X60Y106_SLICE_X91Y106_BO5),
.O6(CLBLM_L_X60Y106_SLICE_X91Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X60Y106_SLICE_X91Y106_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X62Y104_SLICE_X92Y104_BQ),
.O5(CLBLM_L_X60Y106_SLICE_X91Y106_AO5),
.O6(CLBLM_L_X60Y106_SLICE_X91Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y107_SLICE_X90Y107_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y100_SLICE_X90Y100_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X60Y107_SLICE_X90Y107_AO5),
.Q(CLBLM_L_X60Y107_SLICE_X90Y107_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X60Y107_SLICE_X90Y107_CARRY4 (
.CI(CLBLM_L_X60Y106_SLICE_X90Y106_COUT),
.CO({CLBLM_L_X60Y107_SLICE_X90Y107_D_CY, CLBLM_L_X60Y107_SLICE_X90Y107_C_CY, CLBLM_L_X60Y107_SLICE_X90Y107_B_CY, CLBLM_L_X60Y107_SLICE_X90Y107_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_L_X60Y107_SLICE_X90Y107_D_XOR, CLBLM_L_X60Y107_SLICE_X90Y107_C_XOR, CLBLM_L_X60Y107_SLICE_X90Y107_B_XOR, CLBLM_L_X60Y107_SLICE_X90Y107_A_XOR}),
.S({CLBLM_L_X60Y107_SLICE_X90Y107_DO6, CLBLM_L_X60Y107_SLICE_X90Y107_CO6, CLBLM_L_X60Y107_SLICE_X90Y107_BO6, CLBLM_L_X60Y107_SLICE_X90Y107_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X60Y107_SLICE_X90Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X60Y109_SLICE_X91Y109_BQ),
.O5(CLBLM_L_X60Y107_SLICE_X90Y107_DO5),
.O6(CLBLM_L_X60Y107_SLICE_X90Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X60Y107_SLICE_X90Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X62Y107_SLICE_X92Y107_AQ),
.O5(CLBLM_L_X60Y107_SLICE_X90Y107_CO5),
.O6(CLBLM_L_X60Y107_SLICE_X90Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X60Y107_SLICE_X90Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X60Y109_SLICE_X91Y109_AQ),
.O5(CLBLM_L_X60Y107_SLICE_X90Y107_BO5),
.O6(CLBLM_L_X60Y107_SLICE_X90Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ff00ff00)
  ) CLBLM_L_X60Y107_SLICE_X90Y107_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X60Y101_SLICE_X90Y101_AQ),
.I3(CLBLM_L_X62Y107_SLICE_X92Y107_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y107_SLICE_X90Y107_AO5),
.O6(CLBLM_L_X60Y107_SLICE_X90Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y107_SLICE_X91Y107_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y100_SLICE_X90Y100_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X60Y107_SLICE_X91Y107_AO5),
.Q(CLBLM_L_X60Y107_SLICE_X91Y107_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X60Y107_SLICE_X91Y107_CARRY4 (
.CI(CLBLM_L_X60Y106_SLICE_X91Y106_COUT),
.CO({CLBLM_L_X60Y107_SLICE_X91Y107_D_CY, CLBLM_L_X60Y107_SLICE_X91Y107_C_CY, CLBLM_L_X60Y107_SLICE_X91Y107_B_CY, CLBLM_L_X60Y107_SLICE_X91Y107_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_L_X60Y107_SLICE_X91Y107_D_XOR, CLBLM_L_X60Y107_SLICE_X91Y107_C_XOR, CLBLM_L_X60Y107_SLICE_X91Y107_B_XOR, CLBLM_L_X60Y107_SLICE_X91Y107_A_XOR}),
.S({CLBLM_L_X60Y107_SLICE_X91Y107_DO6, CLBLM_L_X60Y107_SLICE_X91Y107_CO6, CLBLM_L_X60Y107_SLICE_X91Y107_BO6, CLBLM_L_X60Y107_SLICE_X91Y107_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y107_SLICE_X91Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y107_SLICE_X91Y107_DO5),
.O6(CLBLM_L_X60Y107_SLICE_X91Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X60Y107_SLICE_X91Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X60Y109_SLICE_X91Y109_BQ),
.O5(CLBLM_L_X60Y107_SLICE_X91Y107_CO5),
.O6(CLBLM_L_X60Y107_SLICE_X91Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X60Y107_SLICE_X91Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X62Y107_SLICE_X92Y107_AQ),
.O5(CLBLM_L_X60Y107_SLICE_X91Y107_BO5),
.O6(CLBLM_L_X60Y107_SLICE_X91Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000cccccccc)
  ) CLBLM_L_X60Y107_SLICE_X91Y107_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X62Y107_SLICE_X92Y107_BO6),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X60Y109_SLICE_X91Y109_AQ),
.I5(1'b1),
.O5(CLBLM_L_X60Y107_SLICE_X91Y107_AO5),
.O6(CLBLM_L_X60Y107_SLICE_X91Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y108_SLICE_X90Y108_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y102_SLICE_X92Y102_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X60Y108_SLICE_X90Y108_BO5),
.Q(CLBLM_L_X60Y108_SLICE_X90Y108_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X60Y108_SLICE_X90Y108_CARRY4 (
.CI(1'b0),
.CO({CLBLM_L_X60Y108_SLICE_X90Y108_D_CY, CLBLM_L_X60Y108_SLICE_X90Y108_C_CY, CLBLM_L_X60Y108_SLICE_X90Y108_B_CY, CLBLM_L_X60Y108_SLICE_X90Y108_A_CY}),
.CYINIT(CLBLM_L_X60Y100_SLICE_X90Y100_AQ),
.DI({1'b0, 1'b0, 1'b0, CLBLM_L_X60Y108_SLICE_X90Y108_AO5}),
.O({CLBLM_L_X60Y108_SLICE_X90Y108_D_XOR, CLBLM_L_X60Y108_SLICE_X90Y108_C_XOR, CLBLM_L_X60Y108_SLICE_X90Y108_B_XOR, CLBLM_L_X60Y108_SLICE_X90Y108_A_XOR}),
.S({CLBLM_L_X60Y108_SLICE_X90Y108_DO6, CLBLM_L_X60Y108_SLICE_X90Y108_CO6, CLBLM_L_X60Y108_SLICE_X90Y108_BO6, CLBLM_L_X60Y108_SLICE_X90Y108_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X60Y108_SLICE_X90Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X60Y104_SLICE_X90Y104_AQ),
.O5(CLBLM_L_X60Y108_SLICE_X90Y108_DO5),
.O6(CLBLM_L_X60Y108_SLICE_X90Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X60Y108_SLICE_X90Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X59Y104_SLICE_X89Y104_CQ),
.O5(CLBLM_L_X60Y108_SLICE_X90Y108_CO5),
.O6(CLBLM_L_X60Y108_SLICE_X90Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccff00ff00)
  ) CLBLM_L_X60Y108_SLICE_X90Y108_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X59Y105_SLICE_X89Y105_CQ),
.I2(1'b1),
.I3(CLBLM_L_X62Y108_SLICE_X92Y108_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y108_SLICE_X90Y108_BO5),
.O6(CLBLM_L_X60Y108_SLICE_X90Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000000000)
  ) CLBLM_L_X60Y108_SLICE_X90Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X59Y106_SLICE_X89Y106_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y108_SLICE_X90Y108_AO5),
.O6(CLBLM_L_X60Y108_SLICE_X90Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y108_SLICE_X91Y108_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y100_SLICE_X90Y100_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X60Y108_SLICE_X91Y108_AO6),
.Q(CLBLM_L_X60Y108_SLICE_X91Y108_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd5dad0df858a808)
  ) CLBLM_L_X60Y108_SLICE_X91Y108_DLUT (
.I0(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I1(CLBLL_R_X57Y106_SLICE_X86Y106_D_XOR),
.I2(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I3(CLBLL_R_X57Y103_SLICE_X87Y103_AQ),
.I4(CLBLL_R_X57Y110_SLICE_X87Y110_A_XOR),
.I5(CLBLM_R_X59Y107_SLICE_X89Y107_BQ),
.O5(CLBLM_L_X60Y108_SLICE_X91Y108_DO5),
.O6(CLBLM_L_X60Y108_SLICE_X91Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffef0f2ff0e00020)
  ) CLBLM_L_X60Y108_SLICE_X91Y108_CLUT (
.I0(CLBLM_L_X60Y105_SLICE_X91Y105_D_XOR),
.I1(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I2(CLBLM_R_X59Y103_SLICE_X89Y103_CQ),
.I3(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I4(CLBLM_L_X60Y102_SLICE_X90Y102_BQ),
.I5(CLBLM_R_X59Y106_SLICE_X89Y106_AO5),
.O5(CLBLM_L_X60Y108_SLICE_X91Y108_CO5),
.O6(CLBLM_L_X60Y108_SLICE_X91Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50fa50eeee4444)
  ) CLBLM_L_X60Y108_SLICE_X91Y108_BLUT (
.I0(CLBLM_L_X62Y106_SLICE_X92Y106_AO5),
.I1(CLBLL_R_X57Y108_SLICE_X87Y108_CO6),
.I2(CLBLL_R_X57Y105_SLICE_X86Y105_AQ),
.I3(CLBLM_R_X59Y108_SLICE_X88Y108_C_XOR),
.I4(CLBLM_L_X60Y108_SLICE_X90Y108_B_XOR),
.I5(CLBLM_R_X59Y106_SLICE_X89Y106_AO6),
.O5(CLBLM_L_X60Y108_SLICE_X91Y108_BO5),
.O6(CLBLM_L_X60Y108_SLICE_X91Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0bb88f0f0ff00)
  ) CLBLM_L_X60Y108_SLICE_X91Y108_ALUT (
.I0(CLBLL_R_X57Y106_SLICE_X87Y106_D_XOR),
.I1(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I2(CLBLM_L_X62Y97_SLICE_X92Y97_AO6),
.I3(CLBLL_R_X57Y107_SLICE_X86Y107_D_XOR),
.I4(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I5(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.O5(CLBLM_L_X60Y108_SLICE_X91Y108_AO5),
.O6(CLBLM_L_X60Y108_SLICE_X91Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X60Y109_SLICE_X90Y109_CARRY4 (
.CI(CLBLM_L_X60Y108_SLICE_X90Y108_COUT),
.CO({CLBLM_L_X60Y109_SLICE_X90Y109_D_CY, CLBLM_L_X60Y109_SLICE_X90Y109_C_CY, CLBLM_L_X60Y109_SLICE_X90Y109_B_CY, CLBLM_L_X60Y109_SLICE_X90Y109_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_L_X60Y109_SLICE_X90Y109_D_XOR, CLBLM_L_X60Y109_SLICE_X90Y109_C_XOR, CLBLM_L_X60Y109_SLICE_X90Y109_B_XOR, CLBLM_L_X60Y109_SLICE_X90Y109_A_XOR}),
.S({CLBLM_L_X60Y109_SLICE_X90Y109_DO6, CLBLM_L_X60Y109_SLICE_X90Y109_CO6, CLBLM_L_X60Y109_SLICE_X90Y109_BO6, CLBLM_L_X60Y109_SLICE_X90Y109_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X60Y109_SLICE_X90Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X59Y111_SLICE_X89Y111_CQ),
.O5(CLBLM_L_X60Y109_SLICE_X90Y109_DO5),
.O6(CLBLM_L_X60Y109_SLICE_X90Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X60Y109_SLICE_X90Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X59Y106_SLICE_X89Y106_BQ),
.O5(CLBLM_L_X60Y109_SLICE_X90Y109_CO5),
.O6(CLBLM_L_X60Y109_SLICE_X90Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X60Y109_SLICE_X90Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X59Y112_SLICE_X89Y112_BQ),
.O5(CLBLM_L_X60Y109_SLICE_X90Y109_BO5),
.O6(CLBLM_L_X60Y109_SLICE_X90Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X60Y109_SLICE_X90Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X59Y112_SLICE_X89Y112_AQ),
.O5(CLBLM_L_X60Y109_SLICE_X90Y109_AO5),
.O6(CLBLM_L_X60Y109_SLICE_X90Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y109_SLICE_X91Y109_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y102_SLICE_X92Y102_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X60Y109_SLICE_X91Y109_AO6),
.Q(CLBLM_L_X60Y109_SLICE_X91Y109_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X60Y109_SLICE_X91Y109_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y102_SLICE_X92Y102_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X60Y109_SLICE_X91Y109_BO6),
.Q(CLBLM_L_X60Y109_SLICE_X91Y109_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaff005500ff00)
  ) CLBLM_L_X60Y109_SLICE_X91Y109_DLUT (
.I0(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X59Y110_SLICE_X89Y110_AQ),
.I4(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I5(CLBLM_L_X60Y107_SLICE_X90Y107_D_XOR),
.O5(CLBLM_L_X60Y109_SLICE_X91Y109_DO5),
.O6(CLBLM_L_X60Y109_SLICE_X91Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000e4ffe400)
  ) CLBLM_L_X60Y109_SLICE_X91Y109_CLUT (
.I0(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I1(CLBLM_L_X60Y107_SLICE_X91Y107_C_XOR),
.I2(CLBLM_L_X60Y109_SLICE_X91Y109_BQ),
.I3(CLBLM_R_X59Y103_SLICE_X89Y103_CQ),
.I4(CLBLM_L_X60Y109_SLICE_X91Y109_DO6),
.I5(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.O5(CLBLM_L_X60Y109_SLICE_X91Y109_CO5),
.O6(CLBLM_L_X60Y109_SLICE_X91Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88d8d8d8d8d8d8)
  ) CLBLM_L_X60Y109_SLICE_X91Y109_BLUT (
.I0(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I1(CLBLM_L_X62Y100_SLICE_X93Y100_BO6),
.I2(CLBLM_L_X60Y107_SLICE_X91Y107_C_XOR),
.I3(CLBLM_L_X60Y104_SLICE_X91Y104_C_XOR),
.I4(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I5(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.O5(CLBLM_L_X60Y109_SLICE_X91Y109_BO5),
.O6(CLBLM_L_X60Y109_SLICE_X91Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafacacaca0acacac)
  ) CLBLM_L_X60Y109_SLICE_X91Y109_ALUT (
.I0(CLBLM_L_X62Y97_SLICE_X92Y97_BO6),
.I1(CLBLM_L_X60Y107_SLICE_X91Y107_A_XOR),
.I2(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I3(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I4(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I5(CLBLM_L_X60Y104_SLICE_X91Y104_A_XOR),
.O5(CLBLM_L_X60Y109_SLICE_X91Y109_AO5),
.O6(CLBLM_L_X60Y109_SLICE_X91Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X60Y110_SLICE_X90Y110_CARRY4 (
.CI(CLBLM_L_X60Y109_SLICE_X90Y109_COUT),
.CO({CLBLM_L_X60Y110_SLICE_X90Y110_D_CY, CLBLM_L_X60Y110_SLICE_X90Y110_C_CY, CLBLM_L_X60Y110_SLICE_X90Y110_B_CY, CLBLM_L_X60Y110_SLICE_X90Y110_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_L_X60Y110_SLICE_X90Y110_D_XOR, CLBLM_L_X60Y110_SLICE_X90Y110_C_XOR, CLBLM_L_X60Y110_SLICE_X90Y110_B_XOR, CLBLM_L_X60Y110_SLICE_X90Y110_A_XOR}),
.S({CLBLM_L_X60Y110_SLICE_X90Y110_DO6, CLBLM_L_X60Y110_SLICE_X90Y110_CO6, CLBLM_L_X60Y110_SLICE_X90Y110_BO6, CLBLM_L_X60Y110_SLICE_X90Y110_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y110_SLICE_X90Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y110_SLICE_X90Y110_DO5),
.O6(CLBLM_L_X60Y110_SLICE_X90Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X60Y110_SLICE_X90Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X59Y110_SLICE_X89Y110_AQ),
.O5(CLBLM_L_X60Y110_SLICE_X90Y110_CO5),
.O6(CLBLM_L_X60Y110_SLICE_X90Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X60Y110_SLICE_X90Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X59Y111_SLICE_X89Y111_BQ),
.O5(CLBLM_L_X60Y110_SLICE_X90Y110_BO5),
.O6(CLBLM_L_X60Y110_SLICE_X90Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X60Y110_SLICE_X90Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X59Y111_SLICE_X89Y111_AQ),
.O5(CLBLM_L_X60Y110_SLICE_X90Y110_AO5),
.O6(CLBLM_L_X60Y110_SLICE_X90Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X60Y110_SLICE_X91Y110_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_R_X59Y99_SLICE_X89Y99_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X60Y110_SLICE_X91Y110_AO6),
.Q(CLBLM_L_X60Y110_SLICE_X91Y110_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbf80bf80bf80bf80)
  ) CLBLM_L_X60Y110_SLICE_X91Y110_DLUT (
.I0(CLBLM_L_X60Y106_SLICE_X90Y106_C_XOR),
.I1(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I2(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I3(CLBLM_R_X59Y112_SLICE_X89Y112_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y110_SLICE_X91Y110_DO5),
.O6(CLBLM_L_X60Y110_SLICE_X91Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbffbbff88008800)
  ) CLBLM_L_X60Y110_SLICE_X91Y110_CLUT (
.I0(CLBLM_L_X60Y107_SLICE_X90Y107_C_XOR),
.I1(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I2(1'b1),
.I3(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I4(1'b1),
.I5(CLBLM_R_X59Y111_SLICE_X89Y111_BQ),
.O5(CLBLM_L_X60Y110_SLICE_X91Y110_CO5),
.O6(CLBLM_L_X60Y110_SLICE_X91Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfecef2c23e0e3202)
  ) CLBLM_L_X60Y110_SLICE_X91Y110_BLUT (
.I0(CLBLM_L_X60Y108_SLICE_X91Y108_DO6),
.I1(CLBLM_R_X59Y106_SLICE_X89Y106_AO6),
.I2(CLBLM_L_X62Y106_SLICE_X92Y106_AO5),
.I3(CLBLM_L_X60Y108_SLICE_X90Y108_D_XOR),
.I4(CLBLL_R_X57Y103_SLICE_X87Y103_AQ),
.I5(CLBLM_R_X59Y109_SLICE_X88Y109_A_XOR),
.O5(CLBLM_L_X60Y110_SLICE_X91Y110_BO5),
.O6(CLBLM_L_X60Y110_SLICE_X91Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddd8ddd88d888d88)
  ) CLBLM_L_X60Y110_SLICE_X91Y110_ALUT (
.I0(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I1(CLBLM_R_X49Y104_SLICE_X75Y104_DQ),
.I2(CLBLM_R_X59Y103_SLICE_X89Y103_DQ),
.I3(CLBLM_L_X60Y110_SLICE_X91Y110_BO6),
.I4(1'b1),
.I5(CLBLM_L_X60Y108_SLICE_X91Y108_CO6),
.O5(CLBLM_L_X60Y110_SLICE_X91Y110_AO5),
.O6(CLBLM_L_X60Y110_SLICE_X91Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X60Y111_SLICE_X90Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_R_X59Y99_SLICE_X89Y99_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X60Y111_SLICE_X90Y111_AO6),
.Q(CLBLM_L_X60Y111_SLICE_X90Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5fff5ffa000a000)
  ) CLBLM_L_X60Y111_SLICE_X90Y111_DLUT (
.I0(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I1(1'b1),
.I2(CLBLM_L_X60Y107_SLICE_X90Y107_B_XOR),
.I3(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I4(1'b1),
.I5(CLBLM_R_X59Y111_SLICE_X89Y111_AQ),
.O5(CLBLM_L_X60Y111_SLICE_X90Y111_DO5),
.O6(CLBLM_L_X60Y111_SLICE_X90Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff37cc04fb33c800)
  ) CLBLM_L_X60Y111_SLICE_X90Y111_CLUT (
.I0(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I1(CLBLM_R_X59Y103_SLICE_X89Y103_CQ),
.I2(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I3(CLBLM_L_X60Y109_SLICE_X91Y109_AQ),
.I4(CLBLM_L_X60Y111_SLICE_X90Y111_DO6),
.I5(CLBLM_L_X60Y107_SLICE_X91Y107_A_XOR),
.O5(CLBLM_L_X60Y111_SLICE_X90Y111_CO5),
.O6(CLBLM_L_X60Y111_SLICE_X90Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffd8aad855d800d8)
  ) CLBLM_L_X60Y111_SLICE_X90Y111_BLUT (
.I0(CLBLM_L_X62Y106_SLICE_X92Y106_AO5),
.I1(CLBLM_L_X60Y109_SLICE_X90Y109_D_XOR),
.I2(CLBLM_R_X59Y111_SLICE_X88Y111_BO6),
.I3(CLBLM_R_X59Y106_SLICE_X89Y106_AO6),
.I4(CLBLM_L_X60Y108_SLICE_X91Y108_AQ),
.I5(CLBLM_R_X59Y110_SLICE_X88Y110_A_XOR),
.O5(CLBLM_L_X60Y111_SLICE_X90Y111_BO5),
.O6(CLBLM_L_X60Y111_SLICE_X90Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe0efe0ef202f202)
  ) CLBLM_L_X60Y111_SLICE_X90Y111_ALUT (
.I0(CLBLM_R_X59Y111_SLICE_X88Y111_CO6),
.I1(CLBLM_R_X59Y103_SLICE_X89Y103_DQ),
.I2(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I3(CLBLM_R_X49Y107_SLICE_X75Y107_DQ),
.I4(1'b1),
.I5(CLBLM_L_X60Y111_SLICE_X90Y111_CO6),
.O5(CLBLM_L_X60Y111_SLICE_X90Y111_AO5),
.O6(CLBLM_L_X60Y111_SLICE_X90Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X60Y111_SLICE_X91Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_R_X59Y99_SLICE_X89Y99_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X60Y111_SLICE_X91Y111_AO6),
.Q(CLBLM_L_X60Y111_SLICE_X91Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X60Y111_SLICE_X91Y111_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_R_X59Y99_SLICE_X89Y99_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X60Y111_SLICE_X91Y111_BO6),
.Q(CLBLM_L_X60Y111_SLICE_X91Y111_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaaaaaaaaaaaa)
  ) CLBLM_L_X60Y111_SLICE_X91Y111_DLUT (
.I0(CLBLM_R_X59Y111_SLICE_X89Y111_CQ),
.I1(CLBLM_L_X60Y107_SLICE_X90Y107_A_XOR),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I5(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.O5(CLBLM_L_X60Y111_SLICE_X91Y111_DO5),
.O6(CLBLM_L_X60Y111_SLICE_X91Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a0f5dda088)
  ) CLBLM_L_X60Y111_SLICE_X91Y111_CLUT (
.I0(CLBLM_R_X59Y103_SLICE_X89Y103_CQ),
.I1(CLBLM_L_X60Y106_SLICE_X91Y106_D_XOR),
.I2(CLBLM_L_X60Y101_SLICE_X90Y101_AQ),
.I3(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I4(CLBLM_L_X60Y111_SLICE_X91Y111_DO6),
.I5(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.O5(CLBLM_L_X60Y111_SLICE_X91Y111_CO5),
.O6(CLBLM_L_X60Y111_SLICE_X91Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaffccaaaa00cc)
  ) CLBLM_L_X60Y111_SLICE_X91Y111_BLUT (
.I0(CLBLM_R_X49Y108_SLICE_X75Y108_DQ),
.I1(CLBLM_L_X60Y111_SLICE_X90Y111_BO6),
.I2(1'b1),
.I3(CLBLM_R_X59Y103_SLICE_X89Y103_DQ),
.I4(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I5(CLBLM_L_X60Y111_SLICE_X91Y111_CO6),
.O5(CLBLM_L_X60Y111_SLICE_X91Y111_BO5),
.O6(CLBLM_L_X60Y111_SLICE_X91Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaaffaaccaa00)
  ) CLBLM_L_X60Y111_SLICE_X91Y111_ALUT (
.I0(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I1(CLBLM_L_X60Y109_SLICE_X91Y109_CO6),
.I2(1'b1),
.I3(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I4(CLBLM_R_X59Y103_SLICE_X89Y103_DQ),
.I5(CLBLM_R_X59Y111_SLICE_X89Y111_DO6),
.O5(CLBLM_L_X60Y111_SLICE_X91Y111_AO5),
.O6(CLBLM_L_X60Y111_SLICE_X91Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y112_SLICE_X90Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y112_SLICE_X90Y112_DO5),
.O6(CLBLM_L_X60Y112_SLICE_X90Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y112_SLICE_X90Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y112_SLICE_X90Y112_CO5),
.O6(CLBLM_L_X60Y112_SLICE_X90Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcfffcfcfffffdd)
  ) CLBLM_L_X60Y112_SLICE_X90Y112_BLUT (
.I0(CLBLM_R_X59Y99_SLICE_X89Y99_A5Q),
.I1(CLBLM_R_X59Y103_SLICE_X89Y103_DQ),
.I2(CLBLM_L_X60Y107_SLICE_X90Y107_AQ),
.I3(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I4(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I5(CLBLM_R_X59Y103_SLICE_X89Y103_CQ),
.O5(CLBLM_L_X60Y112_SLICE_X90Y112_BO5),
.O6(CLBLM_L_X60Y112_SLICE_X90Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff3fff3ff3ffff5)
  ) CLBLM_L_X60Y112_SLICE_X90Y112_ALUT (
.I0(CLBLM_R_X59Y99_SLICE_X89Y99_AQ),
.I1(CLBLM_R_X59Y108_SLICE_X88Y108_AQ),
.I2(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I3(CLBLM_R_X59Y103_SLICE_X89Y103_DQ),
.I4(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I5(CLBLM_R_X59Y103_SLICE_X89Y103_CQ),
.O5(CLBLM_L_X60Y112_SLICE_X90Y112_AO5),
.O6(CLBLM_L_X60Y112_SLICE_X90Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y112_SLICE_X91Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y112_SLICE_X91Y112_DO5),
.O6(CLBLM_L_X60Y112_SLICE_X91Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y112_SLICE_X91Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y112_SLICE_X91Y112_CO5),
.O6(CLBLM_L_X60Y112_SLICE_X91Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y112_SLICE_X91Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y112_SLICE_X91Y112_BO5),
.O6(CLBLM_L_X60Y112_SLICE_X91Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X60Y112_SLICE_X91Y112_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X60Y112_SLICE_X91Y112_AO5),
.O6(CLBLM_L_X60Y112_SLICE_X91Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y95_SLICE_X92Y95_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y98_SLICE_X93Y98_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y95_SLICE_X92Y95_AO5),
.Q(CLBLM_L_X62Y95_SLICE_X92Y95_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y95_SLICE_X92Y95_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y98_SLICE_X93Y98_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y95_SLICE_X92Y95_AO6),
.Q(CLBLM_L_X62Y95_SLICE_X92Y95_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y95_SLICE_X92Y95_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y95_SLICE_X92Y95_DO5),
.O6(CLBLM_L_X62Y95_SLICE_X92Y95_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y95_SLICE_X92Y95_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y95_SLICE_X92Y95_CO5),
.O6(CLBLM_L_X62Y95_SLICE_X92Y95_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff8000fffe0001)
  ) CLBLM_L_X62Y95_SLICE_X92Y95_BLUT (
.I0(CLBLM_L_X56Y98_SLICE_X85Y98_DQ),
.I1(CLBLM_L_X62Y98_SLICE_X92Y98_DQ),
.I2(CLBLM_L_X62Y95_SLICE_X92Y95_AQ),
.I3(CLBLM_L_X62Y98_SLICE_X92Y98_AQ),
.I4(CLBLM_L_X62Y95_SLICE_X92Y95_A5Q),
.I5(CLBLM_L_X62Y98_SLICE_X92Y98_CQ),
.O5(CLBLM_L_X62Y95_SLICE_X92Y95_BO5),
.O6(CLBLM_L_X62Y95_SLICE_X92Y95_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0f0faaaaff00)
  ) CLBLM_L_X62Y95_SLICE_X92Y95_ALUT (
.I0(CLBLM_L_X50Y106_SLICE_X76Y106_AQ),
.I1(CLBLM_L_X50Y104_SLICE_X76Y104_AQ),
.I2(CLBLM_L_X62Y95_SLICE_X92Y95_AQ),
.I3(CLBLM_L_X62Y95_SLICE_X92Y95_BO6),
.I4(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I5(1'b1),
.O5(CLBLM_L_X62Y95_SLICE_X92Y95_AO5),
.O6(CLBLM_L_X62Y95_SLICE_X92Y95_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y95_SLICE_X93Y95_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_AQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y95_SLICE_X93Y95_DO5),
.Q(CLBLM_L_X62Y95_SLICE_X93Y95_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y95_SLICE_X93Y95_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_AQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y95_SLICE_X93Y95_BO5),
.Q(CLBLM_L_X62Y95_SLICE_X93Y95_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y95_SLICE_X93Y95_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_AQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y95_SLICE_X93Y95_AO5),
.Q(CLBLM_L_X62Y95_SLICE_X93Y95_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y95_SLICE_X93Y95_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_AQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y95_SLICE_X93Y95_CO5),
.Q(CLBLM_L_X62Y95_SLICE_X93Y95_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y95_SLICE_X93Y95_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_AQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y95_SLICE_X93Y95_DO6),
.Q(CLBLM_L_X62Y95_SLICE_X93Y95_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555566666666)
  ) CLBLM_L_X62Y95_SLICE_X93Y95_DLUT (
.I0(CLBLM_L_X62Y95_SLICE_X92Y95_AQ),
.I1(CLBLM_L_X62Y98_SLICE_X92Y98_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y95_SLICE_X93Y95_DO5),
.O6(CLBLM_L_X62Y95_SLICE_X93Y95_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000016ccccccc)
  ) CLBLM_L_X62Y95_SLICE_X93Y95_CLUT (
.I0(CLBLM_L_X62Y95_SLICE_X92Y95_AQ),
.I1(CLBLM_L_X62Y95_SLICE_X92Y95_A5Q),
.I2(CLBLM_L_X62Y98_SLICE_X92Y98_AQ),
.I3(CLBLM_L_X62Y98_SLICE_X92Y98_CQ),
.I4(CLBLM_L_X62Y98_SLICE_X92Y98_DQ),
.I5(1'b1),
.O5(CLBLM_L_X62Y95_SLICE_X93Y95_CO5),
.O6(CLBLM_L_X62Y95_SLICE_X93Y95_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000055aaaaaa)
  ) CLBLM_L_X62Y95_SLICE_X93Y95_BLUT (
.I0(CLBLM_L_X62Y98_SLICE_X92Y98_DQ),
.I1(CLBLM_L_X62Y98_SLICE_X92Y98_AQ),
.I2(CLBLM_L_X62Y95_SLICE_X92Y95_A5Q),
.I3(CLBLM_L_X62Y98_SLICE_X92Y98_CQ),
.I4(CLBLM_L_X62Y95_SLICE_X92Y95_AQ),
.I5(1'b1),
.O5(CLBLM_L_X62Y95_SLICE_X93Y95_BO5),
.O6(CLBLM_L_X62Y95_SLICE_X93Y95_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6cccccc96c6ccccc)
  ) CLBLM_L_X62Y95_SLICE_X93Y95_ALUT (
.I0(CLBLM_L_X62Y98_SLICE_X92Y98_CQ),
.I1(CLBLM_L_X62Y98_SLICE_X92Y98_AQ),
.I2(CLBLM_L_X62Y98_SLICE_X92Y98_DQ),
.I3(CLBLM_L_X56Y98_SLICE_X85Y98_DQ),
.I4(CLBLM_L_X62Y95_SLICE_X92Y95_AQ),
.I5(1'b1),
.O5(CLBLM_L_X62Y95_SLICE_X93Y95_AO5),
.O6(CLBLM_L_X62Y95_SLICE_X93Y95_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y96_SLICE_X92Y96_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y99_SLICE_X93Y99_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y96_SLICE_X92Y96_CO6),
.Q(CLBLM_L_X62Y96_SLICE_X92Y96_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y96_SLICE_X92Y96_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y96_SLICE_X92Y96_DO5),
.O6(CLBLM_L_X62Y96_SLICE_X92Y96_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0acacafa0acac)
  ) CLBLM_L_X62Y96_SLICE_X92Y96_CLUT (
.I0(CLBLM_L_X50Y106_SLICE_X76Y106_CQ),
.I1(CLBLM_R_X63Y96_SLICE_X94Y96_AO6),
.I2(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I3(CLBLM_R_X63Y98_SLICE_X95Y98_B5Q),
.I4(CLBLM_L_X56Y98_SLICE_X85Y98_DQ),
.I5(1'b1),
.O5(CLBLM_L_X62Y96_SLICE_X92Y96_CO5),
.O6(CLBLM_L_X62Y96_SLICE_X92Y96_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff0000aaf0aaf0)
  ) CLBLM_L_X62Y96_SLICE_X92Y96_BLUT (
.I0(CLBLM_L_X62Y96_SLICE_X92Y96_CQ),
.I1(1'b1),
.I2(CLBLM_R_X63Y95_SLICE_X95Y95_B5Q),
.I3(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I4(CLBLM_R_X63Y96_SLICE_X95Y96_AQ),
.I5(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.O5(CLBLM_L_X62Y96_SLICE_X92Y96_BO5),
.O6(CLBLM_L_X62Y96_SLICE_X92Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55aa00d8d8d8d8)
  ) CLBLM_L_X62Y96_SLICE_X92Y96_ALUT (
.I0(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I1(CLBLM_R_X63Y98_SLICE_X94Y98_C5Q),
.I2(CLBLM_L_X62Y97_SLICE_X92Y97_C5Q),
.I3(CLBLM_L_X62Y99_SLICE_X93Y99_AQ),
.I4(CLBLM_R_X63Y98_SLICE_X95Y98_C5Q),
.I5(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.O5(CLBLM_L_X62Y96_SLICE_X92Y96_AO5),
.O6(CLBLM_L_X62Y96_SLICE_X92Y96_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X62Y96_SLICE_X92Y96_MUXF7A (
.I0(CLBLM_L_X62Y96_SLICE_X92Y96_BO6),
.I1(CLBLM_L_X62Y96_SLICE_X92Y96_AO6),
.O(CLBLM_L_X62Y96_SLICE_X92Y96_F7AMUX_O),
.S(CLBLM_L_X62Y106_SLICE_X93Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y96_SLICE_X93Y96_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y99_SLICE_X93Y99_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y96_SLICE_X95Y96_AO6),
.Q(CLBLM_L_X62Y96_SLICE_X93Y96_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y96_SLICE_X93Y96_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y99_SLICE_X93Y99_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y96_SLICE_X93Y96_CO6),
.Q(CLBLM_L_X62Y96_SLICE_X93Y96_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y96_SLICE_X93Y96_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y99_SLICE_X93Y99_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y96_SLICE_X93Y96_DO6),
.Q(CLBLM_L_X62Y96_SLICE_X93Y96_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd8ddd8dd888d888)
  ) CLBLM_L_X62Y96_SLICE_X93Y96_DLUT (
.I0(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I1(CLBLM_L_X50Y104_SLICE_X76Y104_AQ),
.I2(CLBLM_L_X56Y98_SLICE_X85Y98_DQ),
.I3(CLBLM_L_X64Y97_SLICE_X96Y97_BQ),
.I4(1'b1),
.I5(CLBLM_R_X63Y96_SLICE_X94Y96_CO5),
.O5(CLBLM_L_X62Y96_SLICE_X93Y96_DO5),
.O6(CLBLM_L_X62Y96_SLICE_X93Y96_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55af05fa50aa00)
  ) CLBLM_L_X62Y96_SLICE_X93Y96_CLUT (
.I0(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I1(1'b1),
.I2(CLBLM_L_X56Y98_SLICE_X85Y98_DQ),
.I3(CLBLM_R_X49Y106_SLICE_X74Y106_AQ),
.I4(CLBLM_R_X63Y100_SLICE_X95Y100_A5Q),
.I5(CLBLM_R_X63Y95_SLICE_X94Y95_AO6),
.O5(CLBLM_L_X62Y96_SLICE_X93Y96_CO5),
.O6(CLBLM_L_X62Y96_SLICE_X93Y96_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaf0ccffcc00)
  ) CLBLM_L_X62Y96_SLICE_X93Y96_BLUT (
.I0(CLBLM_L_X62Y98_SLICE_X93Y98_AQ),
.I1(CLBLM_L_X62Y96_SLICE_X93Y96_BQ),
.I2(CLBLM_R_X63Y94_SLICE_X94Y94_AQ),
.I3(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I4(CLBLM_R_X63Y95_SLICE_X95Y95_D5Q),
.I5(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.O5(CLBLM_L_X62Y96_SLICE_X93Y96_BO5),
.O6(CLBLM_L_X62Y96_SLICE_X93Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbb8888f3c0f3c0)
  ) CLBLM_L_X62Y96_SLICE_X93Y96_ALUT (
.I0(CLBLM_L_X62Y97_SLICE_X93Y97_DQ),
.I1(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I2(CLBLM_R_X63Y98_SLICE_X95Y98_D5Q),
.I3(CLBLM_L_X62Y97_SLICE_X92Y97_D5Q),
.I4(CLBLM_R_X63Y99_SLICE_X94Y99_C5Q),
.I5(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.O5(CLBLM_L_X62Y96_SLICE_X93Y96_AO5),
.O6(CLBLM_L_X62Y96_SLICE_X93Y96_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X62Y96_SLICE_X93Y96_MUXF7A (
.I0(CLBLM_L_X62Y96_SLICE_X93Y96_BO6),
.I1(CLBLM_L_X62Y96_SLICE_X93Y96_AO6),
.O(CLBLM_L_X62Y96_SLICE_X93Y96_F7AMUX_O),
.S(CLBLM_L_X62Y106_SLICE_X93Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y97_SLICE_X92Y97_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y100_SLICE_X92Y100_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y97_SLICE_X92Y97_CO5),
.Q(CLBLM_L_X62Y97_SLICE_X92Y97_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y97_SLICE_X92Y97_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y100_SLICE_X92Y100_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X60Y97_SLICE_X91Y97_AO5),
.Q(CLBLM_L_X62Y97_SLICE_X92Y97_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y97_SLICE_X92Y97_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y100_SLICE_X92Y100_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y97_SLICE_X92Y97_AO5),
.Q(CLBLM_L_X62Y97_SLICE_X92Y97_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y97_SLICE_X92Y97_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y100_SLICE_X92Y100_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y97_SLICE_X92Y97_BO5),
.Q(CLBLM_L_X62Y97_SLICE_X92Y97_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y97_SLICE_X92Y97_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y100_SLICE_X92Y100_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y97_SLICE_X92Y97_CO6),
.Q(CLBLM_L_X62Y97_SLICE_X92Y97_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y97_SLICE_X92Y97_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y100_SLICE_X92Y100_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y97_SLICE_X92Y97_DO6),
.Q(CLBLM_L_X62Y97_SLICE_X92Y97_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0a0a0a0a0)
  ) CLBLM_L_X62Y97_SLICE_X92Y97_DLUT (
.I0(CLBLM_L_X62Y100_SLICE_X92Y100_AO6),
.I1(1'b1),
.I2(CLBLM_L_X50Y107_SLICE_X76Y107_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y97_SLICE_X92Y97_DO5),
.O6(CLBLM_L_X62Y97_SLICE_X92Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55aa0088888888)
  ) CLBLM_L_X62Y97_SLICE_X92Y97_CLUT (
.I0(CLBLM_L_X62Y100_SLICE_X92Y100_AO6),
.I1(CLBLM_L_X50Y106_SLICE_X76Y106_CQ),
.I2(1'b1),
.I3(CLBLM_L_X50Y106_SLICE_X76Y106_AQ),
.I4(CLBLM_L_X60Y97_SLICE_X91Y97_BQ),
.I5(1'b1),
.O5(CLBLM_L_X62Y97_SLICE_X92Y97_CO5),
.O6(CLBLM_L_X62Y97_SLICE_X92Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaf0aaaacccc)
  ) CLBLM_L_X62Y97_SLICE_X92Y97_BLUT (
.I0(CLBLM_L_X50Y105_SLICE_X77Y105_AQ),
.I1(CLBLM_L_X64Y97_SLICE_X96Y97_B5Q),
.I2(CLBLM_L_X62Y100_SLICE_X92Y100_BQ),
.I3(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I4(CLBLM_L_X62Y100_SLICE_X92Y100_AO6),
.I5(1'b1),
.O5(CLBLM_L_X62Y97_SLICE_X92Y97_BO5),
.O6(CLBLM_L_X62Y97_SLICE_X92Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacacacaaaaff00)
  ) CLBLM_L_X62Y97_SLICE_X92Y97_ALUT (
.I0(CLBLM_L_X50Y104_SLICE_X76Y104_AQ),
.I1(CLBLM_L_X62Y100_SLICE_X92Y100_AQ),
.I2(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I3(CLBLM_L_X64Y97_SLICE_X96Y97_BQ),
.I4(CLBLM_L_X62Y100_SLICE_X92Y100_AO6),
.I5(1'b1),
.O5(CLBLM_L_X62Y97_SLICE_X92Y97_AO5),
.O6(CLBLM_L_X62Y97_SLICE_X92Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y97_SLICE_X93Y97_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y100_SLICE_X92Y100_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y97_SLICE_X94Y97_CO6),
.Q(CLBLM_L_X62Y97_SLICE_X93Y97_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y97_SLICE_X93Y97_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y100_SLICE_X92Y100_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y97_SLICE_X93Y97_CO6),
.Q(CLBLM_L_X62Y97_SLICE_X93Y97_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y97_SLICE_X93Y97_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y100_SLICE_X92Y100_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y96_SLICE_X95Y96_AO6),
.Q(CLBLM_L_X62Y97_SLICE_X93Y97_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00dd00cc00000000)
  ) CLBLM_L_X62Y97_SLICE_X93Y97_DLUT (
.I0(CLBLM_L_X62Y96_SLICE_X92Y96_CQ),
.I1(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I2(1'b1),
.I3(CLBLM_L_X56Y97_SLICE_X85Y97_AQ),
.I4(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I5(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.O5(CLBLM_L_X62Y97_SLICE_X93Y97_DO5),
.O6(CLBLM_L_X62Y97_SLICE_X93Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00aafcaa0c)
  ) CLBLM_L_X62Y97_SLICE_X93Y97_CLUT (
.I0(CLBLM_L_X50Y107_SLICE_X76Y107_BQ),
.I1(CLBLM_L_X64Y96_SLICE_X96Y96_AO5),
.I2(CLBLM_L_X56Y98_SLICE_X85Y98_DQ),
.I3(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I4(CLBLM_R_X63Y98_SLICE_X95Y98_DQ),
.I5(1'b1),
.O5(CLBLM_L_X62Y97_SLICE_X93Y97_CO5),
.O6(CLBLM_L_X62Y97_SLICE_X93Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafafc0c0a0afc0c)
  ) CLBLM_L_X62Y97_SLICE_X93Y97_BLUT (
.I0(CLBLM_R_X63Y97_SLICE_X94Y97_CQ),
.I1(CLBLM_R_X63Y95_SLICE_X95Y95_C5Q),
.I2(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I3(CLBLM_L_X64Y97_SLICE_X97Y97_BQ),
.I4(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I5(CLBLM_L_X62Y98_SLICE_X93Y98_BQ),
.O5(CLBLM_L_X62Y97_SLICE_X93Y97_BO5),
.O6(CLBLM_L_X62Y97_SLICE_X93Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hacffacf0ac0fac00)
  ) CLBLM_L_X62Y97_SLICE_X93Y97_ALUT (
.I0(CLBLM_L_X62Y97_SLICE_X93Y97_CQ),
.I1(CLBLM_R_X63Y98_SLICE_X95Y98_DQ),
.I2(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I3(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I4(CLBLM_L_X62Y97_SLICE_X92Y97_DQ),
.I5(CLBLM_R_X63Y99_SLICE_X94Y99_CQ),
.O5(CLBLM_L_X62Y97_SLICE_X93Y97_AO5),
.O6(CLBLM_L_X62Y97_SLICE_X93Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X62Y97_SLICE_X93Y97_MUXF7A (
.I0(CLBLM_L_X62Y97_SLICE_X93Y97_BO6),
.I1(CLBLM_L_X62Y97_SLICE_X93Y97_AO6),
.O(CLBLM_L_X62Y97_SLICE_X93Y97_F7AMUX_O),
.S(CLBLM_L_X62Y106_SLICE_X93Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y98_SLICE_X92Y98_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y98_SLICE_X93Y98_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y98_SLICE_X92Y98_AO5),
.Q(CLBLM_L_X62Y98_SLICE_X92Y98_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y98_SLICE_X92Y98_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y98_SLICE_X93Y98_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y98_SLICE_X92Y98_BO6),
.Q(CLBLM_L_X62Y98_SLICE_X92Y98_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y98_SLICE_X92Y98_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y98_SLICE_X93Y98_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y98_SLICE_X92Y98_CO6),
.Q(CLBLM_L_X62Y98_SLICE_X92Y98_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y98_SLICE_X92Y98_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y98_SLICE_X93Y98_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y98_SLICE_X92Y98_DO6),
.Q(CLBLM_L_X62Y98_SLICE_X92Y98_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff006a6aa9a9)
  ) CLBLM_L_X62Y98_SLICE_X92Y98_DLUT (
.I0(CLBLM_L_X62Y98_SLICE_X92Y98_DQ),
.I1(CLBLM_L_X62Y98_SLICE_X92Y98_CQ),
.I2(CLBLM_L_X56Y98_SLICE_X85Y98_DQ),
.I3(CLBLM_R_X49Y105_SLICE_X75Y105_CQ),
.I4(CLBLM_L_X62Y95_SLICE_X92Y95_AQ),
.I5(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.O5(CLBLM_L_X62Y98_SLICE_X92Y98_DO5),
.O6(CLBLM_L_X62Y98_SLICE_X92Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff003c3cc3c3)
  ) CLBLM_L_X62Y98_SLICE_X92Y98_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X62Y98_SLICE_X92Y98_CQ),
.I2(CLBLM_L_X56Y98_SLICE_X85Y98_DQ),
.I3(CLBLM_L_X50Y105_SLICE_X77Y105_AQ),
.I4(CLBLM_L_X62Y95_SLICE_X92Y95_AQ),
.I5(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.O5(CLBLM_L_X62Y98_SLICE_X92Y98_CO5),
.O6(CLBLM_L_X62Y98_SLICE_X92Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff36ff9c0036009c)
  ) CLBLM_L_X62Y98_SLICE_X92Y98_BLUT (
.I0(CLBLM_L_X56Y98_SLICE_X85Y98_DQ),
.I1(CLBLM_L_X62Y98_SLICE_X92Y98_BQ),
.I2(CLBLM_L_X62Y95_SLICE_X93Y95_CO6),
.I3(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I4(CLBLM_L_X62Y95_SLICE_X93Y95_BO6),
.I5(CLBLM_L_X50Y106_SLICE_X76Y106_CQ),
.O5(CLBLM_L_X62Y98_SLICE_X92Y98_BO5),
.O6(CLBLM_L_X62Y98_SLICE_X92Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc808c808ff33cc00)
  ) CLBLM_L_X62Y98_SLICE_X92Y98_ALUT (
.I0(CLBLM_R_X49Y104_SLICE_X75Y104_CQ),
.I1(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I2(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I3(CLBLM_R_X49Y106_SLICE_X74Y106_AQ),
.I4(CLBLM_L_X62Y95_SLICE_X93Y95_AO6),
.I5(1'b1),
.O5(CLBLM_L_X62Y98_SLICE_X92Y98_AO5),
.O6(CLBLM_L_X62Y98_SLICE_X92Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y98_SLICE_X93Y98_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y98_SLICE_X93Y98_AO6),
.Q(CLBLM_L_X62Y98_SLICE_X93Y98_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y98_SLICE_X93Y98_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y98_SLICE_X93Y98_BO6),
.Q(CLBLM_L_X62Y98_SLICE_X93Y98_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffff7dfd7)
  ) CLBLM_L_X62Y98_SLICE_X93Y98_DLUT (
.I0(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I1(CLBLM_L_X56Y98_SLICE_X85Y98_A5Q),
.I2(CLBLM_L_X56Y98_SLICE_X85Y98_DQ),
.I3(CLBLM_L_X62Y98_SLICE_X93Y98_BQ),
.I4(CLBLM_L_X62Y98_SLICE_X93Y98_AQ),
.I5(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.O5(CLBLM_L_X62Y98_SLICE_X93Y98_DO5),
.O6(CLBLM_L_X62Y98_SLICE_X93Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0200aaaa0000aaaa)
  ) CLBLM_L_X62Y98_SLICE_X93Y98_CLUT (
.I0(CLBLM_L_X62Y99_SLICE_X92Y99_AO6),
.I1(CLBLM_L_X62Y100_SLICE_X93Y100_CO6),
.I2(CLBLM_R_X59Y102_SLICE_X88Y102_AQ),
.I3(CLBLL_R_X57Y101_SLICE_X86Y101_AO5),
.I4(CLBLM_L_X62Y98_SLICE_X93Y98_DO6),
.I5(CLBLM_L_X60Y98_SLICE_X90Y98_BQ),
.O5(CLBLM_L_X62Y98_SLICE_X93Y98_CO5),
.O6(CLBLM_L_X62Y98_SLICE_X93Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4fff4f4f00b00000)
  ) CLBLM_L_X62Y98_SLICE_X93Y98_BLUT (
.I0(CLBLM_R_X49Y119_SLICE_X74Y119_AQ),
.I1(CLBLM_R_X49Y119_SLICE_X74Y119_BQ),
.I2(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I3(CLBLM_L_X62Y98_SLICE_X92Y98_BQ),
.I4(CLBLM_L_X62Y95_SLICE_X93Y95_CO6),
.I5(CLBLM_L_X62Y98_SLICE_X93Y98_BQ),
.O5(CLBLM_L_X62Y98_SLICE_X93Y98_BO5),
.O6(CLBLM_L_X62Y98_SLICE_X93Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h44f4ffff00b00000)
  ) CLBLM_L_X62Y98_SLICE_X93Y98_ALUT (
.I0(CLBLM_R_X49Y119_SLICE_X74Y119_AQ),
.I1(CLBLM_R_X49Y119_SLICE_X74Y119_BQ),
.I2(CLBLM_L_X62Y95_SLICE_X93Y95_BO6),
.I3(CLBLM_L_X62Y98_SLICE_X92Y98_BQ),
.I4(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I5(CLBLM_L_X62Y98_SLICE_X93Y98_AQ),
.O5(CLBLM_L_X62Y98_SLICE_X93Y98_AO5),
.O6(CLBLM_L_X62Y98_SLICE_X93Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y99_SLICE_X92Y99_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y99_SLICE_X92Y99_BO6),
.Q(CLBLM_L_X62Y99_SLICE_X92Y99_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00a000a000a000a0)
  ) CLBLM_L_X62Y99_SLICE_X92Y99_DLUT (
.I0(CLBLL_R_X57Y99_SLICE_X87Y99_AQ),
.I1(1'b1),
.I2(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I3(CLBLM_L_X62Y99_SLICE_X92Y99_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y99_SLICE_X92Y99_DO5),
.O6(CLBLM_L_X62Y99_SLICE_X92Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3230363cfbf3fbbf)
  ) CLBLM_L_X62Y99_SLICE_X92Y99_CLUT (
.I0(CLBLM_L_X62Y104_SLICE_X93Y104_AQ),
.I1(CLBLM_L_X60Y110_SLICE_X91Y110_AQ),
.I2(CLBLM_L_X62Y103_SLICE_X92Y103_AQ),
.I3(CLBLM_R_X59Y102_SLICE_X88Y102_AQ),
.I4(CLBLM_R_X59Y102_SLICE_X89Y102_AQ),
.I5(CLBLM_L_X62Y106_SLICE_X93Y106_AQ),
.O5(CLBLM_L_X62Y99_SLICE_X92Y99_CO5),
.O6(CLBLM_L_X62Y99_SLICE_X92Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0ccccc5c5ccccc)
  ) CLBLM_L_X62Y99_SLICE_X92Y99_BLUT (
.I0(CLBLM_L_X62Y110_SLICE_X92Y110_DO6),
.I1(CLBLM_L_X62Y99_SLICE_X92Y99_BQ),
.I2(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I3(1'b1),
.I4(CLBLL_R_X57Y99_SLICE_X87Y99_AQ),
.I5(CLBLM_L_X62Y99_SLICE_X92Y99_CO6),
.O5(CLBLM_L_X62Y99_SLICE_X92Y99_BO5),
.O6(CLBLM_L_X62Y99_SLICE_X92Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa2222a0a02020)
  ) CLBLM_L_X62Y99_SLICE_X92Y99_ALUT (
.I0(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I1(CLBLM_R_X49Y119_SLICE_X74Y119_BQ),
.I2(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I3(1'b1),
.I4(CLBLM_R_X49Y119_SLICE_X74Y119_AQ),
.I5(1'b1),
.O5(CLBLM_L_X62Y99_SLICE_X92Y99_AO5),
.O6(CLBLM_L_X62Y99_SLICE_X92Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y99_SLICE_X93Y99_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y100_SLICE_X92Y100_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y95_SLICE_X95Y95_AO6),
.Q(CLBLM_L_X62Y99_SLICE_X93Y99_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000044440cc00cc0)
  ) CLBLM_L_X62Y99_SLICE_X93Y99_DLUT (
.I0(CLBLM_L_X60Y99_SLICE_X91Y99_AO6),
.I1(CLBLM_L_X62Y99_SLICE_X92Y99_AO5),
.I2(CLBLM_L_X56Y98_SLICE_X85Y98_DQ),
.I3(CLBLM_L_X56Y98_SLICE_X85Y98_A5Q),
.I4(CLBLM_L_X62Y99_SLICE_X93Y99_BO6),
.I5(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.O5(CLBLM_L_X62Y99_SLICE_X93Y99_DO5),
.O6(CLBLM_L_X62Y99_SLICE_X93Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0404040400cccc00)
  ) CLBLM_L_X62Y99_SLICE_X93Y99_CLUT (
.I0(CLBLM_L_X60Y99_SLICE_X91Y99_AO6),
.I1(CLBLM_L_X62Y99_SLICE_X92Y99_AO5),
.I2(CLBLM_L_X62Y100_SLICE_X93Y100_CO6),
.I3(CLBLM_L_X56Y98_SLICE_X85Y98_A5Q),
.I4(CLBLM_L_X56Y98_SLICE_X85Y98_DQ),
.I5(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.O5(CLBLM_L_X62Y99_SLICE_X93Y99_CO5),
.O6(CLBLM_L_X62Y99_SLICE_X93Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7ffffffffffffff)
  ) CLBLM_L_X62Y99_SLICE_X93Y99_BLUT (
.I0(CLBLM_L_X62Y103_SLICE_X92Y103_AQ),
.I1(CLBLM_L_X62Y106_SLICE_X93Y106_AQ),
.I2(CLBLM_L_X62Y110_SLICE_X92Y110_DO6),
.I3(CLBLM_L_X62Y104_SLICE_X93Y104_AQ),
.I4(CLBLM_R_X59Y102_SLICE_X89Y102_AQ),
.I5(CLBLM_L_X60Y110_SLICE_X91Y110_AQ),
.O5(CLBLM_L_X62Y99_SLICE_X93Y99_BO5),
.O6(CLBLM_L_X62Y99_SLICE_X93Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h10d0101020e02020)
  ) CLBLM_L_X62Y99_SLICE_X93Y99_ALUT (
.I0(CLBLM_L_X56Y98_SLICE_X85Y98_DQ),
.I1(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I2(CLBLM_L_X62Y99_SLICE_X92Y99_AO5),
.I3(CLBLM_L_X62Y99_SLICE_X93Y99_BO6),
.I4(CLBLM_L_X60Y99_SLICE_X90Y99_AO6),
.I5(CLBLM_L_X56Y98_SLICE_X85Y98_A5Q),
.O5(CLBLM_L_X62Y99_SLICE_X93Y99_AO5),
.O6(CLBLM_L_X62Y99_SLICE_X93Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X62Y100_SLICE_X92Y100_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y101_SLICE_X93Y101_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y104_SLICE_X74Y104_AQ),
.Q(CLBLM_L_X62Y100_SLICE_X92Y100_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X62Y100_SLICE_X92Y100_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y101_SLICE_X93Y101_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y104_SLICE_X75Y104_AQ),
.Q(CLBLM_L_X62Y100_SLICE_X92Y100_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X62Y100_SLICE_X92Y100_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y101_SLICE_X93Y101_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y104_SLICE_X75Y104_CQ),
.Q(CLBLM_L_X62Y100_SLICE_X92Y100_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00200000ffff0000)
  ) CLBLM_L_X62Y100_SLICE_X92Y100_DLUT (
.I0(CLBLM_L_X60Y99_SLICE_X90Y99_AO6),
.I1(CLBLM_L_X62Y104_SLICE_X93Y104_AQ),
.I2(CLBLM_R_X59Y102_SLICE_X89Y102_AQ),
.I3(CLBLM_L_X62Y102_SLICE_X93Y102_AO5),
.I4(CLBLM_L_X62Y99_SLICE_X92Y99_AO6),
.I5(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.O5(CLBLM_L_X62Y100_SLICE_X92Y100_DO5),
.O6(CLBLM_L_X62Y100_SLICE_X92Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h02000000ffff0000)
  ) CLBLM_L_X62Y100_SLICE_X92Y100_CLUT (
.I0(CLBLM_L_X60Y99_SLICE_X90Y99_AO6),
.I1(CLBLM_L_X60Y99_SLICE_X91Y99_BO6),
.I2(CLBLM_R_X59Y102_SLICE_X89Y102_AQ),
.I3(CLBLM_L_X62Y104_SLICE_X93Y104_AQ),
.I4(CLBLM_L_X62Y99_SLICE_X92Y99_AO6),
.I5(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.O5(CLBLM_L_X62Y100_SLICE_X92Y100_CO5),
.O6(CLBLM_L_X62Y100_SLICE_X92Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2000000000002000)
  ) CLBLM_L_X62Y100_SLICE_X92Y100_BLUT (
.I0(CLBLM_L_X56Y103_SLICE_X85Y103_CO6),
.I1(CLBLM_L_X62Y102_SLICE_X93Y102_AO5),
.I2(CLBLM_R_X59Y102_SLICE_X89Y102_AQ),
.I3(CLBLM_R_X59Y102_SLICE_X88Y102_AQ),
.I4(CLBLM_L_X60Y98_SLICE_X90Y98_BQ),
.I5(CLBLM_L_X62Y104_SLICE_X93Y104_AQ),
.O5(CLBLM_L_X62Y100_SLICE_X92Y100_BO5),
.O6(CLBLM_L_X62Y100_SLICE_X92Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2000000010000000)
  ) CLBLM_L_X62Y100_SLICE_X92Y100_ALUT (
.I0(CLBLM_R_X59Y102_SLICE_X89Y102_AQ),
.I1(CLBLM_L_X62Y102_SLICE_X93Y102_AO5),
.I2(CLBLM_L_X62Y104_SLICE_X93Y104_AQ),
.I3(CLBLM_R_X59Y102_SLICE_X88Y102_AQ),
.I4(CLBLM_L_X60Y98_SLICE_X90Y98_BQ),
.I5(1'b1),
.O5(CLBLM_L_X62Y100_SLICE_X92Y100_AO5),
.O6(CLBLM_L_X62Y100_SLICE_X92Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y100_SLICE_X93Y100_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y100_SLICE_X92Y100_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y100_SLICE_X93Y100_AO5),
.Q(CLBLM_L_X62Y100_SLICE_X93Y100_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y100_SLICE_X93Y100_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y100_SLICE_X92Y100_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y100_SLICE_X93Y100_BO5),
.Q(CLBLM_L_X62Y100_SLICE_X93Y100_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y100_SLICE_X93Y100_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y100_SLICE_X93Y100_DO5),
.O6(CLBLM_L_X62Y100_SLICE_X93Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffdfffffffffff)
  ) CLBLM_L_X62Y100_SLICE_X93Y100_CLUT (
.I0(CLBLM_L_X62Y103_SLICE_X92Y103_AQ),
.I1(CLBLM_L_X62Y104_SLICE_X93Y104_AQ),
.I2(CLBLM_R_X59Y102_SLICE_X89Y102_AQ),
.I3(CLBLM_L_X60Y110_SLICE_X91Y110_AQ),
.I4(CLBLM_L_X62Y110_SLICE_X92Y110_DO6),
.I5(CLBLM_L_X62Y106_SLICE_X93Y106_AQ),
.O5(CLBLM_L_X62Y100_SLICE_X93Y100_CO5),
.O6(CLBLM_L_X62Y100_SLICE_X93Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc00ccfafa0a0a)
  ) CLBLM_L_X62Y100_SLICE_X93Y100_BLUT (
.I0(CLBLM_R_X63Y100_SLICE_X95Y100_A5Q),
.I1(CLBLM_L_X62Y100_SLICE_X92Y100_CQ),
.I2(CLBLM_L_X62Y100_SLICE_X92Y100_AO6),
.I3(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I4(CLBLM_R_X49Y106_SLICE_X74Y106_AQ),
.I5(1'b1),
.O5(CLBLM_L_X62Y100_SLICE_X93Y100_BO5),
.O6(CLBLM_L_X62Y100_SLICE_X93Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00acacacac)
  ) CLBLM_L_X62Y100_SLICE_X93Y100_ALUT (
.I0(CLBLM_R_X49Y105_SLICE_X75Y105_CQ),
.I1(CLBLM_R_X63Y100_SLICE_X95Y100_AQ),
.I2(CLBLM_L_X62Y100_SLICE_X92Y100_AO6),
.I3(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I4(CLBLM_L_X62Y101_SLICE_X93Y101_AQ),
.I5(1'b1),
.O5(CLBLM_L_X62Y100_SLICE_X93Y100_AO5),
.O6(CLBLM_L_X62Y100_SLICE_X93Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y101_SLICE_X92Y101_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y99_SLICE_X92Y99_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y101_SLICE_X92Y101_AO6),
.Q(CLBLM_L_X62Y101_SLICE_X92Y101_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y101_SLICE_X92Y101_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y99_SLICE_X92Y99_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y101_SLICE_X92Y101_BO6),
.Q(CLBLM_L_X62Y101_SLICE_X92Y101_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y101_SLICE_X92Y101_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y99_SLICE_X92Y99_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y101_SLICE_X92Y101_CO6),
.Q(CLBLM_L_X62Y101_SLICE_X92Y101_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3c0c0bb88bb88)
  ) CLBLM_L_X62Y101_SLICE_X92Y101_DLUT (
.I0(CLBLM_L_X62Y101_SLICE_X92Y101_BQ),
.I1(CLBLM_L_X62Y99_SLICE_X92Y99_BQ),
.I2(CLBLM_L_X62Y101_SLICE_X92Y101_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(1'b1),
.O5(CLBLM_L_X62Y101_SLICE_X92Y101_DO5),
.O6(CLBLM_L_X62Y101_SLICE_X92Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cfc0cfcfc0c0)
  ) CLBLM_L_X62Y101_SLICE_X92Y101_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X62Y96_SLICE_X93Y96_F7AMUX_O),
.I2(CLBLM_L_X60Y99_SLICE_X90Y99_BO5),
.I3(CLBLM_R_X59Y104_SLICE_X89Y104_F7AMUX_O),
.I4(CLBLM_L_X62Y106_SLICE_X93Y106_DO6),
.I5(CLBLM_L_X62Y103_SLICE_X93Y103_BO6),
.O5(CLBLM_L_X62Y101_SLICE_X92Y101_CO5),
.O6(CLBLM_L_X62Y101_SLICE_X92Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0f5a0f5b1b1b1b1)
  ) CLBLM_L_X62Y101_SLICE_X92Y101_BLUT (
.I0(CLBLM_L_X60Y99_SLICE_X90Y99_BO5),
.I1(CLBLM_L_X62Y104_SLICE_X92Y104_DO6),
.I2(CLBLM_L_X62Y96_SLICE_X92Y96_F7AMUX_O),
.I3(CLBLM_R_X59Y105_SLICE_X88Y105_F7AMUX_O),
.I4(1'b1),
.I5(CLBLM_L_X62Y103_SLICE_X93Y103_BO6),
.O5(CLBLM_L_X62Y101_SLICE_X92Y101_BO5),
.O6(CLBLM_L_X62Y101_SLICE_X92Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcaaacaaaaaaaaaaa)
  ) CLBLM_L_X62Y101_SLICE_X92Y101_ALUT (
.I0(CLBLM_L_X60Y103_SLICE_X90Y103_F8MUX_O),
.I1(CLBLM_R_X63Y97_SLICE_X94Y97_F7AMUX_O),
.I2(CLBLM_R_X59Y102_SLICE_X89Y102_AQ),
.I3(CLBLM_L_X62Y106_SLICE_X93Y106_AQ),
.I4(1'b1),
.I5(CLBLM_L_X60Y110_SLICE_X91Y110_AQ),
.O5(CLBLM_L_X62Y101_SLICE_X92Y101_AO5),
.O6(CLBLM_L_X62Y101_SLICE_X92Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X62Y101_SLICE_X93Y101_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y101_SLICE_X93Y101_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y104_SLICE_X75Y104_BQ),
.Q(CLBLM_L_X62Y101_SLICE_X93Y101_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X62Y101_SLICE_X93Y101_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y101_SLICE_X93Y101_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y106_SLICE_X75Y106_DQ),
.Q(CLBLM_L_X62Y101_SLICE_X93Y101_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X62Y101_SLICE_X93Y101_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y101_SLICE_X93Y101_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y107_SLICE_X75Y107_CQ),
.Q(CLBLM_L_X62Y101_SLICE_X93Y101_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y101_SLICE_X93Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y101_SLICE_X93Y101_DO5),
.O6(CLBLM_L_X62Y101_SLICE_X93Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y101_SLICE_X93Y101_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y101_SLICE_X93Y101_CO5),
.O6(CLBLM_L_X62Y101_SLICE_X93Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y101_SLICE_X93Y101_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y101_SLICE_X93Y101_BO5),
.O6(CLBLM_L_X62Y101_SLICE_X93Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c000c0c0c000c0)
  ) CLBLM_L_X62Y101_SLICE_X93Y101_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I2(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I3(CLBLM_R_X49Y119_SLICE_X74Y119_BQ),
.I4(CLBLM_R_X49Y119_SLICE_X74Y119_AQ),
.I5(1'b1),
.O5(CLBLM_L_X62Y101_SLICE_X93Y101_AO5),
.O6(CLBLM_L_X62Y101_SLICE_X93Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y102_SLICE_X92Y102_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y102_SLICE_X92Y102_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y102_SLICE_X92Y102_BO6),
.Q(CLBLM_L_X62Y102_SLICE_X92Y102_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00440000ffff0000)
  ) CLBLM_L_X62Y102_SLICE_X92Y102_DLUT (
.I0(CLBLM_L_X60Y100_SLICE_X91Y100_AO6),
.I1(CLBLM_L_X62Y102_SLICE_X93Y102_AO6),
.I2(1'b1),
.I3(CLBLM_L_X62Y104_SLICE_X93Y104_AQ),
.I4(CLBLM_L_X62Y99_SLICE_X92Y99_AO6),
.I5(CLBLM_L_X60Y101_SLICE_X90Y101_BO6),
.O5(CLBLM_L_X62Y102_SLICE_X92Y102_DO5),
.O6(CLBLM_L_X62Y102_SLICE_X92Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000ffff0000)
  ) CLBLM_L_X62Y102_SLICE_X92Y102_CLUT (
.I0(CLBLM_L_X60Y99_SLICE_X90Y99_AO6),
.I1(CLBLM_L_X62Y102_SLICE_X93Y102_AO6),
.I2(CLBLM_L_X62Y104_SLICE_X93Y104_AQ),
.I3(CLBLL_R_X57Y101_SLICE_X86Y101_AO5),
.I4(CLBLM_L_X62Y99_SLICE_X92Y99_AO6),
.I5(CLBLM_L_X60Y101_SLICE_X90Y101_BO6),
.O5(CLBLM_L_X62Y102_SLICE_X92Y102_CO5),
.O6(CLBLM_L_X62Y102_SLICE_X92Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33f0330f330033)
  ) CLBLM_L_X62Y102_SLICE_X92Y102_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X62Y102_SLICE_X92Y102_BQ),
.I2(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I3(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I4(CLBLM_R_X49Y104_SLICE_X74Y104_AQ),
.I5(CLBLM_L_X50Y104_SLICE_X76Y104_AQ),
.O5(CLBLM_L_X62Y102_SLICE_X92Y102_BO5),
.O6(CLBLM_L_X62Y102_SLICE_X92Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa000000aa00f000)
  ) CLBLM_L_X62Y102_SLICE_X92Y102_ALUT (
.I0(CLBLM_L_X50Y106_SLICE_X76Y106_AQ),
.I1(1'b1),
.I2(CLBLM_R_X49Y104_SLICE_X75Y104_DQ),
.I3(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I4(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X62Y102_SLICE_X92Y102_AO5),
.O6(CLBLM_L_X62Y102_SLICE_X92Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y102_SLICE_X93Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y102_SLICE_X93Y102_DO5),
.O6(CLBLM_L_X62Y102_SLICE_X93Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y102_SLICE_X93Y102_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y102_SLICE_X93Y102_CO5),
.O6(CLBLM_L_X62Y102_SLICE_X93Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y102_SLICE_X93Y102_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y102_SLICE_X93Y102_BO5),
.O6(CLBLM_L_X62Y102_SLICE_X93Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000400faffffff)
  ) CLBLM_L_X62Y102_SLICE_X93Y102_ALUT (
.I0(CLBLM_L_X62Y110_SLICE_X92Y110_DO6),
.I1(CLBLM_R_X59Y102_SLICE_X89Y102_AQ),
.I2(CLBLM_L_X62Y103_SLICE_X92Y103_AQ),
.I3(CLBLM_L_X60Y110_SLICE_X91Y110_AQ),
.I4(CLBLM_L_X62Y106_SLICE_X93Y106_AQ),
.I5(1'b1),
.O5(CLBLM_L_X62Y102_SLICE_X93Y102_AO5),
.O6(CLBLM_L_X62Y102_SLICE_X93Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X62Y103_SLICE_X92Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_R_X59Y99_SLICE_X89Y99_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y103_SLICE_X92Y103_AO6),
.Q(CLBLM_L_X62Y103_SLICE_X92Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y103_SLICE_X92Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y103_SLICE_X92Y103_DO5),
.O6(CLBLM_L_X62Y103_SLICE_X92Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88bb88bb88f3c0)
  ) CLBLM_L_X62Y103_SLICE_X92Y103_CLUT (
.I0(CLBLM_L_X62Y104_SLICE_X92Y104_AQ),
.I1(CLBLM_R_X59Y103_SLICE_X89Y103_CQ),
.I2(CLBLM_L_X60Y105_SLICE_X91Y105_B_XOR),
.I3(CLBLM_L_X60Y101_SLICE_X90Y101_CO6),
.I4(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I5(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.O5(CLBLM_L_X62Y103_SLICE_X92Y103_CO5),
.O6(CLBLM_L_X62Y103_SLICE_X92Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd100c000b3008000)
  ) CLBLM_L_X62Y103_SLICE_X92Y103_BLUT (
.I0(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I1(CLBLM_R_X59Y103_SLICE_X89Y103_CQ),
.I2(CLBLM_L_X60Y102_SLICE_X91Y102_BQ),
.I3(CLBLM_R_X59Y103_SLICE_X89Y103_DQ),
.I4(CLBLM_L_X60Y103_SLICE_X91Y103_AQ),
.I5(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.O5(CLBLM_L_X62Y103_SLICE_X92Y103_BO5),
.O6(CLBLM_L_X62Y103_SLICE_X92Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00ccf0ccf0)
  ) CLBLM_L_X62Y103_SLICE_X92Y103_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X49Y104_SLICE_X75Y104_BQ),
.I2(CLBLM_L_X60Y108_SLICE_X91Y108_BO6),
.I3(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I4(CLBLM_L_X62Y103_SLICE_X92Y103_CO6),
.I5(CLBLM_R_X59Y103_SLICE_X89Y103_DQ),
.O5(CLBLM_L_X62Y103_SLICE_X92Y103_AO5),
.O6(CLBLM_L_X62Y103_SLICE_X92Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y103_SLICE_X93Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y100_SLICE_X92Y100_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y103_SLICE_X93Y103_AO5),
.Q(CLBLM_L_X62Y103_SLICE_X93Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y103_SLICE_X93Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y103_SLICE_X93Y103_DO5),
.O6(CLBLM_L_X62Y103_SLICE_X93Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y103_SLICE_X93Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y103_SLICE_X93Y103_CO5),
.O6(CLBLM_L_X62Y103_SLICE_X93Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa548855aa5488)
  ) CLBLM_L_X62Y103_SLICE_X93Y103_BLUT (
.I0(CLBLM_L_X60Y110_SLICE_X91Y110_AQ),
.I1(CLBLM_L_X62Y104_SLICE_X93Y104_AQ),
.I2(CLBLM_R_X59Y102_SLICE_X88Y102_AQ),
.I3(CLBLM_R_X59Y102_SLICE_X89Y102_AQ),
.I4(CLBLM_L_X62Y103_SLICE_X92Y103_AQ),
.I5(1'b1),
.O5(CLBLM_L_X62Y103_SLICE_X93Y103_BO5),
.O6(CLBLM_L_X62Y103_SLICE_X93Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0cc00e2e2e2e2)
  ) CLBLM_L_X62Y103_SLICE_X93Y103_ALUT (
.I0(CLBLM_R_X63Y110_SLICE_X94Y110_CO6),
.I1(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I2(CLBLM_L_X50Y105_SLICE_X77Y105_AQ),
.I3(CLBLM_R_X49Y104_SLICE_X75Y104_AQ),
.I4(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X62Y103_SLICE_X93Y103_AO5),
.O6(CLBLM_L_X62Y103_SLICE_X93Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y104_SLICE_X92Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y102_SLICE_X92Y102_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y104_SLICE_X92Y104_AO6),
.Q(CLBLM_L_X62Y104_SLICE_X92Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y104_SLICE_X92Y104_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y102_SLICE_X92Y102_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y104_SLICE_X92Y104_BO6),
.Q(CLBLM_L_X62Y104_SLICE_X92Y104_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5ccf5ccf0ccffcc)
  ) CLBLM_L_X62Y104_SLICE_X92Y104_DLUT (
.I0(CLBLM_L_X62Y104_SLICE_X92Y104_BQ),
.I1(CLBLM_L_X60Y104_SLICE_X90Y104_CO6),
.I2(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I3(CLBLM_L_X62Y106_SLICE_X93Y106_CO6),
.I4(CLBLM_L_X62Y107_SLICE_X92Y107_A5Q),
.I5(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.O5(CLBLM_L_X62Y104_SLICE_X92Y104_DO5),
.O6(CLBLM_L_X62Y104_SLICE_X92Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffdfddfcffdfddff)
  ) CLBLM_L_X62Y104_SLICE_X92Y104_CLUT (
.I0(CLBLM_L_X60Y104_SLICE_X91Y104_AQ),
.I1(CLBLM_R_X59Y103_SLICE_X89Y103_DQ),
.I2(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I3(CLBLM_R_X59Y103_SLICE_X89Y103_CQ),
.I4(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I5(CLBLM_R_X59Y99_SLICE_X88Y99_BQ),
.O5(CLBLM_L_X62Y104_SLICE_X92Y104_CO5),
.O6(CLBLM_L_X62Y104_SLICE_X92Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaeefafafa)
  ) CLBLM_L_X62Y104_SLICE_X92Y104_BLUT (
.I0(CLBLM_L_X62Y106_SLICE_X93Y106_BO5),
.I1(CLBLM_L_X60Y103_SLICE_X91Y103_A_XOR),
.I2(CLBLM_L_X60Y106_SLICE_X91Y106_A_XOR),
.I3(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I4(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I5(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.O5(CLBLM_L_X62Y104_SLICE_X92Y104_BO5),
.O6(CLBLM_L_X62Y104_SLICE_X92Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00bfffff0080)
  ) CLBLM_L_X62Y104_SLICE_X92Y104_ALUT (
.I0(CLBLM_L_X60Y102_SLICE_X91Y102_B_XOR),
.I1(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I2(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I3(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I4(CLBLM_L_X62Y105_SLICE_X92Y105_AO6),
.I5(CLBLM_L_X60Y105_SLICE_X91Y105_B_XOR),
.O5(CLBLM_L_X62Y104_SLICE_X92Y104_AO5),
.O6(CLBLM_L_X62Y104_SLICE_X92Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X62Y104_SLICE_X93Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_R_X59Y99_SLICE_X89Y99_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y104_SLICE_X93Y104_AO6),
.Q(CLBLM_L_X62Y104_SLICE_X93Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y104_SLICE_X93Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y104_SLICE_X93Y104_DO5),
.O6(CLBLM_L_X62Y104_SLICE_X93Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y104_SLICE_X93Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y104_SLICE_X93Y104_CO5),
.O6(CLBLM_L_X62Y104_SLICE_X93Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y104_SLICE_X93Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y104_SLICE_X93Y104_BO5),
.O6(CLBLM_L_X62Y104_SLICE_X93Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88d8d8dd88d8d8)
  ) CLBLM_L_X62Y104_SLICE_X93Y104_ALUT (
.I0(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I1(CLBLM_R_X49Y104_SLICE_X75Y104_AQ),
.I2(CLBLM_R_X59Y107_SLICE_X88Y107_AO6),
.I3(CLBLM_L_X60Y104_SLICE_X90Y104_BO6),
.I4(CLBLM_R_X59Y103_SLICE_X89Y103_DQ),
.I5(1'b1),
.O5(CLBLM_L_X62Y104_SLICE_X93Y104_AO5),
.O6(CLBLM_L_X62Y104_SLICE_X93Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y105_SLICE_X92Y105_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y100_SLICE_X92Y100_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y105_SLICE_X92Y105_CO6),
.Q(CLBLM_L_X62Y105_SLICE_X92Y105_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3300fbc833007340)
  ) CLBLM_L_X62Y105_SLICE_X92Y105_DLUT (
.I0(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I1(CLBLM_L_X62Y106_SLICE_X93Y106_CO6),
.I2(CLBLM_L_X60Y108_SLICE_X90Y108_BQ),
.I3(CLBLM_R_X59Y105_SLICE_X89Y105_DO6),
.I4(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I5(CLBLM_L_X62Y106_SLICE_X92Y106_BQ),
.O5(CLBLM_L_X62Y105_SLICE_X92Y105_DO5),
.O6(CLBLM_L_X62Y105_SLICE_X92Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf808fd0dfd0df808)
  ) CLBLM_L_X62Y105_SLICE_X92Y105_CLUT (
.I0(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I1(CLBLM_L_X62Y105_SLICE_X93Y105_AO5),
.I2(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I3(CLBLM_L_X50Y104_SLICE_X76Y104_AQ),
.I4(CLBLM_L_X62Y105_SLICE_X92Y105_BO5),
.I5(CLBLM_L_X62Y105_SLICE_X92Y105_CQ),
.O5(CLBLM_L_X62Y105_SLICE_X92Y105_CO5),
.O6(CLBLM_L_X62Y105_SLICE_X92Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefffea000a000)
  ) CLBLM_L_X62Y105_SLICE_X92Y105_BLUT (
.I0(CLBLM_R_X59Y101_SLICE_X89Y101_AQ),
.I1(CLBLL_R_X57Y102_SLICE_X86Y102_BQ),
.I2(CLBLL_R_X57Y102_SLICE_X86Y102_AQ),
.I3(CLBLM_R_X59Y103_SLICE_X89Y103_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y105_SLICE_X92Y105_BO5),
.O6(CLBLM_L_X62Y105_SLICE_X92Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888a0a0dd88dd88)
  ) CLBLM_L_X62Y105_SLICE_X92Y105_ALUT (
.I0(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I1(CLBLM_R_X49Y105_SLICE_X75Y105_CQ),
.I2(CLBLM_R_X49Y104_SLICE_X75Y104_BQ),
.I3(CLBLM_L_X64Y109_SLICE_X96Y109_CO6),
.I4(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X62Y105_SLICE_X92Y105_AO5),
.O6(CLBLM_L_X62Y105_SLICE_X92Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y105_SLICE_X93Y105_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y100_SLICE_X92Y100_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y105_SLICE_X93Y105_BO6),
.Q(CLBLM_L_X62Y105_SLICE_X93Y105_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0a03020f0a03020)
  ) CLBLM_L_X62Y105_SLICE_X93Y105_DLUT (
.I0(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I1(CLBLM_R_X49Y119_SLICE_X74Y119_BQ),
.I2(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I3(CLBLM_L_X62Y105_SLICE_X92Y105_BO6),
.I4(CLBLM_R_X49Y119_SLICE_X74Y119_AQ),
.I5(1'b1),
.O5(CLBLM_L_X62Y105_SLICE_X93Y105_DO5),
.O6(CLBLM_L_X62Y105_SLICE_X93Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcf4f8f00c040800)
  ) CLBLM_L_X62Y105_SLICE_X93Y105_CLUT (
.I0(CLBLM_L_X62Y105_SLICE_X93Y105_AO6),
.I1(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I2(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I3(CLBLM_R_X63Y106_SLICE_X95Y106_A_XOR),
.I4(CLBLM_R_X63Y106_SLICE_X94Y106_B_XOR),
.I5(CLBLM_L_X50Y106_SLICE_X76Y106_CQ),
.O5(CLBLM_L_X62Y105_SLICE_X93Y105_CO5),
.O6(CLBLM_L_X62Y105_SLICE_X93Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff000a000c)
  ) CLBLM_L_X62Y105_SLICE_X93Y105_BLUT (
.I0(CLBLM_R_X63Y106_SLICE_X95Y106_A_XOR),
.I1(CLBLM_L_X62Y105_SLICE_X93Y105_BQ),
.I2(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I3(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I4(CLBLM_L_X62Y105_SLICE_X92Y105_BO5),
.I5(CLBLM_L_X62Y105_SLICE_X93Y105_CO6),
.O5(CLBLM_L_X62Y105_SLICE_X93Y105_BO5),
.O6(CLBLM_L_X62Y105_SLICE_X93Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f000000a3aaaaaa)
  ) CLBLM_L_X62Y105_SLICE_X93Y105_ALUT (
.I0(CLBLM_R_X63Y105_SLICE_X94Y105_A_XOR),
.I1(CLBLM_L_X62Y105_SLICE_X92Y105_CQ),
.I2(CLBLM_R_X59Y103_SLICE_X89Y103_A5Q),
.I3(CLBLM_R_X59Y101_SLICE_X89Y101_AQ),
.I4(CLBLL_R_X57Y102_SLICE_X86Y102_AQ),
.I5(1'b1),
.O5(CLBLM_L_X62Y105_SLICE_X93Y105_AO5),
.O6(CLBLM_L_X62Y105_SLICE_X93Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y106_SLICE_X92Y106_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y102_SLICE_X92Y102_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y106_SLICE_X92Y106_BO6),
.Q(CLBLM_L_X62Y106_SLICE_X92Y106_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y106_SLICE_X92Y106_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y102_SLICE_X92Y102_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y106_SLICE_X92Y106_CO6),
.Q(CLBLM_L_X62Y106_SLICE_X92Y106_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffc0300aaaaaaaa)
  ) CLBLM_L_X62Y106_SLICE_X92Y106_DLUT (
.I0(CLBLM_L_X62Y106_SLICE_X92Y106_AO6),
.I1(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I2(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I3(CLBLM_L_X60Y106_SLICE_X91Y106_A_XOR),
.I4(CLBLM_L_X62Y104_SLICE_X92Y104_BQ),
.I5(CLBLM_R_X59Y103_SLICE_X89Y103_CQ),
.O5(CLBLM_L_X62Y106_SLICE_X92Y106_DO5),
.O6(CLBLM_L_X62Y106_SLICE_X92Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f1f5f5f4f0f0f0)
  ) CLBLM_L_X62Y106_SLICE_X92Y106_CLUT (
.I0(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I1(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I2(CLBLM_L_X62Y107_SLICE_X92Y107_BO5),
.I3(CLBLM_L_X60Y103_SLICE_X91Y103_C_XOR),
.I4(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I5(CLBLM_L_X60Y106_SLICE_X91Y106_C_XOR),
.O5(CLBLM_L_X62Y106_SLICE_X92Y106_CO5),
.O6(CLBLM_L_X62Y106_SLICE_X92Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbabbaaabaabbaa)
  ) CLBLM_L_X62Y106_SLICE_X92Y106_BLUT (
.I0(CLBLM_L_X62Y108_SLICE_X92Y108_BO5),
.I1(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I2(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I3(CLBLM_L_X60Y106_SLICE_X91Y106_B_XOR),
.I4(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I5(CLBLM_L_X60Y103_SLICE_X91Y103_B_XOR),
.O5(CLBLM_L_X62Y106_SLICE_X92Y106_BO5),
.O6(CLBLM_L_X62Y106_SLICE_X92Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacccccf000f000)
  ) CLBLM_L_X62Y106_SLICE_X92Y106_ALUT (
.I0(CLBLM_L_X60Y106_SLICE_X90Y106_B_XOR),
.I1(CLBLM_R_X59Y112_SLICE_X89Y112_AQ),
.I2(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I3(CLBLM_R_X59Y103_SLICE_X89Y103_CQ),
.I4(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I5(1'b1),
.O5(CLBLM_L_X62Y106_SLICE_X92Y106_AO5),
.O6(CLBLM_L_X62Y106_SLICE_X92Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X62Y106_SLICE_X93Y106_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_R_X59Y99_SLICE_X89Y99_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y106_SLICE_X93Y106_AO6),
.Q(CLBLM_L_X62Y106_SLICE_X93Y106_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h44444444ee4ee444)
  ) CLBLM_L_X62Y106_SLICE_X93Y106_DLUT (
.I0(CLBLM_L_X62Y106_SLICE_X93Y106_CO6),
.I1(CLBLM_L_X62Y107_SLICE_X92Y107_DO6),
.I2(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I3(CLBLM_L_X62Y106_SLICE_X92Y106_CQ),
.I4(CLBLM_L_X62Y107_SLICE_X92Y107_BQ),
.I5(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.O5(CLBLM_L_X62Y106_SLICE_X93Y106_DO5),
.O6(CLBLM_L_X62Y106_SLICE_X93Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00040040fe8cfec8)
  ) CLBLM_L_X62Y106_SLICE_X93Y106_CLUT (
.I0(CLBLM_L_X62Y104_SLICE_X93Y104_AQ),
.I1(CLBLM_L_X60Y110_SLICE_X91Y110_AQ),
.I2(CLBLM_R_X59Y102_SLICE_X88Y102_AQ),
.I3(CLBLM_R_X59Y102_SLICE_X89Y102_AQ),
.I4(CLBLM_L_X62Y106_SLICE_X93Y106_AQ),
.I5(CLBLM_L_X62Y103_SLICE_X92Y103_AQ),
.O5(CLBLM_L_X62Y106_SLICE_X93Y106_CO5),
.O6(CLBLM_L_X62Y106_SLICE_X93Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c00000c0c0f000)
  ) CLBLM_L_X62Y106_SLICE_X93Y106_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X50Y106_SLICE_X76Y106_CQ),
.I2(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I3(CLBLM_R_X49Y106_SLICE_X75Y106_CQ),
.I4(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X62Y106_SLICE_X93Y106_BO5),
.O6(CLBLM_L_X62Y106_SLICE_X93Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfef40e04fef40e04)
  ) CLBLM_L_X62Y106_SLICE_X93Y106_ALUT (
.I0(CLBLM_R_X59Y103_SLICE_X89Y103_DQ),
.I1(CLBLM_R_X59Y110_SLICE_X89Y110_CO6),
.I2(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I3(CLBLM_L_X62Y106_SLICE_X92Y106_DO6),
.I4(CLBLM_R_X49Y106_SLICE_X75Y106_CQ),
.I5(1'b1),
.O5(CLBLM_L_X62Y106_SLICE_X93Y106_AO5),
.O6(CLBLM_L_X62Y106_SLICE_X93Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y107_SLICE_X92Y107_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y102_SLICE_X92Y102_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y106_SLICE_X93Y106_BO6),
.Q(CLBLM_L_X62Y107_SLICE_X92Y107_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y107_SLICE_X92Y107_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y102_SLICE_X92Y102_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y107_SLICE_X92Y107_AO6),
.Q(CLBLM_L_X62Y107_SLICE_X92Y107_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X62Y107_SLICE_X92Y107_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y102_SLICE_X92Y102_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y107_SLICE_X92Y107_BO6),
.Q(CLBLM_L_X62Y107_SLICE_X92Y107_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3bbc0bbf388c088)
  ) CLBLM_L_X62Y107_SLICE_X92Y107_DLUT (
.I0(CLBLM_L_X60Y107_SLICE_X91Y107_AQ),
.I1(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I2(CLBLM_R_X59Y100_SLICE_X89Y100_DQ),
.I3(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I4(CLBLM_R_X59Y106_SLICE_X89Y106_BQ),
.I5(CLBLM_R_X59Y96_SLICE_X89Y96_A5Q),
.O5(CLBLM_L_X62Y107_SLICE_X92Y107_DO5),
.O6(CLBLM_L_X62Y107_SLICE_X92Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hce020000e2220000)
  ) CLBLM_L_X62Y107_SLICE_X92Y107_CLUT (
.I0(CLBLM_L_X60Y106_SLICE_X90Y106_AQ),
.I1(CLBLM_R_X59Y103_SLICE_X89Y103_CQ),
.I2(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I3(CLBLM_L_X62Y107_SLICE_X92Y107_A5Q),
.I4(CLBLM_R_X59Y103_SLICE_X89Y103_DQ),
.I5(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.O5(CLBLM_L_X62Y107_SLICE_X92Y107_CO5),
.O6(CLBLM_L_X62Y107_SLICE_X92Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc000000cc00aa00)
  ) CLBLM_L_X62Y107_SLICE_X92Y107_BLUT (
.I0(CLBLM_R_X49Y107_SLICE_X75Y107_CQ),
.I1(CLBLM_L_X50Y107_SLICE_X77Y107_AQ),
.I2(1'b1),
.I3(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I4(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X62Y107_SLICE_X92Y107_BO5),
.O6(CLBLM_L_X62Y107_SLICE_X92Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccf0aaaaaa)
  ) CLBLM_L_X62Y107_SLICE_X92Y107_ALUT (
.I0(CLBLM_L_X60Y107_SLICE_X91Y107_B_XOR),
.I1(CLBLM_L_X62Y100_SLICE_X93Y100_AO6),
.I2(CLBLM_L_X60Y104_SLICE_X91Y104_B_XOR),
.I3(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I4(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I5(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.O5(CLBLM_L_X62Y107_SLICE_X92Y107_AO5),
.O6(CLBLM_L_X62Y107_SLICE_X92Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y107_SLICE_X93Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y107_SLICE_X93Y107_DO5),
.O6(CLBLM_L_X62Y107_SLICE_X93Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaff2222aaff7777)
  ) CLBLM_L_X62Y107_SLICE_X93Y107_CLUT (
.I0(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I1(CLBLM_L_X64Y105_SLICE_X97Y105_AQ),
.I2(1'b1),
.I3(CLBLM_R_X49Y111_SLICE_X74Y111_BQ),
.I4(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I5(CLBLM_L_X64Y107_SLICE_X97Y107_AQ),
.O5(CLBLM_L_X62Y107_SLICE_X93Y107_CO5),
.O6(CLBLM_L_X62Y107_SLICE_X93Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc3344f3008a44ba)
  ) CLBLM_L_X62Y107_SLICE_X93Y107_BLUT (
.I0(CLBLM_L_X60Y110_SLICE_X91Y110_AQ),
.I1(CLBLM_R_X59Y102_SLICE_X89Y102_AQ),
.I2(CLBLM_L_X62Y106_SLICE_X93Y106_AQ),
.I3(CLBLM_L_X62Y104_SLICE_X93Y104_AQ),
.I4(CLBLM_L_X62Y103_SLICE_X92Y103_AQ),
.I5(CLBLM_R_X59Y102_SLICE_X88Y102_AQ),
.O5(CLBLM_L_X62Y107_SLICE_X93Y107_BO5),
.O6(CLBLM_L_X62Y107_SLICE_X93Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f6f6fb383b3b3)
  ) CLBLM_L_X62Y107_SLICE_X93Y107_ALUT (
.I0(CLBLM_L_X60Y110_SLICE_X91Y110_AQ),
.I1(CLBLM_R_X59Y102_SLICE_X89Y102_AQ),
.I2(CLBLM_L_X62Y106_SLICE_X93Y106_AQ),
.I3(CLBLM_L_X62Y104_SLICE_X93Y104_AQ),
.I4(CLBLM_L_X62Y103_SLICE_X92Y103_AQ),
.I5(CLBLM_R_X59Y102_SLICE_X88Y102_AQ),
.O5(CLBLM_L_X62Y107_SLICE_X93Y107_AO5),
.O6(CLBLM_L_X62Y107_SLICE_X93Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X62Y108_SLICE_X92Y108_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_R_X59Y99_SLICE_X89Y99_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y108_SLICE_X92Y108_AO5),
.Q(CLBLM_L_X62Y108_SLICE_X92Y108_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X62Y108_SLICE_X92Y108_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_R_X59Y99_SLICE_X89Y99_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y108_SLICE_X92Y108_AO6),
.Q(CLBLM_L_X62Y108_SLICE_X92Y108_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y108_SLICE_X92Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y108_SLICE_X92Y108_DO5),
.O6(CLBLM_L_X62Y108_SLICE_X92Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc85fc80000000000)
  ) CLBLM_L_X62Y108_SLICE_X92Y108_CLUT (
.I0(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I1(CLBLM_L_X60Y108_SLICE_X90Y108_BQ),
.I2(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I3(CLBLM_R_X59Y103_SLICE_X89Y103_CQ),
.I4(CLBLM_R_X59Y108_SLICE_X89Y108_AQ),
.I5(CLBLM_R_X59Y103_SLICE_X89Y103_DQ),
.O5(CLBLM_L_X62Y108_SLICE_X92Y108_CO5),
.O6(CLBLM_L_X62Y108_SLICE_X92Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a00000aaa00a00)
  ) CLBLM_L_X62Y108_SLICE_X92Y108_BLUT (
.I0(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I1(1'b1),
.I2(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I3(CLBLM_R_X49Y106_SLICE_X75Y106_DQ),
.I4(CLBLM_L_X50Y107_SLICE_X76Y107_BQ),
.I5(1'b1),
.O5(CLBLM_L_X62Y108_SLICE_X92Y108_BO5),
.O6(CLBLM_L_X62Y108_SLICE_X92Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5500555551515151)
  ) CLBLM_L_X62Y108_SLICE_X92Y108_ALUT (
.I0(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I1(CLBLM_R_X59Y105_SLICE_X88Y105_CO6),
.I2(CLBLM_L_X62Y107_SLICE_X92Y107_CO6),
.I3(CLBLM_L_X62Y103_SLICE_X92Y103_BO6),
.I4(CLBLM_L_X62Y104_SLICE_X92Y104_CO6),
.I5(1'b1),
.O5(CLBLM_L_X62Y108_SLICE_X92Y108_AO5),
.O6(CLBLM_L_X62Y108_SLICE_X92Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X62Y108_SLICE_X93Y108_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_R_X59Y99_SLICE_X89Y99_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y108_SLICE_X93Y108_AO6),
.Q(CLBLM_L_X62Y108_SLICE_X93Y108_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44cccccccc)
  ) CLBLM_L_X62Y108_SLICE_X93Y108_DLUT (
.I0(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I1(CLBLM_R_X59Y106_SLICE_X89Y106_BQ),
.I2(1'b1),
.I3(CLBLM_L_X60Y106_SLICE_X90Y106_D_XOR),
.I4(1'b1),
.I5(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.O5(CLBLM_L_X62Y108_SLICE_X93Y108_DO5),
.O6(CLBLM_L_X62Y108_SLICE_X93Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0df8fd080)
  ) CLBLM_L_X62Y108_SLICE_X93Y108_CLUT (
.I0(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I1(CLBLM_L_X62Y106_SLICE_X92Y106_CQ),
.I2(CLBLM_R_X59Y103_SLICE_X89Y103_CQ),
.I3(CLBLM_L_X60Y106_SLICE_X91Y106_C_XOR),
.I4(CLBLM_L_X62Y108_SLICE_X93Y108_DO6),
.I5(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.O5(CLBLM_L_X62Y108_SLICE_X93Y108_CO5),
.O6(CLBLM_L_X62Y108_SLICE_X93Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8080a280a2802200)
  ) CLBLM_L_X62Y108_SLICE_X93Y108_BLUT (
.I0(CLBLM_R_X59Y103_SLICE_X89Y103_DQ),
.I1(CLBLM_R_X59Y103_SLICE_X89Y103_CQ),
.I2(CLBLM_L_X62Y107_SLICE_X92Y107_BQ),
.I3(CLBLM_L_X60Y107_SLICE_X91Y107_AQ),
.I4(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I5(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.O5(CLBLM_L_X62Y108_SLICE_X93Y108_BO5),
.O6(CLBLM_L_X62Y108_SLICE_X93Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0eef0eef022f022)
  ) CLBLM_L_X62Y108_SLICE_X93Y108_ALUT (
.I0(CLBLM_R_X59Y107_SLICE_X88Y107_CO6),
.I1(CLBLM_R_X59Y103_SLICE_X89Y103_DQ),
.I2(CLBLM_R_X49Y107_SLICE_X75Y107_CQ),
.I3(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I4(1'b1),
.I5(CLBLM_L_X62Y108_SLICE_X93Y108_CO6),
.O5(CLBLM_L_X62Y108_SLICE_X93Y108_AO5),
.O6(CLBLM_L_X62Y108_SLICE_X93Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y109_SLICE_X92Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y109_SLICE_X92Y109_DO5),
.O6(CLBLM_L_X62Y109_SLICE_X92Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffff7ff)
  ) CLBLM_L_X62Y109_SLICE_X92Y109_CLUT (
.I0(CLBLM_L_X62Y103_SLICE_X92Y103_AQ),
.I1(CLBLM_L_X62Y106_SLICE_X93Y106_AQ),
.I2(CLBLM_L_X62Y104_SLICE_X93Y104_AQ),
.I3(CLBLM_L_X60Y110_SLICE_X91Y110_AQ),
.I4(CLBLM_L_X62Y110_SLICE_X92Y110_DO6),
.I5(CLBLM_R_X59Y102_SLICE_X89Y102_AQ),
.O5(CLBLM_L_X62Y109_SLICE_X92Y109_CO5),
.O6(CLBLM_L_X62Y109_SLICE_X92Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aa00c000ea00)
  ) CLBLM_L_X62Y109_SLICE_X92Y109_BLUT (
.I0(CLBLL_R_X57Y102_SLICE_X86Y102_AQ),
.I1(CLBLM_L_X60Y98_SLICE_X90Y98_BQ),
.I2(CLBLM_R_X59Y102_SLICE_X88Y102_AQ),
.I3(CLBLM_L_X56Y103_SLICE_X85Y103_CO6),
.I4(CLBLL_R_X57Y102_SLICE_X86Y102_BQ),
.I5(CLBLM_L_X62Y109_SLICE_X92Y109_CO6),
.O5(CLBLM_L_X62Y109_SLICE_X92Y109_BO5),
.O6(CLBLM_L_X62Y109_SLICE_X92Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeff02fffe000200)
  ) CLBLM_L_X62Y109_SLICE_X92Y109_ALUT (
.I0(CLBLM_L_X60Y107_SLICE_X91Y107_B_XOR),
.I1(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I2(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I3(CLBLM_R_X59Y103_SLICE_X89Y103_CQ),
.I4(CLBLM_L_X62Y107_SLICE_X92Y107_AQ),
.I5(CLBLM_L_X60Y110_SLICE_X91Y110_CO6),
.O5(CLBLM_L_X62Y109_SLICE_X92Y109_AO5),
.O6(CLBLM_L_X62Y109_SLICE_X92Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y109_SLICE_X93Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y109_SLICE_X93Y109_DO5),
.O6(CLBLM_L_X62Y109_SLICE_X93Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y109_SLICE_X93Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y109_SLICE_X93Y109_CO5),
.O6(CLBLM_L_X62Y109_SLICE_X93Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y109_SLICE_X93Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y109_SLICE_X93Y109_BO5),
.O6(CLBLM_L_X62Y109_SLICE_X93Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y109_SLICE_X93Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y109_SLICE_X93Y109_AO5),
.O6(CLBLM_L_X62Y109_SLICE_X93Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X62Y110_SLICE_X92Y110_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_R_X59Y99_SLICE_X89Y99_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y110_SLICE_X92Y110_AO6),
.Q(CLBLM_L_X62Y110_SLICE_X92Y110_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X62Y110_SLICE_X92Y110_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_R_X59Y99_SLICE_X89Y99_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y110_SLICE_X92Y110_BO6),
.Q(CLBLM_L_X62Y110_SLICE_X92Y110_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff5fffffffffffff)
  ) CLBLM_L_X62Y110_SLICE_X92Y110_DLUT (
.I0(CLBLM_L_X62Y108_SLICE_X92Y108_AQ),
.I1(1'b1),
.I2(CLBLM_L_X62Y110_SLICE_X92Y110_BQ),
.I3(CLBLM_L_X62Y111_SLICE_X92Y111_CO6),
.I4(CLBLM_L_X62Y108_SLICE_X93Y108_AQ),
.I5(CLBLM_L_X60Y111_SLICE_X91Y111_AQ),
.O5(CLBLM_L_X62Y110_SLICE_X92Y110_DO5),
.O6(CLBLM_L_X62Y110_SLICE_X92Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000e2ffe200)
  ) CLBLM_L_X62Y110_SLICE_X92Y110_CLUT (
.I0(CLBLM_L_X60Y106_SLICE_X91Y106_B_XOR),
.I1(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I2(CLBLM_L_X62Y106_SLICE_X92Y106_BQ),
.I3(CLBLM_R_X59Y103_SLICE_X89Y103_CQ),
.I4(CLBLM_L_X60Y110_SLICE_X91Y110_DO6),
.I5(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.O5(CLBLM_L_X62Y110_SLICE_X92Y110_CO5),
.O6(CLBLM_L_X62Y110_SLICE_X92Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccaaffaa00)
  ) CLBLM_L_X62Y110_SLICE_X92Y110_BLUT (
.I0(CLBLM_L_X62Y109_SLICE_X92Y109_AO6),
.I1(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.I2(1'b1),
.I3(CLBLM_R_X59Y103_SLICE_X89Y103_DQ),
.I4(CLBLM_R_X59Y110_SLICE_X89Y110_BO6),
.I5(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.O5(CLBLM_L_X62Y110_SLICE_X92Y110_BO5),
.O6(CLBLM_L_X62Y110_SLICE_X92Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcacfcac0cac0ca)
  ) CLBLM_L_X62Y110_SLICE_X92Y110_ALUT (
.I0(CLBLM_R_X59Y112_SLICE_X89Y112_CO6),
.I1(CLBLM_R_X49Y106_SLICE_X75Y106_DQ),
.I2(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I3(CLBLM_R_X59Y103_SLICE_X89Y103_DQ),
.I4(1'b1),
.I5(CLBLM_L_X62Y110_SLICE_X92Y110_CO6),
.O5(CLBLM_L_X62Y110_SLICE_X92Y110_AO5),
.O6(CLBLM_L_X62Y110_SLICE_X92Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X62Y110_SLICE_X93Y110_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y110_SLICE_X93Y110_AO6),
.Q(CLBLM_L_X62Y110_SLICE_X93Y110_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y110_SLICE_X93Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y110_SLICE_X93Y110_DO5),
.O6(CLBLM_L_X62Y110_SLICE_X93Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000aaaaaaaa)
  ) CLBLM_L_X62Y110_SLICE_X93Y110_CLUT (
.I0(CLBLM_R_X49Y119_SLICE_X74Y119_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X49Y119_SLICE_X74Y119_AQ),
.O5(CLBLM_L_X62Y110_SLICE_X93Y110_CO5),
.O6(CLBLM_L_X62Y110_SLICE_X93Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8282414100820041)
  ) CLBLM_L_X62Y110_SLICE_X93Y110_BLUT (
.I0(CLBLL_R_X57Y99_SLICE_X87Y99_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(CLBLM_L_X62Y110_SLICE_X93Y110_AQ),
.I3(CLBLM_R_X49Y119_SLICE_X74Y119_BQ),
.I4(LIOB33_X0Y121_IOB_X0Y122_I),
.I5(CLBLM_R_X49Y119_SLICE_X74Y119_AQ),
.O5(CLBLM_L_X62Y110_SLICE_X93Y110_BO5),
.O6(CLBLM_L_X62Y110_SLICE_X93Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ccccf0f08800)
  ) CLBLM_L_X62Y110_SLICE_X93Y110_ALUT (
.I0(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I1(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I2(CLBLM_L_X62Y110_SLICE_X93Y110_AQ),
.I3(CLBLM_L_X62Y105_SLICE_X92Y105_BO6),
.I4(CLBLM_L_X62Y110_SLICE_X93Y110_CO6),
.I5(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.O5(CLBLM_L_X62Y110_SLICE_X93Y110_AO5),
.O6(CLBLM_L_X62Y110_SLICE_X93Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X62Y111_SLICE_X92Y111_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_R_X59Y99_SLICE_X89Y99_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y111_SLICE_X92Y111_AO5),
.Q(CLBLM_L_X62Y111_SLICE_X92Y111_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X62Y111_SLICE_X92Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_R_X59Y99_SLICE_X89Y99_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y111_SLICE_X92Y111_AO6),
.Q(CLBLM_L_X62Y111_SLICE_X92Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f7fffffffffffff)
  ) CLBLM_L_X62Y111_SLICE_X92Y111_DLUT (
.I0(CLBLM_L_X62Y110_SLICE_X92Y110_BQ),
.I1(CLBLM_L_X60Y111_SLICE_X90Y111_AQ),
.I2(CLBLM_L_X62Y108_SLICE_X93Y108_AQ),
.I3(1'b1),
.I4(CLBLM_L_X62Y110_SLICE_X92Y110_AQ),
.I5(CLBLM_L_X60Y111_SLICE_X91Y111_BQ),
.O5(CLBLM_L_X62Y111_SLICE_X92Y111_DO5),
.O6(CLBLM_L_X62Y111_SLICE_X92Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffffffffffffff)
  ) CLBLM_L_X62Y111_SLICE_X92Y111_CLUT (
.I0(CLBLM_L_X60Y111_SLICE_X91Y111_BQ),
.I1(CLBLM_L_X62Y111_SLICE_X92Y111_AQ),
.I2(CLBLM_L_X60Y111_SLICE_X90Y111_AQ),
.I3(CLBLM_L_X62Y111_SLICE_X92Y111_A5Q),
.I4(CLBLM_L_X62Y110_SLICE_X92Y110_AQ),
.I5(CLBLM_L_X62Y108_SLICE_X92Y108_A5Q),
.O5(CLBLM_L_X62Y111_SLICE_X92Y111_CO5),
.O6(CLBLM_L_X62Y111_SLICE_X92Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfffffffffffffff)
  ) CLBLM_L_X62Y111_SLICE_X92Y111_BLUT (
.I0(CLBLM_L_X62Y111_SLICE_X92Y111_DO6),
.I1(CLBLM_L_X60Y111_SLICE_X91Y111_AQ),
.I2(CLBLM_L_X62Y111_SLICE_X92Y111_AQ),
.I3(CLBLM_L_X62Y108_SLICE_X92Y108_A5Q),
.I4(CLBLM_L_X62Y108_SLICE_X92Y108_AQ),
.I5(CLBLM_L_X62Y111_SLICE_X92Y111_A5Q),
.O5(CLBLM_L_X62Y111_SLICE_X92Y111_BO5),
.O6(CLBLM_L_X62Y111_SLICE_X92Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0f0c0f0f0f0505)
  ) CLBLM_L_X62Y111_SLICE_X92Y111_ALUT (
.I0(CLBLM_L_X60Y112_SLICE_X90Y112_BO6),
.I1(CLBLM_L_X62Y108_SLICE_X92Y108_CO6),
.I2(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I3(CLBLM_L_X60Y112_SLICE_X90Y112_AO6),
.I4(CLBLM_L_X62Y108_SLICE_X93Y108_BO6),
.I5(1'b1),
.O5(CLBLM_L_X62Y111_SLICE_X92Y111_AO5),
.O6(CLBLM_L_X62Y111_SLICE_X92Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y111_SLICE_X93Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y111_SLICE_X93Y111_DO5),
.O6(CLBLM_L_X62Y111_SLICE_X93Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y111_SLICE_X93Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y111_SLICE_X93Y111_CO5),
.O6(CLBLM_L_X62Y111_SLICE_X93Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y111_SLICE_X93Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y111_SLICE_X93Y111_BO5),
.O6(CLBLM_L_X62Y111_SLICE_X93Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y111_SLICE_X93Y111_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y111_SLICE_X93Y111_AO5),
.O6(CLBLM_L_X62Y111_SLICE_X93Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X62Y112_SLICE_X92Y112_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y110_SLICE_X93Y110_BO6),
.D(CLBLM_L_X62Y112_SLICE_X92Y112_AO6),
.PRE(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.Q(CLBLM_L_X62Y112_SLICE_X92Y112_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y112_SLICE_X92Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y112_SLICE_X92Y112_DO5),
.O6(CLBLM_L_X62Y112_SLICE_X92Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y112_SLICE_X92Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y112_SLICE_X92Y112_CO5),
.O6(CLBLM_L_X62Y112_SLICE_X92Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y112_SLICE_X92Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y112_SLICE_X92Y112_BO5),
.O6(CLBLM_L_X62Y112_SLICE_X92Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0f0f0f)
  ) CLBLM_L_X62Y112_SLICE_X92Y112_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y112_SLICE_X92Y112_AO5),
.O6(CLBLM_L_X62Y112_SLICE_X92Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y112_SLICE_X93Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y112_SLICE_X93Y112_DO5),
.O6(CLBLM_L_X62Y112_SLICE_X93Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y112_SLICE_X93Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y112_SLICE_X93Y112_CO5),
.O6(CLBLM_L_X62Y112_SLICE_X93Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y112_SLICE_X93Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y112_SLICE_X93Y112_BO5),
.O6(CLBLM_L_X62Y112_SLICE_X93Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X62Y112_SLICE_X93Y112_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X62Y112_SLICE_X93Y112_AO5),
.O6(CLBLM_L_X62Y112_SLICE_X93Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y95_SLICE_X97Y95_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y95_SLICE_X97Y95_DO5),
.O6(CLBLM_L_X64Y95_SLICE_X97Y95_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y95_SLICE_X97Y95_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y95_SLICE_X97Y95_CO5),
.O6(CLBLM_L_X64Y95_SLICE_X97Y95_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y95_SLICE_X97Y95_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y95_SLICE_X97Y95_BO5),
.O6(CLBLM_L_X64Y95_SLICE_X97Y95_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y95_SLICE_X97Y95_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y95_SLICE_X97Y95_AO5),
.O6(CLBLM_L_X64Y95_SLICE_X97Y95_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y96_SLICE_X97Y96_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y99_SLICE_X93Y99_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X64Y96_SLICE_X97Y96_AO6),
.Q(CLBLM_L_X64Y96_SLICE_X97Y96_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y96_SLICE_X97Y96_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y99_SLICE_X93Y99_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X64Y96_SLICE_X97Y96_BO6),
.Q(CLBLM_L_X64Y96_SLICE_X97Y96_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y96_SLICE_X97Y96_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y99_SLICE_X93Y99_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X64Y96_SLICE_X97Y96_CO6),
.Q(CLBLM_L_X64Y96_SLICE_X97Y96_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y96_SLICE_X97Y96_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y99_SLICE_X93Y99_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X64Y96_SLICE_X97Y96_DO6),
.Q(CLBLM_L_X64Y96_SLICE_X97Y96_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55fa50aa00fa50)
  ) CLBLM_L_X64Y96_SLICE_X97Y96_DLUT (
.I0(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I1(1'b1),
.I2(CLBLM_L_X64Y96_SLICE_X96Y96_BO5),
.I3(CLBLM_L_X50Y104_SLICE_X76Y104_AQ),
.I4(CLBLM_L_X56Y98_SLICE_X85Y98_DQ),
.I5(CLBLM_R_X63Y98_SLICE_X95Y98_AQ),
.O5(CLBLM_L_X64Y96_SLICE_X97Y96_DO5),
.O6(CLBLM_L_X64Y96_SLICE_X97Y96_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50ee44fa50ee44)
  ) CLBLM_L_X64Y96_SLICE_X97Y96_CLUT (
.I0(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I1(CLBLM_L_X64Y96_SLICE_X96Y96_CO6),
.I2(CLBLM_L_X64Y97_SLICE_X96Y97_A5Q),
.I3(CLBLM_R_X49Y106_SLICE_X74Y106_AQ),
.I4(CLBLM_L_X56Y98_SLICE_X85Y98_DQ),
.I5(1'b1),
.O5(CLBLM_L_X64Y96_SLICE_X97Y96_CO5),
.O6(CLBLM_L_X64Y96_SLICE_X97Y96_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffd8d80000d8d8)
  ) CLBLM_L_X64Y96_SLICE_X97Y96_BLUT (
.I0(CLBLM_L_X56Y98_SLICE_X85Y98_DQ),
.I1(CLBLM_L_X64Y97_SLICE_X96Y97_AQ),
.I2(CLBLM_L_X64Y96_SLICE_X96Y96_CO5),
.I3(1'b1),
.I4(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I5(CLBLM_R_X49Y105_SLICE_X75Y105_CQ),
.O5(CLBLM_L_X64Y96_SLICE_X97Y96_BO5),
.O6(CLBLM_L_X64Y96_SLICE_X97Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffee440000ee44)
  ) CLBLM_L_X64Y96_SLICE_X97Y96_ALUT (
.I0(CLBLM_L_X56Y98_SLICE_X85Y98_DQ),
.I1(CLBLM_L_X64Y96_SLICE_X96Y96_BO6),
.I2(1'b1),
.I3(CLBLM_R_X63Y98_SLICE_X95Y98_A5Q),
.I4(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I5(CLBLM_L_X50Y105_SLICE_X77Y105_AQ),
.O5(CLBLM_L_X64Y96_SLICE_X97Y96_AO5),
.O6(CLBLM_L_X64Y96_SLICE_X97Y96_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X64Y97_SLICE_X96Y97_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X64Y97_SLICE_X96Y97_AO5),
.Q(CLBLM_L_X64Y97_SLICE_X96Y97_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X64Y97_SLICE_X96Y97_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X64Y97_SLICE_X96Y97_BO5),
.Q(CLBLM_L_X64Y97_SLICE_X96Y97_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X64Y97_SLICE_X96Y97_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X64Y97_SLICE_X96Y97_AO6),
.Q(CLBLM_L_X64Y97_SLICE_X96Y97_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X64Y97_SLICE_X96Y97_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X64Y97_SLICE_X96Y97_BO6),
.Q(CLBLM_L_X64Y97_SLICE_X96Y97_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y97_SLICE_X96Y97_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y97_SLICE_X96Y97_DO5),
.O6(CLBLM_L_X64Y97_SLICE_X96Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ff5000000000)
  ) CLBLM_L_X64Y97_SLICE_X96Y97_CLUT (
.I0(CLBLM_L_X64Y96_SLICE_X97Y96_AQ),
.I1(1'b1),
.I2(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I3(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I4(CLBLM_L_X56Y97_SLICE_X85Y97_AQ),
.I5(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.O5(CLBLM_L_X64Y97_SLICE_X96Y97_CO5),
.O6(CLBLM_L_X64Y97_SLICE_X96Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a0dd88dd88)
  ) CLBLM_L_X64Y97_SLICE_X96Y97_BLUT (
.I0(CLBLM_R_X63Y99_SLICE_X94Y99_DO5),
.I1(CLBLM_L_X62Y97_SLICE_X92Y97_BQ),
.I2(CLBLM_L_X62Y97_SLICE_X92Y97_AQ),
.I3(CLBLM_R_X65Y104_SLICE_X99Y104_BQ),
.I4(CLBLM_R_X65Y103_SLICE_X99Y103_BQ),
.I5(1'b1),
.O5(CLBLM_L_X64Y97_SLICE_X96Y97_BO5),
.O6(CLBLM_L_X64Y97_SLICE_X96Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00aaf0aaf0)
  ) CLBLM_L_X64Y97_SLICE_X96Y97_ALUT (
.I0(CLBLM_R_X63Y97_SLICE_X95Y97_D5Q),
.I1(CLBLM_R_X63Y97_SLICE_X95Y97_DQ),
.I2(CLBLM_L_X64Y99_SLICE_X96Y99_AQ),
.I3(CLBLM_R_X63Y99_SLICE_X94Y99_DO5),
.I4(CLBLM_R_X65Y102_SLICE_X99Y102_AQ),
.I5(1'b1),
.O5(CLBLM_L_X64Y97_SLICE_X96Y97_AO5),
.O6(CLBLM_L_X64Y97_SLICE_X96Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y97_SLICE_X97Y97_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y99_SLICE_X93Y99_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X64Y97_SLICE_X97Y97_AO6),
.Q(CLBLM_L_X64Y97_SLICE_X97Y97_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y97_SLICE_X97Y97_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y99_SLICE_X93Y99_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X64Y97_SLICE_X97Y97_BO6),
.Q(CLBLM_L_X64Y97_SLICE_X97Y97_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y97_SLICE_X97Y97_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y97_SLICE_X97Y97_DO5),
.O6(CLBLM_L_X64Y97_SLICE_X97Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000f0c00000c0c0)
  ) CLBLM_L_X64Y97_SLICE_X97Y97_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I2(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I3(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I4(CLBLM_L_X56Y97_SLICE_X85Y97_AQ),
.I5(CLBLM_R_X63Y95_SLICE_X95Y95_AQ),
.O5(CLBLM_L_X64Y97_SLICE_X97Y97_CO5),
.O6(CLBLM_L_X64Y97_SLICE_X97Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacfcac0cacfcac0)
  ) CLBLM_L_X64Y97_SLICE_X97Y97_BLUT (
.I0(CLBLM_R_X63Y99_SLICE_X95Y99_AQ),
.I1(CLBLM_L_X50Y107_SLICE_X76Y107_BQ),
.I2(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I3(CLBLM_L_X56Y98_SLICE_X85Y98_DQ),
.I4(CLBLM_R_X63Y96_SLICE_X94Y96_BO5),
.I5(1'b1),
.O5(CLBLM_L_X64Y97_SLICE_X97Y97_BO5),
.O6(CLBLM_L_X64Y97_SLICE_X97Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa3afa3aca0aca0)
  ) CLBLM_L_X64Y97_SLICE_X97Y97_ALUT (
.I0(CLBLM_L_X50Y106_SLICE_X76Y106_AQ),
.I1(CLBLM_L_X56Y98_SLICE_X85Y98_DQ),
.I2(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I3(CLBLM_R_X63Y98_SLICE_X95Y98_BQ),
.I4(1'b1),
.I5(CLBLM_R_X63Y96_SLICE_X94Y96_AO5),
.O5(CLBLM_L_X64Y97_SLICE_X97Y97_AO5),
.O6(CLBLM_L_X64Y97_SLICE_X97Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X64Y98_SLICE_X96Y98_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_BQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X64Y98_SLICE_X96Y98_AO6),
.Q(CLBLM_L_X64Y98_SLICE_X96Y98_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h80002000f0f0f0f0)
  ) CLBLM_L_X64Y98_SLICE_X96Y98_DLUT (
.I0(CLBLM_L_X60Y98_SLICE_X90Y98_AQ),
.I1(CLBLM_L_X62Y100_SLICE_X92Y100_AQ),
.I2(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I3(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I4(CLBLM_R_X65Y100_SLICE_X99Y100_CQ),
.I5(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.O5(CLBLM_L_X64Y98_SLICE_X96Y98_DO5),
.O6(CLBLM_L_X64Y98_SLICE_X96Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffbb0000f7b3)
  ) CLBLM_L_X64Y98_SLICE_X96Y98_CLUT (
.I0(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I1(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I2(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I3(CLBLM_L_X64Y100_SLICE_X97Y100_A_XOR),
.I4(CLBLM_L_X64Y98_SLICE_X96Y98_DO6),
.I5(CLBLM_L_X62Y100_SLICE_X92Y100_AQ),
.O5(CLBLM_L_X64Y98_SLICE_X96Y98_CO5),
.O6(CLBLM_L_X64Y98_SLICE_X96Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00dc0000ffdcff00)
  ) CLBLM_L_X64Y98_SLICE_X96Y98_BLUT (
.I0(CLBLM_R_X63Y95_SLICE_X95Y95_DQ),
.I1(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I2(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I3(CLBLM_L_X56Y97_SLICE_X85Y97_AQ),
.I4(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I5(CLBLM_L_X64Y98_SLICE_X96Y98_CO6),
.O5(CLBLM_L_X64Y98_SLICE_X96Y98_BO5),
.O6(CLBLM_L_X64Y98_SLICE_X96Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0c0e0e0c000e00)
  ) CLBLM_L_X64Y98_SLICE_X96Y98_ALUT (
.I0(CLBLM_R_X63Y101_SLICE_X95Y101_DO6),
.I1(CLBLM_R_X65Y97_SLICE_X98Y97_AO6),
.I2(CLBLM_L_X64Y97_SLICE_X96Y97_CO6),
.I3(CLBLM_L_X64Y101_SLICE_X96Y101_D_XOR),
.I4(CLBLM_R_X65Y98_SLICE_X98Y98_DO6),
.I5(CLBLM_R_X65Y97_SLICE_X98Y97_AO5),
.O5(CLBLM_L_X64Y98_SLICE_X96Y98_AO5),
.O6(CLBLM_L_X64Y98_SLICE_X96Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X64Y98_SLICE_X97Y98_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_BQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X64Y98_SLICE_X97Y98_AO6),
.Q(CLBLM_L_X64Y98_SLICE_X97Y98_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff3bfb3fff3bfb3)
  ) CLBLM_L_X64Y98_SLICE_X97Y98_DLUT (
.I0(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I1(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I2(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I3(CLBLM_L_X64Y101_SLICE_X97Y101_D_XOR),
.I4(CLBLM_L_X62Y101_SLICE_X93Y101_CQ),
.I5(1'b1),
.O5(CLBLM_L_X64Y98_SLICE_X97Y98_DO5),
.O6(CLBLM_L_X64Y98_SLICE_X97Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33330000bb330000)
  ) CLBLM_L_X64Y98_SLICE_X97Y98_CLUT (
.I0(CLBLM_L_X60Y98_SLICE_X90Y98_AQ),
.I1(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I2(1'b1),
.I3(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I4(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I5(CLBLM_R_X65Y101_SLICE_X98Y101_D_XOR),
.O5(CLBLM_L_X64Y98_SLICE_X97Y98_CO5),
.O6(CLBLM_L_X64Y98_SLICE_X97Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3010301030003000)
  ) CLBLM_L_X64Y98_SLICE_X97Y98_BLUT (
.I0(CLBLM_L_X64Y96_SLICE_X97Y96_DQ),
.I1(CLBLM_L_X56Y97_SLICE_X85Y97_AQ),
.I2(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I3(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I4(1'b1),
.I5(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.O5(CLBLM_L_X64Y98_SLICE_X97Y98_BO5),
.O6(CLBLM_L_X64Y98_SLICE_X97Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00e000e000ee00e0)
  ) CLBLM_L_X64Y98_SLICE_X97Y98_ALUT (
.I0(CLBLM_L_X64Y101_SLICE_X96Y101_C_XOR),
.I1(CLBLM_R_X65Y97_SLICE_X98Y97_AO5),
.I2(CLBLM_R_X65Y97_SLICE_X98Y97_AO6),
.I3(CLBLM_L_X64Y98_SLICE_X97Y98_BO6),
.I4(CLBLM_L_X64Y98_SLICE_X97Y98_DO6),
.I5(CLBLM_L_X64Y98_SLICE_X97Y98_CO6),
.O5(CLBLM_L_X64Y98_SLICE_X97Y98_AO5),
.O6(CLBLM_L_X64Y98_SLICE_X97Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X64Y99_SLICE_X96Y99_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_BQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X64Y99_SLICE_X96Y99_AO6),
.Q(CLBLM_L_X64Y99_SLICE_X96Y99_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X64Y99_SLICE_X96Y99_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_BQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X64Y99_SLICE_X96Y99_BO6),
.Q(CLBLM_L_X64Y99_SLICE_X96Y99_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55005500f5005500)
  ) CLBLM_L_X64Y99_SLICE_X96Y99_DLUT (
.I0(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I1(1'b1),
.I2(CLBLM_L_X60Y98_SLICE_X90Y98_AQ),
.I3(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I4(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I5(CLBLM_R_X65Y101_SLICE_X98Y101_C_XOR),
.O5(CLBLM_L_X64Y99_SLICE_X96Y99_DO5),
.O6(CLBLM_L_X64Y99_SLICE_X96Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2200220022202220)
  ) CLBLM_L_X64Y99_SLICE_X96Y99_CLUT (
.I0(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I1(CLBLM_L_X56Y97_SLICE_X85Y97_AQ),
.I2(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I3(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I4(1'b1),
.I5(CLBLM_L_X64Y96_SLICE_X97Y96_CQ),
.O5(CLBLM_L_X64Y99_SLICE_X96Y99_CO5),
.O6(CLBLM_L_X64Y99_SLICE_X96Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000fcfc00005400)
  ) CLBLM_L_X64Y99_SLICE_X96Y99_BLUT (
.I0(CLBLM_L_X64Y99_SLICE_X96Y99_DO6),
.I1(CLBLM_L_X64Y101_SLICE_X96Y101_B_XOR),
.I2(CLBLM_R_X65Y97_SLICE_X98Y97_AO5),
.I3(CLBLM_L_X64Y99_SLICE_X97Y99_CO6),
.I4(CLBLM_R_X65Y96_SLICE_X98Y96_BO6),
.I5(CLBLM_R_X65Y97_SLICE_X98Y97_AO6),
.O5(CLBLM_L_X64Y99_SLICE_X96Y99_BO5),
.O6(CLBLM_L_X64Y99_SLICE_X96Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ff22f020)
  ) CLBLM_L_X64Y99_SLICE_X96Y99_ALUT (
.I0(CLBLM_R_X63Y101_SLICE_X95Y101_CO6),
.I1(CLBLM_L_X64Y99_SLICE_X97Y99_BO6),
.I2(CLBLM_R_X65Y97_SLICE_X98Y97_AO5),
.I3(CLBLM_R_X65Y97_SLICE_X98Y97_AO6),
.I4(CLBLM_L_X64Y102_SLICE_X96Y102_B_XOR),
.I5(CLBLM_L_X64Y99_SLICE_X96Y99_CO6),
.O5(CLBLM_L_X64Y99_SLICE_X96Y99_AO5),
.O6(CLBLM_L_X64Y99_SLICE_X96Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X64Y99_SLICE_X97Y99_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_BQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X64Y99_SLICE_X97Y99_AO6),
.Q(CLBLM_L_X64Y99_SLICE_X97Y99_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cc000000fc0000)
  ) CLBLM_L_X64Y99_SLICE_X97Y99_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I2(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I3(CLBLM_L_X56Y97_SLICE_X85Y97_AQ),
.I4(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I5(CLBLM_L_X64Y96_SLICE_X97Y96_BQ),
.O5(CLBLM_L_X64Y99_SLICE_X97Y99_DO5),
.O6(CLBLM_L_X64Y99_SLICE_X97Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hefefefefef2fef2f)
  ) CLBLM_L_X64Y99_SLICE_X97Y99_CLUT (
.I0(CLBLM_L_X64Y101_SLICE_X97Y101_C_XOR),
.I1(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I2(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I3(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I4(1'b1),
.I5(CLBLM_L_X62Y101_SLICE_X93Y101_BQ),
.O5(CLBLM_L_X64Y99_SLICE_X97Y99_CO5),
.O6(CLBLM_L_X64Y99_SLICE_X97Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f8f8f00000000)
  ) CLBLM_L_X64Y99_SLICE_X97Y99_BLUT (
.I0(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I1(CLBLM_L_X60Y98_SLICE_X90Y98_AQ),
.I2(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I3(1'b1),
.I4(CLBLM_R_X65Y102_SLICE_X98Y102_C_XOR),
.I5(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.O5(CLBLM_L_X64Y99_SLICE_X97Y99_BO5),
.O6(CLBLM_L_X64Y99_SLICE_X97Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff4f4fffff444f)
  ) CLBLM_L_X64Y99_SLICE_X97Y99_ALUT (
.I0(CLBLM_R_X65Y97_SLICE_X98Y97_AO5),
.I1(CLBLM_L_X64Y100_SLICE_X96Y100_C_XOR),
.I2(CLBLM_R_X65Y97_SLICE_X98Y97_AO6),
.I3(CLBLM_R_X63Y100_SLICE_X95Y100_BO6),
.I4(CLBLM_L_X64Y97_SLICE_X97Y97_CO6),
.I5(CLBLM_R_X65Y99_SLICE_X99Y99_DO6),
.O5(CLBLM_L_X64Y99_SLICE_X97Y99_AO5),
.O6(CLBLM_L_X64Y99_SLICE_X97Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X64Y100_SLICE_X96Y100_CARRY4 (
.CI(1'b0),
.CO({CLBLM_L_X64Y100_SLICE_X96Y100_D_CY, CLBLM_L_X64Y100_SLICE_X96Y100_C_CY, CLBLM_L_X64Y100_SLICE_X96Y100_B_CY, CLBLM_L_X64Y100_SLICE_X96Y100_A_CY}),
.CYINIT(CLBLM_R_X65Y100_SLICE_X99Y100_CQ),
.DI({1'b0, 1'b0, 1'b0, CLBLM_L_X64Y100_SLICE_X96Y100_AO5}),
.O({CLBLM_L_X64Y100_SLICE_X96Y100_D_XOR, CLBLM_L_X64Y100_SLICE_X96Y100_C_XOR, CLBLM_L_X64Y100_SLICE_X96Y100_B_XOR, CLBLM_L_X64Y100_SLICE_X96Y100_A_XOR}),
.S({CLBLM_L_X64Y100_SLICE_X96Y100_DO6, CLBLM_L_X64Y100_SLICE_X96Y100_CO6, CLBLM_L_X64Y100_SLICE_X96Y100_BO6, CLBLM_L_X64Y100_SLICE_X96Y100_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X64Y100_SLICE_X96Y100_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X65Y100_SLICE_X99Y100_BQ),
.O5(CLBLM_L_X64Y100_SLICE_X96Y100_DO5),
.O6(CLBLM_L_X64Y100_SLICE_X96Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X64Y100_SLICE_X96Y100_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X64Y106_SLICE_X97Y106_DQ),
.O5(CLBLM_L_X64Y100_SLICE_X96Y100_CO5),
.O6(CLBLM_L_X64Y100_SLICE_X96Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X64Y100_SLICE_X96Y100_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X65Y106_SLICE_X98Y106_CQ),
.O5(CLBLM_L_X64Y100_SLICE_X96Y100_BO5),
.O6(CLBLM_L_X64Y100_SLICE_X96Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0000000000)
  ) CLBLM_L_X64Y100_SLICE_X96Y100_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X65Y100_SLICE_X99Y100_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y100_SLICE_X96Y100_AO5),
.O6(CLBLM_L_X64Y100_SLICE_X96Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X64Y100_SLICE_X97Y100_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y101_SLICE_X93Y101_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X64Y100_SLICE_X97Y100_AO5),
.Q(CLBLM_L_X64Y100_SLICE_X97Y100_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X64Y100_SLICE_X97Y100_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y101_SLICE_X93Y101_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X64Y100_SLICE_X97Y100_BO5),
.Q(CLBLM_L_X64Y100_SLICE_X97Y100_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X64Y100_SLICE_X97Y100_CARRY4 (
.CI(1'b0),
.CO({CLBLM_L_X64Y100_SLICE_X97Y100_D_CY, CLBLM_L_X64Y100_SLICE_X97Y100_C_CY, CLBLM_L_X64Y100_SLICE_X97Y100_B_CY, CLBLM_L_X64Y100_SLICE_X97Y100_A_CY}),
.CYINIT(1'b0),
.DI({CLBLM_L_X64Y106_SLICE_X97Y106_DQ, CLBLM_R_X65Y106_SLICE_X98Y106_CQ, CLBLM_R_X65Y100_SLICE_X99Y100_AQ, CLBLM_R_X65Y100_SLICE_X99Y100_CQ}),
.O({CLBLM_L_X64Y100_SLICE_X97Y100_D_XOR, CLBLM_L_X64Y100_SLICE_X97Y100_C_XOR, CLBLM_L_X64Y100_SLICE_X97Y100_B_XOR, CLBLM_L_X64Y100_SLICE_X97Y100_A_XOR}),
.S({CLBLM_L_X64Y100_SLICE_X97Y100_DO6, CLBLM_L_X64Y100_SLICE_X97Y100_CO6, CLBLM_L_X64Y100_SLICE_X97Y100_BO6, CLBLM_L_X64Y100_SLICE_X97Y100_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6666666666666666)
  ) CLBLM_L_X64Y100_SLICE_X97Y100_DLUT (
.I0(CLBLM_L_X64Y106_SLICE_X97Y106_DQ),
.I1(CLBLM_L_X62Y100_SLICE_X92Y100_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y100_SLICE_X97Y100_DO5),
.O6(CLBLM_L_X64Y100_SLICE_X97Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5a5a5a5a5a)
  ) CLBLM_L_X64Y100_SLICE_X97Y100_CLUT (
.I0(CLBLM_L_X62Y101_SLICE_X93Y101_AQ),
.I1(1'b1),
.I2(CLBLM_R_X65Y106_SLICE_X98Y106_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y100_SLICE_X97Y100_CO5),
.O6(CLBLM_L_X64Y100_SLICE_X97Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cc33ccf0f0f0f0)
  ) CLBLM_L_X64Y100_SLICE_X97Y100_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X65Y100_SLICE_X99Y100_AQ),
.I2(CLBLM_R_X49Y106_SLICE_X75Y106_CQ),
.I3(CLBLM_L_X62Y100_SLICE_X92Y100_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y100_SLICE_X97Y100_BO5),
.O6(CLBLM_L_X64Y100_SLICE_X97Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5aff00ff00)
  ) CLBLM_L_X64Y100_SLICE_X97Y100_ALUT (
.I0(CLBLM_R_X65Y100_SLICE_X99Y100_CQ),
.I1(1'b1),
.I2(CLBLM_L_X62Y100_SLICE_X92Y100_AQ),
.I3(CLBLM_R_X49Y104_SLICE_X75Y104_DQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y100_SLICE_X97Y100_AO5),
.O6(CLBLM_L_X64Y100_SLICE_X97Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X64Y101_SLICE_X96Y101_CARRY4 (
.CI(CLBLM_L_X64Y100_SLICE_X96Y100_COUT),
.CO({CLBLM_L_X64Y101_SLICE_X96Y101_D_CY, CLBLM_L_X64Y101_SLICE_X96Y101_C_CY, CLBLM_L_X64Y101_SLICE_X96Y101_B_CY, CLBLM_L_X64Y101_SLICE_X96Y101_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_L_X64Y101_SLICE_X96Y101_D_XOR, CLBLM_L_X64Y101_SLICE_X96Y101_C_XOR, CLBLM_L_X64Y101_SLICE_X96Y101_B_XOR, CLBLM_L_X64Y101_SLICE_X96Y101_A_XOR}),
.S({CLBLM_L_X64Y101_SLICE_X96Y101_DO6, CLBLM_L_X64Y101_SLICE_X96Y101_CO6, CLBLM_L_X64Y101_SLICE_X96Y101_BO6, CLBLM_L_X64Y101_SLICE_X96Y101_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X64Y101_SLICE_X96Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X63Y103_SLICE_X95Y103_CQ),
.O5(CLBLM_L_X64Y101_SLICE_X96Y101_DO5),
.O6(CLBLM_L_X64Y101_SLICE_X96Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X64Y101_SLICE_X96Y101_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X63Y101_SLICE_X95Y101_AQ),
.O5(CLBLM_L_X64Y101_SLICE_X96Y101_CO5),
.O6(CLBLM_L_X64Y101_SLICE_X96Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X64Y101_SLICE_X96Y101_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X63Y103_SLICE_X95Y103_BQ),
.O5(CLBLM_L_X64Y101_SLICE_X96Y101_BO5),
.O6(CLBLM_L_X64Y101_SLICE_X96Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X64Y101_SLICE_X96Y101_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X65Y106_SLICE_X98Y106_DQ),
.O5(CLBLM_L_X64Y101_SLICE_X96Y101_AO5),
.O6(CLBLM_L_X64Y101_SLICE_X96Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X64Y101_SLICE_X97Y101_CARRY4 (
.CI(CLBLM_L_X64Y100_SLICE_X97Y100_COUT),
.CO({CLBLM_L_X64Y101_SLICE_X97Y101_D_CY, CLBLM_L_X64Y101_SLICE_X97Y101_C_CY, CLBLM_L_X64Y101_SLICE_X97Y101_B_CY, CLBLM_L_X64Y101_SLICE_X97Y101_A_CY}),
.CYINIT(1'b0),
.DI({CLBLM_R_X63Y101_SLICE_X95Y101_AQ, CLBLM_R_X63Y103_SLICE_X95Y103_BQ, CLBLM_R_X65Y106_SLICE_X98Y106_DQ, CLBLM_R_X65Y100_SLICE_X99Y100_BQ}),
.O({CLBLM_L_X64Y101_SLICE_X97Y101_D_XOR, CLBLM_L_X64Y101_SLICE_X97Y101_C_XOR, CLBLM_L_X64Y101_SLICE_X97Y101_B_XOR, CLBLM_L_X64Y101_SLICE_X97Y101_A_XOR}),
.S({CLBLM_L_X64Y101_SLICE_X97Y101_DO6, CLBLM_L_X64Y101_SLICE_X97Y101_CO6, CLBLM_L_X64Y101_SLICE_X97Y101_BO6, CLBLM_L_X64Y101_SLICE_X97Y101_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333333cccccccc)
  ) CLBLM_L_X64Y101_SLICE_X97Y101_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X62Y101_SLICE_X93Y101_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X63Y101_SLICE_X95Y101_AQ),
.O5(CLBLM_L_X64Y101_SLICE_X97Y101_DO5),
.O6(CLBLM_L_X64Y101_SLICE_X97Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555555aaaaaaaa)
  ) CLBLM_L_X64Y101_SLICE_X97Y101_CLUT (
.I0(CLBLM_R_X63Y103_SLICE_X95Y103_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X62Y101_SLICE_X93Y101_BQ),
.O5(CLBLM_L_X64Y101_SLICE_X97Y101_CO5),
.O6(CLBLM_L_X64Y101_SLICE_X97Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3c3c3c3c3c)
  ) CLBLM_L_X64Y101_SLICE_X97Y101_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X65Y106_SLICE_X98Y106_DQ),
.I2(CLBLM_L_X64Y100_SLICE_X97Y100_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y101_SLICE_X97Y101_BO5),
.O6(CLBLM_L_X64Y101_SLICE_X97Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff00ff00ff00ff0)
  ) CLBLM_L_X64Y101_SLICE_X97Y101_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X64Y100_SLICE_X97Y100_AQ),
.I3(CLBLM_R_X65Y100_SLICE_X99Y100_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y101_SLICE_X97Y101_AO5),
.O6(CLBLM_L_X64Y101_SLICE_X97Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X64Y102_SLICE_X96Y102_CARRY4 (
.CI(CLBLM_L_X64Y101_SLICE_X96Y101_COUT),
.CO({CLBLM_L_X64Y102_SLICE_X96Y102_D_CY, CLBLM_L_X64Y102_SLICE_X96Y102_C_CY, CLBLM_L_X64Y102_SLICE_X96Y102_B_CY, CLBLM_L_X64Y102_SLICE_X96Y102_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_L_X64Y102_SLICE_X96Y102_D_XOR, CLBLM_L_X64Y102_SLICE_X96Y102_C_XOR, CLBLM_L_X64Y102_SLICE_X96Y102_B_XOR, CLBLM_L_X64Y102_SLICE_X96Y102_A_XOR}),
.S({CLBLM_L_X64Y102_SLICE_X96Y102_DO6, CLBLM_L_X64Y102_SLICE_X96Y102_CO6, CLBLM_L_X64Y102_SLICE_X96Y102_BO6, CLBLM_L_X64Y102_SLICE_X96Y102_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X64Y102_SLICE_X96Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X65Y107_SLICE_X98Y107_CQ),
.O5(CLBLM_L_X64Y102_SLICE_X96Y102_DO5),
.O6(CLBLM_L_X64Y102_SLICE_X96Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X64Y102_SLICE_X96Y102_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X65Y107_SLICE_X98Y107_BQ),
.O5(CLBLM_L_X64Y102_SLICE_X96Y102_CO5),
.O6(CLBLM_L_X64Y102_SLICE_X96Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X64Y102_SLICE_X96Y102_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X65Y107_SLICE_X98Y107_AQ),
.O5(CLBLM_L_X64Y102_SLICE_X96Y102_BO5),
.O6(CLBLM_L_X64Y102_SLICE_X96Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X64Y102_SLICE_X96Y102_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X65Y107_SLICE_X98Y107_DQ),
.O5(CLBLM_L_X64Y102_SLICE_X96Y102_AO5),
.O6(CLBLM_L_X64Y102_SLICE_X96Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X64Y102_SLICE_X97Y102_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y101_SLICE_X93Y101_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X64Y102_SLICE_X97Y102_AO5),
.Q(CLBLM_L_X64Y102_SLICE_X97Y102_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X64Y102_SLICE_X97Y102_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y101_SLICE_X93Y101_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X64Y102_SLICE_X97Y102_BO5),
.Q(CLBLM_L_X64Y102_SLICE_X97Y102_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X64Y102_SLICE_X97Y102_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y101_SLICE_X93Y101_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X64Y102_SLICE_X97Y102_CO5),
.Q(CLBLM_L_X64Y102_SLICE_X97Y102_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X64Y102_SLICE_X97Y102_CARRY4 (
.CI(CLBLM_L_X64Y101_SLICE_X97Y101_COUT),
.CO({CLBLM_L_X64Y102_SLICE_X97Y102_D_CY, CLBLM_L_X64Y102_SLICE_X97Y102_C_CY, CLBLM_L_X64Y102_SLICE_X97Y102_B_CY, CLBLM_L_X64Y102_SLICE_X97Y102_A_CY}),
.CYINIT(1'b0),
.DI({CLBLM_L_X64Y102_SLICE_X97Y102_DO5, CLBLM_L_X64Y102_SLICE_X97Y102_AQ, CLBLM_R_X65Y107_SLICE_X98Y107_DQ, CLBLM_R_X63Y103_SLICE_X95Y103_CQ}),
.O({CLBLM_L_X64Y102_SLICE_X97Y102_D_XOR, CLBLM_L_X64Y102_SLICE_X97Y102_C_XOR, CLBLM_L_X64Y102_SLICE_X97Y102_B_XOR, CLBLM_L_X64Y102_SLICE_X97Y102_A_XOR}),
.S({CLBLM_L_X64Y102_SLICE_X97Y102_DO6, CLBLM_L_X64Y102_SLICE_X97Y102_CO6, CLBLM_L_X64Y102_SLICE_X97Y102_BO6, CLBLM_L_X64Y102_SLICE_X97Y102_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555aaaa0000ffff)
  ) CLBLM_L_X64Y102_SLICE_X97Y102_DLUT (
.I0(CLBLM_R_X65Y107_SLICE_X98Y107_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X64Y102_SLICE_X97Y102_AQ),
.I5(1'b1),
.O5(CLBLM_L_X64Y102_SLICE_X97Y102_DO5),
.O6(CLBLM_L_X64Y102_SLICE_X97Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ccccf0f0f0f0)
  ) CLBLM_L_X64Y102_SLICE_X97Y102_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X65Y107_SLICE_X98Y107_AQ),
.I2(CLBLM_R_X49Y107_SLICE_X75Y107_DQ),
.I3(1'b1),
.I4(CLBLM_L_X64Y102_SLICE_X97Y102_AQ),
.I5(1'b1),
.O5(CLBLM_L_X64Y102_SLICE_X97Y102_CO5),
.O6(CLBLM_L_X64Y102_SLICE_X97Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3cffff0000)
  ) CLBLM_L_X64Y102_SLICE_X97Y102_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X65Y107_SLICE_X98Y107_DQ),
.I2(CLBLM_L_X64Y102_SLICE_X97Y102_CQ),
.I3(1'b1),
.I4(CLBLM_R_X49Y108_SLICE_X75Y108_DQ),
.I5(1'b1),
.O5(CLBLM_L_X64Y102_SLICE_X97Y102_BO5),
.O6(CLBLM_L_X64Y102_SLICE_X97Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3cff00ff00)
  ) CLBLM_L_X64Y102_SLICE_X97Y102_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X64Y102_SLICE_X97Y102_BQ),
.I2(CLBLM_R_X63Y103_SLICE_X95Y103_CQ),
.I3(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y102_SLICE_X97Y102_AO5),
.O6(CLBLM_L_X64Y102_SLICE_X97Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X64Y103_SLICE_X96Y103_CARRY4 (
.CI(CLBLM_L_X64Y102_SLICE_X96Y102_COUT),
.CO({CLBLM_L_X64Y103_SLICE_X96Y103_D_CY, CLBLM_L_X64Y103_SLICE_X96Y103_C_CY, CLBLM_L_X64Y103_SLICE_X96Y103_B_CY, CLBLM_L_X64Y103_SLICE_X96Y103_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_L_X64Y103_SLICE_X96Y103_D_XOR, CLBLM_L_X64Y103_SLICE_X96Y103_C_XOR, CLBLM_L_X64Y103_SLICE_X96Y103_B_XOR, CLBLM_L_X64Y103_SLICE_X96Y103_A_XOR}),
.S({CLBLM_L_X64Y103_SLICE_X96Y103_DO6, CLBLM_L_X64Y103_SLICE_X96Y103_CO6, CLBLM_L_X64Y103_SLICE_X96Y103_BO6, CLBLM_L_X64Y103_SLICE_X96Y103_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X64Y103_SLICE_X96Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X65Y106_SLICE_X98Y106_BQ),
.O5(CLBLM_L_X64Y103_SLICE_X96Y103_DO5),
.O6(CLBLM_L_X64Y103_SLICE_X96Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X64Y103_SLICE_X96Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X63Y103_SLICE_X95Y103_AQ),
.O5(CLBLM_L_X64Y103_SLICE_X96Y103_CO5),
.O6(CLBLM_L_X64Y103_SLICE_X96Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X64Y103_SLICE_X96Y103_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X64Y106_SLICE_X97Y106_AQ),
.O5(CLBLM_L_X64Y103_SLICE_X96Y103_BO5),
.O6(CLBLM_L_X64Y103_SLICE_X96Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X64Y103_SLICE_X96Y103_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X65Y106_SLICE_X98Y106_AQ),
.O5(CLBLM_L_X64Y103_SLICE_X96Y103_AO5),
.O6(CLBLM_L_X64Y103_SLICE_X96Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X64Y103_SLICE_X97Y103_CARRY4 (
.CI(CLBLM_L_X64Y102_SLICE_X97Y102_COUT),
.CO({CLBLM_L_X64Y103_SLICE_X97Y103_D_CY, CLBLM_L_X64Y103_SLICE_X97Y103_C_CY, CLBLM_L_X64Y103_SLICE_X97Y103_B_CY, CLBLM_L_X64Y103_SLICE_X97Y103_A_CY}),
.CYINIT(1'b0),
.DI({CLBLM_L_X64Y106_SLICE_X97Y106_AQ, CLBLM_R_X65Y106_SLICE_X98Y106_AQ, CLBLM_R_X65Y107_SLICE_X98Y107_CQ, CLBLM_R_X65Y107_SLICE_X98Y107_BQ}),
.O({CLBLM_L_X64Y103_SLICE_X97Y103_D_XOR, CLBLM_L_X64Y103_SLICE_X97Y103_C_XOR, CLBLM_L_X64Y103_SLICE_X97Y103_B_XOR, CLBLM_L_X64Y103_SLICE_X97Y103_A_XOR}),
.S({CLBLM_L_X64Y103_SLICE_X97Y103_DO6, CLBLM_L_X64Y103_SLICE_X97Y103_CO6, CLBLM_L_X64Y103_SLICE_X97Y103_BO6, CLBLM_L_X64Y103_SLICE_X97Y103_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa55555555)
  ) CLBLM_L_X64Y103_SLICE_X97Y103_DLUT (
.I0(CLBLM_L_X64Y106_SLICE_X97Y106_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X63Y103_SLICE_X95Y103_AQ),
.O5(CLBLM_L_X64Y103_SLICE_X97Y103_DO5),
.O6(CLBLM_L_X64Y103_SLICE_X97Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9999999999999999)
  ) CLBLM_L_X64Y103_SLICE_X97Y103_CLUT (
.I0(CLBLM_L_X64Y106_SLICE_X97Y106_AQ),
.I1(CLBLM_R_X65Y106_SLICE_X98Y106_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y103_SLICE_X97Y103_CO5),
.O6(CLBLM_L_X64Y103_SLICE_X97Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0000ff00ff)
  ) CLBLM_L_X64Y103_SLICE_X97Y103_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X65Y106_SLICE_X98Y106_AQ),
.I4(1'b1),
.I5(CLBLM_R_X65Y107_SLICE_X98Y107_CQ),
.O5(CLBLM_L_X64Y103_SLICE_X97Y103_BO5),
.O6(CLBLM_L_X64Y103_SLICE_X97Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0000ff00ff)
  ) CLBLM_L_X64Y103_SLICE_X97Y103_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X65Y107_SLICE_X98Y107_BQ),
.I4(1'b1),
.I5(CLBLM_R_X65Y107_SLICE_X98Y107_CQ),
.O5(CLBLM_L_X64Y103_SLICE_X97Y103_AO5),
.O6(CLBLM_L_X64Y103_SLICE_X97Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X64Y104_SLICE_X96Y104_CARRY4 (
.CI(CLBLM_L_X64Y103_SLICE_X96Y103_COUT),
.CO({CLBLM_L_X64Y104_SLICE_X96Y104_D_CY, CLBLM_L_X64Y104_SLICE_X96Y104_C_CY, CLBLM_L_X64Y104_SLICE_X96Y104_B_CY, CLBLM_L_X64Y104_SLICE_X96Y104_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_L_X64Y104_SLICE_X96Y104_D_XOR, CLBLM_L_X64Y104_SLICE_X96Y104_C_XOR, CLBLM_L_X64Y104_SLICE_X96Y104_B_XOR, CLBLM_L_X64Y104_SLICE_X96Y104_A_XOR}),
.S({CLBLM_L_X64Y104_SLICE_X96Y104_DO6, CLBLM_L_X64Y104_SLICE_X96Y104_CO6, CLBLM_L_X64Y104_SLICE_X96Y104_BO6, CLBLM_L_X64Y104_SLICE_X96Y104_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y104_SLICE_X96Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y104_SLICE_X96Y104_DO5),
.O6(CLBLM_L_X64Y104_SLICE_X96Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y104_SLICE_X96Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y104_SLICE_X96Y104_CO5),
.O6(CLBLM_L_X64Y104_SLICE_X96Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X64Y104_SLICE_X96Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X64Y106_SLICE_X97Y106_CQ),
.O5(CLBLM_L_X64Y104_SLICE_X96Y104_BO5),
.O6(CLBLM_L_X64Y104_SLICE_X96Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X64Y104_SLICE_X96Y104_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X64Y106_SLICE_X97Y106_BQ),
.O5(CLBLM_L_X64Y104_SLICE_X96Y104_AO5),
.O6(CLBLM_L_X64Y104_SLICE_X96Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X64Y104_SLICE_X97Y104_CARRY4 (
.CI(CLBLM_L_X64Y103_SLICE_X97Y103_COUT),
.CO({CLBLM_L_X64Y104_SLICE_X97Y104_D_CY, CLBLM_L_X64Y104_SLICE_X97Y104_C_CY, CLBLM_L_X64Y104_SLICE_X97Y104_B_CY, CLBLM_L_X64Y104_SLICE_X97Y104_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, CLBLM_R_X65Y106_SLICE_X98Y106_BQ, CLBLM_R_X63Y103_SLICE_X95Y103_AQ}),
.O({CLBLM_L_X64Y104_SLICE_X97Y104_D_XOR, CLBLM_L_X64Y104_SLICE_X97Y104_C_XOR, CLBLM_L_X64Y104_SLICE_X97Y104_B_XOR, CLBLM_L_X64Y104_SLICE_X97Y104_A_XOR}),
.S({CLBLM_L_X64Y104_SLICE_X97Y104_DO6, CLBLM_L_X64Y104_SLICE_X97Y104_CO6, CLBLM_L_X64Y104_SLICE_X97Y104_BO6, CLBLM_L_X64Y104_SLICE_X97Y104_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y104_SLICE_X97Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y104_SLICE_X97Y104_DO5),
.O6(CLBLM_L_X64Y104_SLICE_X97Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc33cc33cc33cc33)
  ) CLBLM_L_X64Y104_SLICE_X97Y104_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X64Y106_SLICE_X97Y106_BQ),
.I2(1'b1),
.I3(CLBLM_L_X64Y106_SLICE_X97Y106_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y104_SLICE_X97Y104_CO5),
.O6(CLBLM_L_X64Y104_SLICE_X97Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc33cc33cc33cc33)
  ) CLBLM_L_X64Y104_SLICE_X97Y104_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X64Y106_SLICE_X97Y106_BQ),
.I2(1'b1),
.I3(CLBLM_R_X65Y106_SLICE_X98Y106_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y104_SLICE_X97Y104_BO5),
.O6(CLBLM_L_X64Y104_SLICE_X97Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc3c3c3c3c3c3c3c3)
  ) CLBLM_L_X64Y104_SLICE_X97Y104_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X65Y106_SLICE_X98Y106_BQ),
.I2(CLBLM_R_X63Y103_SLICE_X95Y103_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y104_SLICE_X97Y104_AO5),
.O6(CLBLM_L_X64Y104_SLICE_X97Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y105_SLICE_X96Y105_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y100_SLICE_X92Y100_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X64Y105_SLICE_X96Y105_AO6),
.Q(CLBLM_L_X64Y105_SLICE_X96Y105_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd0c0cdddd3f3f)
  ) CLBLM_L_X64Y105_SLICE_X96Y105_DLUT (
.I0(CLBLM_R_X49Y111_SLICE_X74Y111_AQ),
.I1(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I2(CLBLM_L_X64Y105_SLICE_X96Y105_AQ),
.I3(1'b1),
.I4(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I5(CLBLM_L_X64Y107_SLICE_X96Y107_BQ),
.O5(CLBLM_L_X64Y105_SLICE_X96Y105_DO5),
.O6(CLBLM_L_X64Y105_SLICE_X96Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaafffff0aaffff)
  ) CLBLM_L_X64Y105_SLICE_X96Y105_CLUT (
.I0(CLBLM_L_X64Y103_SLICE_X97Y103_C_XOR),
.I1(1'b1),
.I2(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I3(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I4(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I5(CLBLM_R_X49Y106_SLICE_X75Y106_DQ),
.O5(CLBLM_L_X64Y105_SLICE_X96Y105_CO5),
.O6(CLBLM_L_X64Y105_SLICE_X96Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd8d8888d8888888)
  ) CLBLM_L_X64Y105_SLICE_X96Y105_BLUT (
.I0(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I1(CLBLM_R_X49Y105_SLICE_X75Y105_CQ),
.I2(CLBLM_L_X62Y105_SLICE_X93Y105_AO6),
.I3(CLBLM_R_X63Y105_SLICE_X95Y105_B_XOR),
.I4(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I5(CLBLM_R_X63Y105_SLICE_X94Y105_C_XOR),
.O5(CLBLM_L_X64Y105_SLICE_X96Y105_BO5),
.O6(CLBLM_L_X64Y105_SLICE_X96Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff54ff00ff10)
  ) CLBLM_L_X64Y105_SLICE_X96Y105_ALUT (
.I0(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I1(CLBLM_L_X62Y105_SLICE_X92Y105_BO5),
.I2(CLBLM_L_X64Y105_SLICE_X96Y105_AQ),
.I3(CLBLM_L_X64Y105_SLICE_X96Y105_BO6),
.I4(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I5(CLBLM_R_X63Y105_SLICE_X95Y105_B_XOR),
.O5(CLBLM_L_X64Y105_SLICE_X96Y105_AO5),
.O6(CLBLM_L_X64Y105_SLICE_X96Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y105_SLICE_X97Y105_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y100_SLICE_X92Y100_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X64Y105_SLICE_X97Y105_AO6),
.Q(CLBLM_L_X64Y105_SLICE_X97Y105_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hefefefefefef2f2f)
  ) CLBLM_L_X64Y105_SLICE_X97Y105_DLUT (
.I0(CLBLM_L_X64Y104_SLICE_X97Y104_C_XOR),
.I1(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I2(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I3(1'b1),
.I4(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I5(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.O5(CLBLM_L_X64Y105_SLICE_X97Y105_DO5),
.O6(CLBLM_L_X64Y105_SLICE_X97Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffddffddf7d5f7d5)
  ) CLBLM_L_X64Y105_SLICE_X97Y105_CLUT (
.I0(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I1(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I2(CLBLM_R_X49Y104_SLICE_X75Y104_DQ),
.I3(CLBLM_L_X64Y103_SLICE_X97Y103_A_XOR),
.I4(1'b1),
.I5(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.O5(CLBLM_L_X64Y105_SLICE_X97Y105_CO5),
.O6(CLBLM_L_X64Y105_SLICE_X97Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hec20fc30ec20cc00)
  ) CLBLM_L_X64Y105_SLICE_X97Y105_BLUT (
.I0(CLBLM_R_X63Y105_SLICE_X95Y105_C_XOR),
.I1(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I2(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I3(CLBLM_R_X49Y106_SLICE_X74Y106_AQ),
.I4(CLBLM_L_X62Y105_SLICE_X93Y105_AO6),
.I5(CLBLM_R_X63Y105_SLICE_X94Y105_D_XOR),
.O5(CLBLM_L_X64Y105_SLICE_X97Y105_BO5),
.O6(CLBLM_L_X64Y105_SLICE_X97Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff22ff00ff30)
  ) CLBLM_L_X64Y105_SLICE_X97Y105_ALUT (
.I0(CLBLM_R_X63Y105_SLICE_X95Y105_C_XOR),
.I1(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I2(CLBLM_L_X64Y105_SLICE_X97Y105_AQ),
.I3(CLBLM_L_X64Y105_SLICE_X97Y105_BO6),
.I4(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I5(CLBLM_L_X62Y105_SLICE_X92Y105_BO5),
.O5(CLBLM_L_X64Y105_SLICE_X97Y105_AO5),
.O6(CLBLM_L_X64Y105_SLICE_X97Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y106_SLICE_X96Y106_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y100_SLICE_X92Y100_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X64Y106_SLICE_X96Y106_AO6),
.Q(CLBLM_L_X64Y106_SLICE_X96Y106_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y106_SLICE_X96Y106_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y100_SLICE_X92Y100_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X64Y106_SLICE_X96Y106_BO6),
.Q(CLBLM_L_X64Y106_SLICE_X96Y106_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0aa882200)
  ) CLBLM_L_X64Y106_SLICE_X96Y106_DLUT (
.I0(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I1(CLBLM_L_X62Y105_SLICE_X93Y105_AO6),
.I2(CLBLM_L_X50Y107_SLICE_X77Y107_AQ),
.I3(CLBLM_R_X63Y106_SLICE_X94Y106_D_XOR),
.I4(CLBLM_R_X63Y106_SLICE_X95Y106_C_XOR),
.I5(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.O5(CLBLM_L_X64Y106_SLICE_X96Y106_DO5),
.O6(CLBLM_L_X64Y106_SLICE_X96Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa3aca0a0a0a0a0)
  ) CLBLM_L_X64Y106_SLICE_X96Y106_CLUT (
.I0(CLBLM_L_X50Y107_SLICE_X76Y107_BQ),
.I1(CLBLM_L_X62Y105_SLICE_X93Y105_AO6),
.I2(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I3(CLBLM_R_X63Y106_SLICE_X95Y106_B_XOR),
.I4(CLBLM_R_X63Y106_SLICE_X94Y106_C_XOR),
.I5(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.O5(CLBLM_L_X64Y106_SLICE_X96Y106_CO5),
.O6(CLBLM_L_X64Y106_SLICE_X96Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00ff0aff0c)
  ) CLBLM_L_X64Y106_SLICE_X96Y106_BLUT (
.I0(CLBLM_R_X63Y106_SLICE_X95Y106_C_XOR),
.I1(CLBLM_L_X64Y106_SLICE_X96Y106_BQ),
.I2(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I3(CLBLM_L_X64Y106_SLICE_X96Y106_DO6),
.I4(CLBLM_L_X62Y105_SLICE_X92Y105_BO5),
.I5(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.O5(CLBLM_L_X64Y106_SLICE_X96Y106_BO5),
.O6(CLBLM_L_X64Y106_SLICE_X96Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0054ffff0010)
  ) CLBLM_L_X64Y106_SLICE_X96Y106_ALUT (
.I0(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I1(CLBLM_L_X62Y105_SLICE_X92Y105_BO5),
.I2(CLBLM_L_X64Y106_SLICE_X96Y106_AQ),
.I3(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I4(CLBLM_L_X64Y106_SLICE_X96Y106_CO6),
.I5(CLBLM_R_X63Y106_SLICE_X95Y106_B_XOR),
.O5(CLBLM_L_X64Y106_SLICE_X96Y106_AO5),
.O6(CLBLM_L_X64Y106_SLICE_X96Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X64Y106_SLICE_X97Y106_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y105_SLICE_X93Y105_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X64Y106_SLICE_X97Y106_AO6),
.Q(CLBLM_L_X64Y106_SLICE_X97Y106_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X64Y106_SLICE_X97Y106_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y105_SLICE_X93Y105_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X64Y106_SLICE_X97Y106_BO6),
.Q(CLBLM_L_X64Y106_SLICE_X97Y106_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X64Y106_SLICE_X97Y106_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y105_SLICE_X93Y105_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X64Y106_SLICE_X97Y106_CO6),
.Q(CLBLM_L_X64Y106_SLICE_X97Y106_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_L_X64Y106_SLICE_X97Y106_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y105_SLICE_X93Y105_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X64Y106_SLICE_X97Y106_DO6),
.Q(CLBLM_L_X64Y106_SLICE_X97Y106_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf775f775a220a220)
  ) CLBLM_L_X64Y106_SLICE_X97Y106_DLUT (
.I0(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I1(CLBLL_R_X57Y103_SLICE_X86Y103_A5Q),
.I2(CLBLM_L_X64Y99_SLICE_X97Y99_AQ),
.I3(CLBLL_R_X57Y103_SLICE_X86Y103_AQ),
.I4(1'b1),
.I5(CLBLM_R_X63Y104_SLICE_X94Y104_BQ),
.O5(CLBLM_L_X64Y106_SLICE_X97Y106_DO5),
.O6(CLBLM_L_X64Y106_SLICE_X97Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8725050d8725050)
  ) CLBLM_L_X64Y106_SLICE_X97Y106_CLUT (
.I0(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I1(CLBLL_R_X57Y103_SLICE_X86Y103_A5Q),
.I2(CLBLM_L_X64Y109_SLICE_X96Y109_A5Q),
.I3(CLBLL_R_X57Y103_SLICE_X86Y103_AQ),
.I4(CLBLM_R_X65Y105_SLICE_X99Y105_AQ),
.I5(1'b1),
.O5(CLBLM_L_X64Y106_SLICE_X97Y106_CO5),
.O6(CLBLM_L_X64Y106_SLICE_X97Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00f0f05500f0f0)
  ) CLBLM_L_X64Y106_SLICE_X97Y106_BLUT (
.I0(CLBLL_R_X57Y103_SLICE_X86Y103_AQ),
.I1(1'b1),
.I2(CLBLM_R_X63Y105_SLICE_X94Y105_AQ),
.I3(CLBLM_R_X65Y105_SLICE_X98Y105_BQ),
.I4(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I5(CLBLL_R_X57Y103_SLICE_X86Y103_A5Q),
.O5(CLBLM_L_X64Y106_SLICE_X97Y106_BO5),
.O6(CLBLM_L_X64Y106_SLICE_X97Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa00f005f500f00)
  ) CLBLM_L_X64Y106_SLICE_X97Y106_ALUT (
.I0(CLBLL_R_X57Y103_SLICE_X86Y103_AQ),
.I1(1'b1),
.I2(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I3(CLBLM_L_X64Y108_SLICE_X96Y108_BQ),
.I4(CLBLM_R_X65Y103_SLICE_X99Y103_AQ),
.I5(CLBLL_R_X57Y103_SLICE_X86Y103_A5Q),
.O5(CLBLM_L_X64Y106_SLICE_X97Y106_AO5),
.O6(CLBLM_L_X64Y106_SLICE_X97Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y107_SLICE_X96Y107_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_R_X63Y100_SLICE_X94Y100_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X64Y107_SLICE_X96Y107_AO6),
.Q(CLBLM_L_X64Y107_SLICE_X96Y107_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y107_SLICE_X96Y107_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_R_X63Y100_SLICE_X94Y100_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X64Y107_SLICE_X96Y107_BO6),
.Q(CLBLM_L_X64Y107_SLICE_X96Y107_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaf0f8f80a000808)
  ) CLBLM_L_X64Y107_SLICE_X96Y107_DLUT (
.I0(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I1(CLBLM_R_X63Y107_SLICE_X94Y107_C_XOR),
.I2(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I3(CLBLM_R_X63Y107_SLICE_X95Y107_B_XOR),
.I4(CLBLM_L_X62Y105_SLICE_X93Y105_AO6),
.I5(CLBLM_R_X49Y105_SLICE_X75Y105_CQ),
.O5(CLBLM_L_X64Y107_SLICE_X96Y107_DO5),
.O6(CLBLM_L_X64Y107_SLICE_X96Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfacc0acc00cc00)
  ) CLBLM_L_X64Y107_SLICE_X96Y107_CLUT (
.I0(CLBLM_R_X63Y107_SLICE_X94Y107_B_XOR),
.I1(CLBLM_L_X50Y105_SLICE_X77Y105_AQ),
.I2(CLBLM_L_X62Y105_SLICE_X93Y105_AO6),
.I3(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I4(CLBLM_R_X63Y107_SLICE_X95Y107_A_XOR),
.I5(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.O5(CLBLM_L_X64Y107_SLICE_X96Y107_CO5),
.O6(CLBLM_L_X64Y107_SLICE_X96Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f5f0f4f0f0f0f4)
  ) CLBLM_L_X64Y107_SLICE_X96Y107_BLUT (
.I0(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I1(CLBLM_L_X64Y107_SLICE_X96Y107_BQ),
.I2(CLBLM_L_X64Y107_SLICE_X96Y107_DO6),
.I3(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I4(CLBLM_L_X62Y105_SLICE_X92Y105_BO5),
.I5(CLBLM_R_X63Y107_SLICE_X95Y107_B_XOR),
.O5(CLBLM_L_X64Y107_SLICE_X96Y107_BO5),
.O6(CLBLM_L_X64Y107_SLICE_X96Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00220030)
  ) CLBLM_L_X64Y107_SLICE_X96Y107_ALUT (
.I0(CLBLM_R_X63Y107_SLICE_X95Y107_A_XOR),
.I1(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I2(CLBLM_L_X64Y107_SLICE_X96Y107_AQ),
.I3(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I4(CLBLM_L_X62Y105_SLICE_X92Y105_BO5),
.I5(CLBLM_L_X64Y107_SLICE_X96Y107_CO6),
.O5(CLBLM_L_X64Y107_SLICE_X96Y107_AO5),
.O6(CLBLM_L_X64Y107_SLICE_X96Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y107_SLICE_X97Y107_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_R_X63Y100_SLICE_X94Y100_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X64Y107_SLICE_X97Y107_AO6),
.Q(CLBLM_L_X64Y107_SLICE_X97Y107_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y107_SLICE_X97Y107_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_R_X63Y100_SLICE_X94Y100_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X64Y107_SLICE_X97Y107_BO6),
.Q(CLBLM_L_X64Y107_SLICE_X97Y107_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0aca0a0a0aca0)
  ) CLBLM_L_X64Y107_SLICE_X97Y107_DLUT (
.I0(CLBLM_R_X49Y106_SLICE_X74Y106_AQ),
.I1(CLBLM_R_X63Y107_SLICE_X94Y107_D_XOR),
.I2(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I3(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I4(CLBLM_L_X62Y105_SLICE_X93Y105_AO6),
.I5(CLBLM_R_X63Y107_SLICE_X95Y107_C_XOR),
.O5(CLBLM_L_X64Y107_SLICE_X97Y107_DO5),
.O6(CLBLM_L_X64Y107_SLICE_X97Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cac0c0c0cac0)
  ) CLBLM_L_X64Y107_SLICE_X97Y107_CLUT (
.I0(CLBLM_R_X63Y107_SLICE_X94Y107_A_XOR),
.I1(CLBLM_L_X50Y104_SLICE_X76Y104_AQ),
.I2(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I3(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I4(CLBLM_L_X62Y105_SLICE_X93Y105_AO6),
.I5(CLBLM_R_X63Y106_SLICE_X95Y106_D_XOR),
.O5(CLBLM_L_X64Y107_SLICE_X97Y107_CO5),
.O6(CLBLM_L_X64Y107_SLICE_X97Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff05000404)
  ) CLBLM_L_X64Y107_SLICE_X97Y107_BLUT (
.I0(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I1(CLBLM_L_X64Y107_SLICE_X97Y107_BQ),
.I2(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I3(CLBLM_R_X63Y106_SLICE_X95Y106_D_XOR),
.I4(CLBLM_L_X62Y105_SLICE_X92Y105_BO5),
.I5(CLBLM_L_X64Y107_SLICE_X97Y107_CO6),
.O5(CLBLM_L_X64Y107_SLICE_X97Y107_BO5),
.O6(CLBLM_L_X64Y107_SLICE_X97Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff44ff00ff50)
  ) CLBLM_L_X64Y107_SLICE_X97Y107_ALUT (
.I0(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I1(CLBLM_R_X63Y107_SLICE_X95Y107_C_XOR),
.I2(CLBLM_L_X64Y107_SLICE_X97Y107_AQ),
.I3(CLBLM_L_X64Y107_SLICE_X97Y107_DO6),
.I4(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I5(CLBLM_L_X62Y105_SLICE_X92Y105_BO5),
.O5(CLBLM_L_X64Y107_SLICE_X97Y107_AO5),
.O6(CLBLM_L_X64Y107_SLICE_X97Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y108_SLICE_X96Y108_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_R_X63Y100_SLICE_X94Y100_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X64Y108_SLICE_X96Y108_AO6),
.Q(CLBLM_L_X64Y108_SLICE_X96Y108_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y108_SLICE_X96Y108_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_R_X63Y100_SLICE_X94Y100_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X64Y108_SLICE_X96Y108_BO6),
.Q(CLBLM_L_X64Y108_SLICE_X96Y108_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc5c5c5c0c0c5c0c0)
  ) CLBLM_L_X64Y108_SLICE_X96Y108_DLUT (
.I0(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I1(CLBLM_L_X50Y107_SLICE_X77Y107_AQ),
.I2(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I3(CLBLM_L_X62Y105_SLICE_X92Y105_BO5),
.I4(CLBLM_L_X64Y108_SLICE_X96Y108_BQ),
.I5(CLBLM_R_X63Y108_SLICE_X95Y108_C_XOR),
.O5(CLBLM_L_X64Y108_SLICE_X96Y108_DO5),
.O6(CLBLM_L_X64Y108_SLICE_X96Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcac0cac0cacac0c0)
  ) CLBLM_L_X64Y108_SLICE_X96Y108_CLUT (
.I0(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I1(CLBLM_L_X50Y106_SLICE_X76Y106_AQ),
.I2(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I3(CLBLM_R_X63Y107_SLICE_X95Y107_D_XOR),
.I4(CLBLM_R_X63Y108_SLICE_X94Y108_A_XOR),
.I5(CLBLM_L_X62Y105_SLICE_X93Y105_AO6),
.O5(CLBLM_L_X64Y108_SLICE_X96Y108_CO5),
.O6(CLBLM_L_X64Y108_SLICE_X96Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdcdcdcccccdccccc)
  ) CLBLM_L_X64Y108_SLICE_X96Y108_BLUT (
.I0(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I1(CLBLM_L_X64Y108_SLICE_X96Y108_DO6),
.I2(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I3(CLBLM_L_X62Y105_SLICE_X93Y105_AO6),
.I4(CLBLM_R_X63Y108_SLICE_X94Y108_D_XOR),
.I5(CLBLM_R_X63Y108_SLICE_X95Y108_C_XOR),
.O5(CLBLM_L_X64Y108_SLICE_X96Y108_BO5),
.O6(CLBLM_L_X64Y108_SLICE_X96Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00005410)
  ) CLBLM_L_X64Y108_SLICE_X96Y108_ALUT (
.I0(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I1(CLBLM_L_X62Y105_SLICE_X92Y105_BO5),
.I2(CLBLM_L_X64Y108_SLICE_X96Y108_AQ),
.I3(CLBLM_R_X63Y107_SLICE_X95Y107_D_XOR),
.I4(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I5(CLBLM_L_X64Y108_SLICE_X96Y108_CO6),
.O5(CLBLM_L_X64Y108_SLICE_X96Y108_AO5),
.O6(CLBLM_L_X64Y108_SLICE_X96Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y108_SLICE_X97Y108_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_R_X63Y100_SLICE_X94Y100_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X64Y108_SLICE_X97Y108_AO6),
.Q(CLBLM_L_X64Y108_SLICE_X97Y108_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y108_SLICE_X97Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y108_SLICE_X97Y108_DO5),
.O6(CLBLM_L_X64Y108_SLICE_X97Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y108_SLICE_X97Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y108_SLICE_X97Y108_CO5),
.O6(CLBLM_L_X64Y108_SLICE_X97Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50ba10ea40aa00)
  ) CLBLM_L_X64Y108_SLICE_X97Y108_BLUT (
.I0(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I1(CLBLM_L_X62Y105_SLICE_X93Y105_AO6),
.I2(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I3(CLBLM_L_X50Y106_SLICE_X76Y106_CQ),
.I4(CLBLM_R_X63Y108_SLICE_X95Y108_A_XOR),
.I5(CLBLM_R_X63Y108_SLICE_X94Y108_B_XOR),
.O5(CLBLM_L_X64Y108_SLICE_X97Y108_BO5),
.O6(CLBLM_L_X64Y108_SLICE_X97Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00ff44ff50)
  ) CLBLM_L_X64Y108_SLICE_X97Y108_ALUT (
.I0(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I1(CLBLM_R_X63Y108_SLICE_X95Y108_A_XOR),
.I2(CLBLM_L_X64Y108_SLICE_X97Y108_AQ),
.I3(CLBLM_L_X64Y108_SLICE_X97Y108_BO6),
.I4(CLBLM_L_X62Y105_SLICE_X92Y105_BO5),
.I5(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.O5(CLBLM_L_X64Y108_SLICE_X97Y108_AO5),
.O6(CLBLM_L_X64Y108_SLICE_X97Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y109_SLICE_X96Y109_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y100_SLICE_X92Y100_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X64Y109_SLICE_X96Y109_AO5),
.Q(CLBLM_L_X64Y109_SLICE_X96Y109_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X64Y109_SLICE_X96Y109_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y100_SLICE_X92Y100_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X64Y109_SLICE_X96Y109_AO6),
.Q(CLBLM_L_X64Y109_SLICE_X96Y109_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcffaa0c0c5500)
  ) CLBLM_L_X64Y109_SLICE_X96Y109_DLUT (
.I0(CLBLM_L_X62Y105_SLICE_X92Y105_BO5),
.I1(CLBLM_R_X63Y109_SLICE_X94Y109_D_XOR),
.I2(CLBLM_L_X62Y105_SLICE_X93Y105_AO6),
.I3(CLBLM_L_X64Y109_SLICE_X96Y109_A5Q),
.I4(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I5(CLBLM_R_X63Y109_SLICE_X95Y109_C_XOR),
.O5(CLBLM_L_X64Y109_SLICE_X96Y109_DO5),
.O6(CLBLM_L_X64Y109_SLICE_X96Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33cc00fa50fa50)
  ) CLBLM_L_X64Y109_SLICE_X96Y109_CLUT (
.I0(CLBLM_L_X62Y105_SLICE_X92Y105_BO5),
.I1(CLBLM_L_X62Y105_SLICE_X93Y105_AO6),
.I2(CLBLM_R_X63Y105_SLICE_X94Y105_AQ),
.I3(CLBLM_R_X63Y109_SLICE_X95Y109_B_XOR),
.I4(CLBLM_R_X63Y109_SLICE_X94Y109_C_XOR),
.I5(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.O5(CLBLM_L_X64Y109_SLICE_X96Y109_CO5),
.O6(CLBLM_L_X64Y109_SLICE_X96Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbbfcb8008830b8)
  ) CLBLM_L_X64Y109_SLICE_X96Y109_BLUT (
.I0(CLBLM_R_X63Y109_SLICE_X94Y109_A_XOR),
.I1(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I2(CLBLM_L_X64Y109_SLICE_X96Y109_AQ),
.I3(CLBLM_L_X62Y105_SLICE_X93Y105_AO6),
.I4(CLBLM_L_X62Y105_SLICE_X92Y105_BO5),
.I5(CLBLM_R_X63Y108_SLICE_X95Y108_D_XOR),
.O5(CLBLM_L_X64Y109_SLICE_X96Y109_BO5),
.O6(CLBLM_L_X64Y109_SLICE_X96Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff00ccccaaaa)
  ) CLBLM_L_X64Y109_SLICE_X96Y109_ALUT (
.I0(CLBLM_L_X64Y109_SLICE_X96Y109_DO6),
.I1(CLBLM_R_X49Y106_SLICE_X74Y106_AQ),
.I2(CLBLM_L_X50Y104_SLICE_X76Y104_AQ),
.I3(CLBLM_L_X64Y109_SLICE_X96Y109_BO6),
.I4(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I5(1'b1),
.O5(CLBLM_L_X64Y109_SLICE_X96Y109_AO5),
.O6(CLBLM_L_X64Y109_SLICE_X96Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y109_SLICE_X97Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y109_SLICE_X97Y109_DO5),
.O6(CLBLM_L_X64Y109_SLICE_X97Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y109_SLICE_X97Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y109_SLICE_X97Y109_CO5),
.O6(CLBLM_L_X64Y109_SLICE_X97Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y109_SLICE_X97Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y109_SLICE_X97Y109_BO5),
.O6(CLBLM_L_X64Y109_SLICE_X97Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X64Y109_SLICE_X97Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X64Y109_SLICE_X97Y109_AO5),
.O6(CLBLM_L_X64Y109_SLICE_X97Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y122_SLICE_X20Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y122_SLICE_X20Y122_DO5),
.O6(CLBLM_R_X15Y122_SLICE_X20Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y122_SLICE_X20Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y122_SLICE_X20Y122_CO5),
.O6(CLBLM_R_X15Y122_SLICE_X20Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y122_SLICE_X20Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y122_SLICE_X20Y122_BO5),
.O6(CLBLM_R_X15Y122_SLICE_X20Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555555)
  ) CLBLM_R_X15Y122_SLICE_X20Y122_ALUT (
.I0(LIOB33_X0Y123_IOB_X0Y123_I),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y122_SLICE_X20Y122_AO5),
.O6(CLBLM_R_X15Y122_SLICE_X20Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y122_SLICE_X21Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y122_SLICE_X21Y122_DO5),
.O6(CLBLM_R_X15Y122_SLICE_X21Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y122_SLICE_X21Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y122_SLICE_X21Y122_CO5),
.O6(CLBLM_R_X15Y122_SLICE_X21Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y122_SLICE_X21Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y122_SLICE_X21Y122_BO5),
.O6(CLBLM_R_X15Y122_SLICE_X21Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y122_SLICE_X21Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y122_SLICE_X21Y122_AO5),
.O6(CLBLM_R_X15Y122_SLICE_X21Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X47Y119_SLICE_X72Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X47Y119_SLICE_X72Y119_DO5),
.O6(CLBLM_R_X47Y119_SLICE_X72Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X47Y119_SLICE_X72Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X47Y119_SLICE_X72Y119_CO5),
.O6(CLBLM_R_X47Y119_SLICE_X72Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X47Y119_SLICE_X72Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X47Y119_SLICE_X72Y119_BO5),
.O6(CLBLM_R_X47Y119_SLICE_X72Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X47Y119_SLICE_X72Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X47Y119_SLICE_X72Y119_AO5),
.O6(CLBLM_R_X47Y119_SLICE_X72Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X47Y119_SLICE_X73Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(CLBLM_R_X15Y122_SLICE_X20Y122_AO6),
.D(CLBLM_L_X32Y119_SLICE_X46Y119_AQ),
.Q(CLBLM_R_X47Y119_SLICE_X73Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X47Y119_SLICE_X73Y119_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(CLBLM_R_X15Y122_SLICE_X20Y122_AO6),
.D(CLBLM_R_X47Y119_SLICE_X73Y119_AQ),
.Q(CLBLM_R_X47Y119_SLICE_X73Y119_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X47Y119_SLICE_X73Y119_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(CLBLM_R_X15Y122_SLICE_X20Y122_AO6),
.D(CLBLM_L_X32Y119_SLICE_X46Y119_BQ),
.Q(CLBLM_R_X47Y119_SLICE_X73Y119_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X47Y119_SLICE_X73Y119_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(CLBLM_R_X15Y122_SLICE_X20Y122_AO6),
.D(CLBLM_R_X47Y119_SLICE_X73Y119_CQ),
.Q(CLBLM_R_X47Y119_SLICE_X73Y119_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X47Y119_SLICE_X73Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X47Y119_SLICE_X73Y119_DO5),
.O6(CLBLM_R_X47Y119_SLICE_X73Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X47Y119_SLICE_X73Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X47Y119_SLICE_X73Y119_CO5),
.O6(CLBLM_R_X47Y119_SLICE_X73Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3000300030003000)
  ) CLBLM_R_X47Y119_SLICE_X73Y119_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X47Y119_SLICE_X73Y119_BQ),
.I2(CLBLM_R_X47Y119_SLICE_X73Y119_AQ),
.I3(CLBLM_L_X32Y119_SLICE_X46Y119_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X47Y119_SLICE_X73Y119_BO5),
.O6(CLBLM_R_X47Y119_SLICE_X73Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ffff00a00000)
  ) CLBLM_R_X47Y119_SLICE_X73Y119_ALUT (
.I0(CLBLM_R_X47Y119_SLICE_X73Y119_CQ),
.I1(1'b1),
.I2(LIOB33_X0Y119_IOB_X0Y120_I),
.I3(CLBLM_R_X47Y119_SLICE_X73Y119_DQ),
.I4(CLBLM_L_X32Y119_SLICE_X46Y119_BQ),
.I5(1'b1),
.O5(CLBLM_R_X47Y119_SLICE_X73Y119_AO5),
.O6(CLBLM_R_X47Y119_SLICE_X73Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X49Y104_SLICE_X74Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X49Y104_SLICE_X75Y104_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X49Y104_SLICE_X74Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X49Y104_SLICE_X74Y104_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X49Y104_SLICE_X75Y104_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(LIOB33_X0Y113_IOB_X0Y114_I),
.Q(CLBLM_R_X49Y104_SLICE_X74Y104_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y104_SLICE_X74Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y104_SLICE_X74Y104_DO5),
.O6(CLBLM_R_X49Y104_SLICE_X74Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y104_SLICE_X74Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y104_SLICE_X74Y104_CO5),
.O6(CLBLM_R_X49Y104_SLICE_X74Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y104_SLICE_X74Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y104_SLICE_X74Y104_BO5),
.O6(CLBLM_R_X49Y104_SLICE_X74Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y104_SLICE_X74Y104_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y104_SLICE_X74Y104_AO5),
.O6(CLBLM_R_X49Y104_SLICE_X74Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X49Y104_SLICE_X75Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X49Y104_SLICE_X75Y104_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(LIOB33_X0Y101_IOB_X0Y101_I),
.Q(CLBLM_R_X49Y104_SLICE_X75Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X49Y104_SLICE_X75Y104_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X49Y104_SLICE_X75Y104_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(LIOB33_X0Y101_IOB_X0Y102_I),
.Q(CLBLM_R_X49Y104_SLICE_X75Y104_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X49Y104_SLICE_X75Y104_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X49Y104_SLICE_X75Y104_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(LIOB33_X0Y103_IOB_X0Y103_I),
.Q(CLBLM_R_X49Y104_SLICE_X75Y104_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X49Y104_SLICE_X75Y104_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X49Y104_SLICE_X75Y104_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(LIOB33_X0Y103_IOB_X0Y104_I),
.Q(CLBLM_R_X49Y104_SLICE_X75Y104_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y104_SLICE_X75Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y104_SLICE_X75Y104_DO5),
.O6(CLBLM_R_X49Y104_SLICE_X75Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y104_SLICE_X75Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y104_SLICE_X75Y104_CO5),
.O6(CLBLM_R_X49Y104_SLICE_X75Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y104_SLICE_X75Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y104_SLICE_X75Y104_BO5),
.O6(CLBLM_R_X49Y104_SLICE_X75Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0303000303030003)
  ) CLBLM_R_X49Y104_SLICE_X75Y104_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I2(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I3(CLBLM_R_X49Y119_SLICE_X74Y119_BQ),
.I4(CLBLM_R_X49Y119_SLICE_X74Y119_AQ),
.I5(1'b1),
.O5(CLBLM_R_X49Y104_SLICE_X75Y104_AO5),
.O6(CLBLM_R_X49Y104_SLICE_X75Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y105_SLICE_X74Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y105_SLICE_X74Y105_DO5),
.O6(CLBLM_R_X49Y105_SLICE_X74Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y105_SLICE_X74Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y105_SLICE_X74Y105_CO5),
.O6(CLBLM_R_X49Y105_SLICE_X74Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y105_SLICE_X74Y105_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y105_SLICE_X74Y105_BO5),
.O6(CLBLM_R_X49Y105_SLICE_X74Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y105_SLICE_X74Y105_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y105_SLICE_X74Y105_AO5),
.O6(CLBLM_R_X49Y105_SLICE_X74Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X49Y105_SLICE_X75Y105_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X56Y98_SLICE_X84Y98_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y105_SLICE_X75Y105_CO6),
.Q(CLBLM_R_X49Y105_SLICE_X75Y105_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y105_SLICE_X75Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y105_SLICE_X75Y105_DO5),
.O6(CLBLM_R_X49Y105_SLICE_X75Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacacacacacacac)
  ) CLBLM_R_X49Y105_SLICE_X75Y105_CLUT (
.I0(CLBLM_R_X49Y105_SLICE_X75Y105_F7AMUX_O),
.I1(CLBLM_R_X49Y107_SLICE_X75Y107_F7AMUX_O),
.I2(CLBLM_R_X53Y100_SLICE_X81Y100_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y105_SLICE_X75Y105_CO5),
.O6(CLBLM_R_X49Y105_SLICE_X75Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7b7b7b4848487b48)
  ) CLBLM_R_X49Y105_SLICE_X75Y105_BLUT (
.I0(CLBLM_L_X56Y101_SLICE_X85Y101_CQ),
.I1(CLBLM_L_X50Y106_SLICE_X77Y106_AO5),
.I2(CLBLM_L_X56Y101_SLICE_X85Y101_AQ),
.I3(CLBLL_R_X57Y100_SLICE_X86Y100_CQ),
.I4(CLBLL_L_X54Y100_SLICE_X82Y100_BQ),
.I5(CLBLL_R_X57Y100_SLICE_X87Y100_CQ),
.O5(CLBLM_R_X49Y105_SLICE_X75Y105_BO5),
.O6(CLBLM_R_X49Y105_SLICE_X75Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h56565656569a569a)
  ) CLBLM_R_X49Y105_SLICE_X75Y105_ALUT (
.I0(CLBLM_L_X56Y101_SLICE_X85Y101_CQ),
.I1(CLBLM_L_X50Y106_SLICE_X77Y106_AO5),
.I2(CLBLM_L_X56Y101_SLICE_X85Y101_AQ),
.I3(CLBLL_R_X57Y100_SLICE_X86Y100_CQ),
.I4(1'b1),
.I5(CLBLL_R_X57Y100_SLICE_X86Y100_DQ),
.O5(CLBLM_R_X49Y105_SLICE_X75Y105_AO5),
.O6(CLBLM_R_X49Y105_SLICE_X75Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X49Y105_SLICE_X75Y105_MUXF7A (
.I0(CLBLM_R_X49Y105_SLICE_X75Y105_BO6),
.I1(CLBLM_R_X49Y105_SLICE_X75Y105_AO6),
.O(CLBLM_R_X49Y105_SLICE_X75Y105_F7AMUX_O),
.S(CLBLM_R_X49Y106_SLICE_X74Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X49Y106_SLICE_X74Y106_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X56Y98_SLICE_X84Y98_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y106_SLICE_X74Y106_AO6),
.Q(CLBLM_R_X49Y106_SLICE_X74Y106_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y106_SLICE_X74Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y106_SLICE_X74Y106_DO5),
.O6(CLBLM_R_X49Y106_SLICE_X74Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555000055550000)
  ) CLBLM_R_X49Y106_SLICE_X74Y106_CLUT (
.I0(CLBLL_L_X54Y100_SLICE_X82Y100_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X53Y101_SLICE_X81Y101_AQ),
.I5(1'b1),
.O5(CLBLM_R_X49Y106_SLICE_X74Y106_CO5),
.O6(CLBLM_R_X49Y106_SLICE_X74Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h503c503c53f353f3)
  ) CLBLM_R_X49Y106_SLICE_X74Y106_BLUT (
.I0(CLBLL_R_X57Y99_SLICE_X86Y99_BQ),
.I1(CLBLL_R_X57Y100_SLICE_X87Y100_CQ),
.I2(CLBLL_L_X54Y100_SLICE_X82Y100_BQ),
.I3(CLBLM_R_X53Y101_SLICE_X80Y101_BQ),
.I4(1'b1),
.I5(CLBLL_R_X57Y100_SLICE_X87Y100_AQ),
.O5(CLBLM_R_X49Y106_SLICE_X74Y106_BO5),
.O6(CLBLM_R_X49Y106_SLICE_X74Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f44770f0f4477)
  ) CLBLM_R_X49Y106_SLICE_X74Y106_ALUT (
.I0(CLBLM_R_X49Y107_SLICE_X75Y107_DO6),
.I1(CLBLM_R_X53Y101_SLICE_X81Y101_AQ),
.I2(CLBLM_R_X49Y106_SLICE_X75Y106_F7AMUX_O),
.I3(CLBLM_R_X49Y106_SLICE_X74Y106_BO6),
.I4(CLBLM_R_X53Y100_SLICE_X81Y100_AQ),
.I5(1'b1),
.O5(CLBLM_R_X49Y106_SLICE_X74Y106_AO5),
.O6(CLBLM_R_X49Y106_SLICE_X74Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X49Y106_SLICE_X75Y106_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X49Y104_SLICE_X75Y104_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(LIOB33_X0Y115_IOB_X0Y115_I),
.Q(CLBLM_R_X49Y106_SLICE_X75Y106_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X49Y106_SLICE_X75Y106_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X49Y104_SLICE_X75Y104_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(LIOB33_X0Y105_IOB_X0Y105_I),
.Q(CLBLM_R_X49Y106_SLICE_X75Y106_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X49Y106_SLICE_X75Y106_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X49Y104_SLICE_X75Y104_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_R_X49Y106_SLICE_X75Y106_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X49Y106_SLICE_X75Y106_DLUT (
.I0(CLBLL_R_X57Y100_SLICE_X87Y100_CQ),
.I1(CLBLM_L_X56Y101_SLICE_X85Y101_DQ),
.I2(CLBLL_R_X57Y101_SLICE_X87Y101_CQ),
.I3(CLBLL_R_X57Y100_SLICE_X86Y100_CQ),
.I4(CLBLM_L_X56Y101_SLICE_X85Y101_CQ),
.I5(CLBLL_R_X57Y100_SLICE_X86Y100_DQ),
.O5(CLBLM_R_X49Y106_SLICE_X75Y106_DO5),
.O6(CLBLM_R_X49Y106_SLICE_X75Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcf301dd103fc1dd1)
  ) CLBLM_R_X49Y106_SLICE_X75Y106_CLUT (
.I0(CLBLM_L_X50Y105_SLICE_X76Y105_BO6),
.I1(CLBLM_R_X49Y106_SLICE_X74Y106_CO6),
.I2(CLBLL_R_X57Y100_SLICE_X87Y100_BQ),
.I3(CLBLL_R_X57Y101_SLICE_X87Y101_DQ),
.I4(CLBLM_L_X50Y106_SLICE_X77Y106_AO5),
.I5(CLBLM_R_X49Y106_SLICE_X75Y106_DO6),
.O5(CLBLM_R_X49Y106_SLICE_X75Y106_CO5),
.O6(CLBLM_R_X49Y106_SLICE_X75Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88dd22778d8d2727)
  ) CLBLM_R_X49Y106_SLICE_X75Y106_BLUT (
.I0(CLBLM_L_X50Y106_SLICE_X77Y106_AO5),
.I1(CLBLL_R_X57Y100_SLICE_X87Y100_AQ),
.I2(CLBLM_L_X56Y101_SLICE_X85Y101_CQ),
.I3(CLBLL_R_X57Y101_SLICE_X87Y101_CQ),
.I4(CLBLL_R_X57Y100_SLICE_X87Y100_CQ),
.I5(CLBLL_L_X54Y100_SLICE_X82Y100_BQ),
.O5(CLBLM_R_X49Y106_SLICE_X75Y106_BO5),
.O6(CLBLM_R_X49Y106_SLICE_X75Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeeeee41111111b)
  ) CLBLM_R_X49Y106_SLICE_X75Y106_ALUT (
.I0(CLBLM_L_X50Y106_SLICE_X77Y106_AO5),
.I1(CLBLL_R_X57Y100_SLICE_X87Y100_AQ),
.I2(CLBLM_L_X56Y101_SLICE_X85Y101_CQ),
.I3(CLBLL_R_X57Y100_SLICE_X86Y100_DQ),
.I4(CLBLL_R_X57Y100_SLICE_X86Y100_CQ),
.I5(CLBLL_R_X57Y100_SLICE_X87Y100_CQ),
.O5(CLBLM_R_X49Y106_SLICE_X75Y106_AO5),
.O6(CLBLM_R_X49Y106_SLICE_X75Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X49Y106_SLICE_X75Y106_MUXF7A (
.I0(CLBLM_R_X49Y106_SLICE_X75Y106_BO6),
.I1(CLBLM_R_X49Y106_SLICE_X75Y106_AO6),
.O(CLBLM_R_X49Y106_SLICE_X75Y106_F7AMUX_O),
.S(CLBLM_R_X49Y106_SLICE_X74Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X49Y107_SLICE_X74Y107_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X62Y109_SLICE_X92Y109_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y107_SLICE_X74Y107_AO6),
.Q(CLBLM_R_X49Y107_SLICE_X74Y107_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4000000000000000)
  ) CLBLM_R_X49Y107_SLICE_X74Y107_DLUT (
.I0(CLBLM_L_X50Y105_SLICE_X76Y105_CO6),
.I1(CLBLM_R_X49Y108_SLICE_X75Y108_A_XOR),
.I2(CLBLM_R_X49Y108_SLICE_X75Y108_D_XOR),
.I3(CLBLM_R_X49Y109_SLICE_X75Y109_A_XOR),
.I4(CLBLM_R_X49Y108_SLICE_X75Y108_B_XOR),
.I5(CLBLM_R_X49Y108_SLICE_X75Y108_C_XOR),
.O5(CLBLM_R_X49Y107_SLICE_X74Y107_DO5),
.O6(CLBLM_R_X49Y107_SLICE_X74Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffffffffffffff)
  ) CLBLM_R_X49Y107_SLICE_X74Y107_CLUT (
.I0(CLBLL_R_X57Y97_SLICE_X86Y97_AQ),
.I1(CLBLM_R_X53Y101_SLICE_X80Y101_BQ),
.I2(CLBLM_R_X49Y108_SLICE_X75Y108_D_XOR),
.I3(CLBLM_R_X49Y108_SLICE_X75Y108_A_XOR),
.I4(CLBLM_R_X49Y108_SLICE_X75Y108_B_XOR),
.I5(CLBLM_R_X49Y108_SLICE_X75Y108_C_XOR),
.O5(CLBLM_R_X49Y107_SLICE_X74Y107_CO5),
.O6(CLBLM_R_X49Y107_SLICE_X74Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b8fc308b8bcf03)
  ) CLBLM_R_X49Y107_SLICE_X74Y107_BLUT (
.I0(CLBLM_L_X50Y109_SLICE_X77Y109_A_XOR),
.I1(CLBLL_L_X54Y100_SLICE_X82Y100_BQ),
.I2(CLBLM_R_X49Y109_SLICE_X75Y109_A_XOR),
.I3(CLBLM_L_X50Y109_SLICE_X76Y109_A_XOR),
.I4(CLBLM_R_X53Y101_SLICE_X80Y101_BQ),
.I5(CLBLM_R_X49Y107_SLICE_X74Y107_CO6),
.O5(CLBLM_R_X49Y107_SLICE_X74Y107_BO5),
.O6(CLBLM_R_X49Y107_SLICE_X74Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0b8f0b8f0b8f0b8)
  ) CLBLM_R_X49Y107_SLICE_X74Y107_ALUT (
.I0(CLBLM_R_X49Y108_SLICE_X74Y108_A5Q),
.I1(CLBLL_R_X57Y102_SLICE_X86Y102_AQ),
.I2(CLBLM_L_X50Y105_SLICE_X77Y105_AQ),
.I3(CLBLL_R_X57Y102_SLICE_X86Y102_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y107_SLICE_X74Y107_AO5),
.O6(CLBLM_R_X49Y107_SLICE_X74Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X49Y107_SLICE_X75Y107_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X49Y104_SLICE_X75Y104_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(LIOB33_X0Y113_IOB_X0Y113_I),
.Q(CLBLM_R_X49Y107_SLICE_X75Y107_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X49Y107_SLICE_X75Y107_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X49Y104_SLICE_X75Y104_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(LIOB33_X0Y107_IOB_X0Y107_I),
.Q(CLBLM_R_X49Y107_SLICE_X75Y107_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X49Y107_SLICE_X75Y107_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X49Y104_SLICE_X75Y104_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(LIOB33_X0Y109_IOB_X0Y109_I),
.Q(CLBLM_R_X49Y107_SLICE_X75Y107_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h043737048cbfbf8c)
  ) CLBLM_R_X49Y107_SLICE_X75Y107_DLUT (
.I0(CLBLM_R_X53Y101_SLICE_X80Y101_BQ),
.I1(CLBLL_L_X54Y100_SLICE_X82Y100_BQ),
.I2(CLBLM_L_X50Y108_SLICE_X76Y108_D_XOR),
.I3(CLBLM_R_X49Y107_SLICE_X75Y107_CO5),
.I4(CLBLM_R_X49Y108_SLICE_X75Y108_D_XOR),
.I5(CLBLM_L_X50Y108_SLICE_X77Y108_D_XOR),
.O5(CLBLM_R_X49Y107_SLICE_X75Y107_DO5),
.O6(CLBLM_R_X49Y107_SLICE_X75Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5fffffff7fffffff)
  ) CLBLM_R_X49Y107_SLICE_X75Y107_CLUT (
.I0(CLBLM_R_X53Y101_SLICE_X80Y101_BQ),
.I1(CLBLM_R_X49Y108_SLICE_X75Y108_C_XOR),
.I2(CLBLL_R_X57Y97_SLICE_X86Y97_AQ),
.I3(CLBLM_R_X49Y108_SLICE_X75Y108_A_XOR),
.I4(CLBLM_R_X49Y108_SLICE_X75Y108_B_XOR),
.I5(1'b1),
.O5(CLBLM_R_X49Y107_SLICE_X75Y107_CO5),
.O6(CLBLM_R_X49Y107_SLICE_X75Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddaa55dd885500)
  ) CLBLM_R_X49Y107_SLICE_X75Y107_BLUT (
.I0(CLBLL_L_X54Y100_SLICE_X82Y100_BQ),
.I1(CLBLL_R_X57Y101_SLICE_X87Y101_DQ),
.I2(1'b1),
.I3(CLBLM_L_X56Y101_SLICE_X85Y101_AQ),
.I4(CLBLM_R_X53Y101_SLICE_X80Y101_BQ),
.I5(CLBLM_L_X56Y101_SLICE_X85Y101_CQ),
.O5(CLBLM_R_X49Y107_SLICE_X75Y107_BO5),
.O6(CLBLM_R_X49Y107_SLICE_X75Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee4ee444bb1bb111)
  ) CLBLM_R_X49Y107_SLICE_X75Y107_ALUT (
.I0(CLBLL_L_X54Y100_SLICE_X82Y100_BQ),
.I1(CLBLM_R_X49Y108_SLICE_X75Y108_C_XOR),
.I2(CLBLM_R_X53Y101_SLICE_X80Y101_BQ),
.I3(CLBLM_L_X50Y108_SLICE_X77Y108_C_XOR),
.I4(CLBLM_L_X50Y108_SLICE_X76Y108_C_XOR),
.I5(CLBLM_R_X49Y107_SLICE_X75Y107_CO6),
.O5(CLBLM_R_X49Y107_SLICE_X75Y107_AO5),
.O6(CLBLM_R_X49Y107_SLICE_X75Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X49Y107_SLICE_X75Y107_MUXF7A (
.I0(CLBLM_R_X49Y107_SLICE_X75Y107_BO6),
.I1(CLBLM_R_X49Y107_SLICE_X75Y107_AO6),
.O(CLBLM_R_X49Y107_SLICE_X75Y107_F7AMUX_O),
.S(CLBLM_R_X53Y101_SLICE_X81Y101_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X49Y108_SLICE_X74Y108_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X49Y110_SLICE_X74Y110_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y108_SLICE_X74Y108_AO5),
.Q(CLBLM_R_X49Y108_SLICE_X74Y108_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X49Y108_SLICE_X74Y108_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X49Y110_SLICE_X74Y110_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y108_SLICE_X74Y108_BO5),
.Q(CLBLM_R_X49Y108_SLICE_X74Y108_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X49Y108_SLICE_X74Y108_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X49Y110_SLICE_X74Y110_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y108_SLICE_X74Y108_CO5),
.Q(CLBLM_R_X49Y108_SLICE_X74Y108_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X49Y108_SLICE_X74Y108_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X49Y110_SLICE_X74Y110_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y108_SLICE_X74Y108_AO6),
.Q(CLBLM_R_X49Y108_SLICE_X74Y108_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X49Y108_SLICE_X74Y108_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X49Y110_SLICE_X74Y110_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y108_SLICE_X74Y108_BO6),
.Q(CLBLM_R_X49Y108_SLICE_X74Y108_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X49Y108_SLICE_X74Y108_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X49Y110_SLICE_X74Y110_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y108_SLICE_X74Y108_CO6),
.Q(CLBLM_R_X49Y108_SLICE_X74Y108_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8b8bb8b8cf03fc30)
  ) CLBLM_R_X49Y108_SLICE_X74Y108_DLUT (
.I0(CLBLM_L_X50Y109_SLICE_X77Y109_B_XOR),
.I1(CLBLL_L_X54Y100_SLICE_X82Y100_BQ),
.I2(CLBLM_R_X49Y107_SLICE_X74Y107_DO6),
.I3(CLBLM_L_X50Y109_SLICE_X76Y109_B_XOR),
.I4(CLBLM_R_X49Y109_SLICE_X75Y109_B_XOR),
.I5(CLBLM_R_X53Y101_SLICE_X80Y101_BQ),
.O5(CLBLM_R_X49Y108_SLICE_X74Y108_DO5),
.O6(CLBLM_R_X49Y108_SLICE_X74Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc3300e2e2e2e2)
  ) CLBLM_R_X49Y108_SLICE_X74Y108_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLM_L_X62Y105_SLICE_X92Y105_CQ),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(1'b1),
.O5(CLBLM_R_X49Y108_SLICE_X74Y108_CO5),
.O6(CLBLM_R_X49Y108_SLICE_X74Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacacacfff00f00)
  ) CLBLM_R_X49Y108_SLICE_X74Y108_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(CLBLM_L_X62Y105_SLICE_X92Y105_CQ),
.I3(LIOB33_X0Y113_IOB_X0Y113_I),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X49Y108_SLICE_X74Y108_BO5),
.O6(CLBLM_R_X49Y108_SLICE_X74Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00f0aaf0aa)
  ) CLBLM_R_X49Y108_SLICE_X74Y108_ALUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(CLBLM_L_X62Y105_SLICE_X92Y105_CQ),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(1'b1),
.O5(CLBLM_R_X49Y108_SLICE_X74Y108_AO5),
.O6(CLBLM_R_X49Y108_SLICE_X74Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X49Y108_SLICE_X75Y108_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X49Y104_SLICE_X75Y104_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y108_SLICE_X75Y108_AO5),
.Q(CLBLM_R_X49Y108_SLICE_X75Y108_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X49Y108_SLICE_X75Y108_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X49Y104_SLICE_X75Y104_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y108_SLICE_X75Y108_BO5),
.Q(CLBLM_R_X49Y108_SLICE_X75Y108_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X49Y108_SLICE_X75Y108_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X49Y104_SLICE_X75Y104_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y108_SLICE_X75Y108_CO5),
.Q(CLBLM_R_X49Y108_SLICE_X75Y108_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X49Y108_SLICE_X75Y108_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X49Y104_SLICE_X75Y104_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y108_SLICE_X75Y108_DO5),
.Q(CLBLM_R_X49Y108_SLICE_X75Y108_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X49Y108_SLICE_X75Y108_CARRY4 (
.CI(1'b0),
.CO({CLBLM_R_X49Y108_SLICE_X75Y108_D_CY, CLBLM_R_X49Y108_SLICE_X75Y108_C_CY, CLBLM_R_X49Y108_SLICE_X75Y108_B_CY, CLBLM_R_X49Y108_SLICE_X75Y108_A_CY}),
.CYINIT(1'b0),
.DI({CLBLL_R_X57Y100_SLICE_X87Y100_AQ, CLBLM_L_X56Y101_SLICE_X85Y101_AQ, CLBLL_R_X57Y100_SLICE_X86Y100_BQ, CLBLL_R_X57Y100_SLICE_X86Y100_AQ}),
.O({CLBLM_R_X49Y108_SLICE_X75Y108_D_XOR, CLBLM_R_X49Y108_SLICE_X75Y108_C_XOR, CLBLM_R_X49Y108_SLICE_X75Y108_B_XOR, CLBLM_R_X49Y108_SLICE_X75Y108_A_XOR}),
.S({CLBLM_R_X49Y108_SLICE_X75Y108_DO6, CLBLM_R_X49Y108_SLICE_X75Y108_CO6, CLBLM_R_X49Y108_SLICE_X75Y108_BO6, CLBLM_R_X49Y108_SLICE_X75Y108_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0ff0f0aaaaaaaa)
  ) CLBLM_R_X49Y108_SLICE_X75Y108_DLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(1'b1),
.I2(CLBLL_R_X57Y100_SLICE_X87Y100_CQ),
.I3(1'b1),
.I4(CLBLL_R_X57Y100_SLICE_X87Y100_AQ),
.I5(1'b1),
.O5(CLBLM_R_X49Y108_SLICE_X75Y108_DO5),
.O6(CLBLM_R_X49Y108_SLICE_X75Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ccccaaaaaaaa)
  ) CLBLM_R_X49Y108_SLICE_X75Y108_CLUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(CLBLM_L_X56Y101_SLICE_X85Y101_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X56Y101_SLICE_X85Y101_AQ),
.I5(1'b1),
.O5(CLBLM_R_X49Y108_SLICE_X75Y108_CO5),
.O6(CLBLM_R_X49Y108_SLICE_X75Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3cff00ff00)
  ) CLBLM_R_X49Y108_SLICE_X75Y108_BLUT (
.I0(1'b1),
.I1(CLBLL_R_X57Y100_SLICE_X86Y100_BQ),
.I2(CLBLL_R_X57Y100_SLICE_X86Y100_CQ),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y108_SLICE_X75Y108_BO5),
.O6(CLBLM_R_X49Y108_SLICE_X75Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3caaaaaaaa)
  ) CLBLM_R_X49Y108_SLICE_X75Y108_ALUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(CLBLL_R_X57Y100_SLICE_X86Y100_DQ),
.I2(CLBLL_R_X57Y100_SLICE_X86Y100_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y108_SLICE_X75Y108_AO5),
.O6(CLBLM_R_X49Y108_SLICE_X75Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X49Y109_SLICE_X74Y109_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X62Y109_SLICE_X92Y109_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y109_SLICE_X74Y109_AO6),
.Q(CLBLM_R_X49Y109_SLICE_X74Y109_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X49Y109_SLICE_X74Y109_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X62Y109_SLICE_X92Y109_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y109_SLICE_X74Y109_BO6),
.Q(CLBLM_R_X49Y109_SLICE_X74Y109_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X49Y109_SLICE_X74Y109_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X62Y109_SLICE_X92Y109_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y109_SLICE_X74Y109_CO6),
.Q(CLBLM_R_X49Y109_SLICE_X74Y109_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X49Y109_SLICE_X74Y109_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X62Y109_SLICE_X92Y109_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y109_SLICE_X74Y109_DO6),
.Q(CLBLM_R_X49Y109_SLICE_X74Y109_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaafafa0a0a)
  ) CLBLM_R_X49Y109_SLICE_X74Y109_DLUT (
.I0(CLBLM_L_X50Y104_SLICE_X76Y104_AQ),
.I1(1'b1),
.I2(CLBLL_R_X57Y102_SLICE_X86Y102_AQ),
.I3(1'b1),
.I4(CLBLM_R_X49Y108_SLICE_X74Y108_AQ),
.I5(CLBLL_R_X57Y102_SLICE_X86Y102_BQ),
.O5(CLBLM_R_X49Y109_SLICE_X74Y109_DO5),
.O6(CLBLM_R_X49Y109_SLICE_X74Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0f0f0aaf0f0)
  ) CLBLM_R_X49Y109_SLICE_X74Y109_CLUT (
.I0(CLBLM_R_X49Y108_SLICE_X74Y108_C5Q),
.I1(1'b1),
.I2(CLBLM_L_X50Y107_SLICE_X77Y107_AQ),
.I3(CLBLL_R_X57Y102_SLICE_X86Y102_BQ),
.I4(CLBLL_R_X57Y102_SLICE_X86Y102_AQ),
.I5(1'b1),
.O5(CLBLM_R_X49Y109_SLICE_X74Y109_CO5),
.O6(CLBLM_R_X49Y109_SLICE_X74Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0faf0faf050f050)
  ) CLBLM_R_X49Y109_SLICE_X74Y109_BLUT (
.I0(CLBLL_R_X57Y102_SLICE_X86Y102_AQ),
.I1(1'b1),
.I2(CLBLM_L_X50Y106_SLICE_X76Y106_CQ),
.I3(CLBLL_R_X57Y102_SLICE_X86Y102_BQ),
.I4(1'b1),
.I5(CLBLM_R_X49Y108_SLICE_X74Y108_B5Q),
.O5(CLBLM_R_X49Y109_SLICE_X74Y109_BO5),
.O6(CLBLM_R_X49Y109_SLICE_X74Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffdd0088ffdd0088)
  ) CLBLM_R_X49Y109_SLICE_X74Y109_ALUT (
.I0(CLBLL_R_X57Y102_SLICE_X86Y102_AQ),
.I1(CLBLM_R_X49Y108_SLICE_X74Y108_BQ),
.I2(1'b1),
.I3(CLBLL_R_X57Y102_SLICE_X86Y102_BQ),
.I4(CLBLM_L_X50Y106_SLICE_X76Y106_AQ),
.I5(1'b1),
.O5(CLBLM_R_X49Y109_SLICE_X74Y109_AO5),
.O6(CLBLM_R_X49Y109_SLICE_X74Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X49Y109_SLICE_X75Y109_CARRY4 (
.CI(CLBLM_R_X49Y108_SLICE_X75Y108_COUT),
.CO({CLBLM_R_X49Y109_SLICE_X75Y109_D_CY, CLBLM_R_X49Y109_SLICE_X75Y109_C_CY, CLBLM_R_X49Y109_SLICE_X75Y109_B_CY, CLBLM_R_X49Y109_SLICE_X75Y109_A_CY}),
.CYINIT(1'b0),
.DI({CLBLL_R_X57Y99_SLICE_X86Y99_AQ, CLBLL_R_X57Y100_SLICE_X87Y100_BQ, CLBLM_L_X56Y101_SLICE_X85Y101_BQ, CLBLL_R_X57Y101_SLICE_X87Y101_AQ}),
.O({CLBLM_R_X49Y109_SLICE_X75Y109_D_XOR, CLBLM_R_X49Y109_SLICE_X75Y109_C_XOR, CLBLM_R_X49Y109_SLICE_X75Y109_B_XOR, CLBLM_R_X49Y109_SLICE_X75Y109_A_XOR}),
.S({CLBLM_R_X49Y109_SLICE_X75Y109_DO6, CLBLM_R_X49Y109_SLICE_X75Y109_CO6, CLBLM_R_X49Y109_SLICE_X75Y109_BO6, CLBLM_R_X49Y109_SLICE_X75Y109_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555aaaa5555aaaa)
  ) CLBLM_R_X49Y109_SLICE_X75Y109_DLUT (
.I0(CLBLL_R_X57Y99_SLICE_X86Y99_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_R_X57Y99_SLICE_X86Y99_AQ),
.I5(1'b1),
.O5(CLBLM_R_X49Y109_SLICE_X75Y109_DO5),
.O6(CLBLM_R_X49Y109_SLICE_X75Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cc33cc33cc33cc)
  ) CLBLM_R_X49Y109_SLICE_X75Y109_CLUT (
.I0(1'b1),
.I1(CLBLL_R_X57Y100_SLICE_X87Y100_BQ),
.I2(1'b1),
.I3(CLBLL_R_X57Y101_SLICE_X87Y101_DQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y109_SLICE_X75Y109_CO5),
.O6(CLBLM_R_X49Y109_SLICE_X75Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffff0000ffff00)
  ) CLBLM_R_X49Y109_SLICE_X75Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X56Y101_SLICE_X85Y101_DQ),
.I4(CLBLM_L_X56Y101_SLICE_X85Y101_BQ),
.I5(1'b1),
.O5(CLBLM_R_X49Y109_SLICE_X75Y109_BO5),
.O6(CLBLM_R_X49Y109_SLICE_X75Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0ff0f00f0ff0f0)
  ) CLBLM_R_X49Y109_SLICE_X75Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_R_X57Y101_SLICE_X87Y101_CQ),
.I3(1'b1),
.I4(CLBLL_R_X57Y101_SLICE_X87Y101_AQ),
.I5(1'b1),
.O5(CLBLM_R_X49Y109_SLICE_X75Y109_AO5),
.O6(CLBLM_R_X49Y109_SLICE_X75Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X49Y110_SLICE_X74Y110_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X49Y110_SLICE_X74Y110_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y110_SLICE_X74Y110_AO5),
.Q(CLBLM_R_X49Y110_SLICE_X74Y110_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X49Y110_SLICE_X74Y110_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X49Y110_SLICE_X74Y110_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y110_SLICE_X74Y110_AO6),
.Q(CLBLM_R_X49Y110_SLICE_X74Y110_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y110_SLICE_X74Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y110_SLICE_X74Y110_DO5),
.O6(CLBLM_R_X49Y110_SLICE_X74Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y110_SLICE_X74Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y110_SLICE_X74Y110_CO5),
.O6(CLBLM_R_X49Y110_SLICE_X74Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000f0ff0000)
  ) CLBLM_R_X49Y110_SLICE_X74Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X49Y119_SLICE_X74Y119_AQ),
.I3(CLBLM_R_X49Y119_SLICE_X74Y119_BQ),
.I4(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I5(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.O5(CLBLM_R_X49Y110_SLICE_X74Y110_BO5),
.O6(CLBLM_R_X49Y110_SLICE_X74Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ccccf0f0aaaa)
  ) CLBLM_R_X49Y110_SLICE_X74Y110_ALUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(CLBLM_L_X62Y105_SLICE_X92Y105_CQ),
.I5(1'b1),
.O5(CLBLM_R_X49Y110_SLICE_X74Y110_AO5),
.O6(CLBLM_R_X49Y110_SLICE_X74Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X49Y110_SLICE_X75Y110_CARRY4 (
.CI(CLBLM_R_X49Y109_SLICE_X75Y109_COUT),
.CO({CLBLM_R_X49Y110_SLICE_X75Y110_D_CY, CLBLM_R_X49Y110_SLICE_X75Y110_C_CY, CLBLM_R_X49Y110_SLICE_X75Y110_B_CY, CLBLM_R_X49Y110_SLICE_X75Y110_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X49Y110_SLICE_X75Y110_D_XOR, CLBLM_R_X49Y110_SLICE_X75Y110_C_XOR, CLBLM_R_X49Y110_SLICE_X75Y110_B_XOR, CLBLM_R_X49Y110_SLICE_X75Y110_A_XOR}),
.S({CLBLM_R_X49Y110_SLICE_X75Y110_DO6, CLBLM_R_X49Y110_SLICE_X75Y110_CO6, CLBLM_R_X49Y110_SLICE_X75Y110_BO6, CLBLM_R_X49Y110_SLICE_X75Y110_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y110_SLICE_X75Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y110_SLICE_X75Y110_DO5),
.O6(CLBLM_R_X49Y110_SLICE_X75Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y110_SLICE_X75Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y110_SLICE_X75Y110_CO5),
.O6(CLBLM_R_X49Y110_SLICE_X75Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y110_SLICE_X75Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y110_SLICE_X75Y110_BO5),
.O6(CLBLM_R_X49Y110_SLICE_X75Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffff)
  ) CLBLM_R_X49Y110_SLICE_X75Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y110_SLICE_X75Y110_AO5),
.O6(CLBLM_R_X49Y110_SLICE_X75Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X49Y111_SLICE_X74Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X62Y109_SLICE_X92Y109_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y111_SLICE_X74Y111_AO6),
.Q(CLBLM_R_X49Y111_SLICE_X74Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X49Y111_SLICE_X74Y111_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X62Y109_SLICE_X92Y109_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y111_SLICE_X74Y111_BO6),
.Q(CLBLM_R_X49Y111_SLICE_X74Y111_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X49Y111_SLICE_X74Y111_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X62Y109_SLICE_X92Y109_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y111_SLICE_X74Y111_CO6),
.Q(CLBLM_R_X49Y111_SLICE_X74Y111_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y111_SLICE_X74Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y111_SLICE_X74Y111_DO5),
.O6(CLBLM_R_X49Y111_SLICE_X74Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haacaaacaaacaaaca)
  ) CLBLM_R_X49Y111_SLICE_X74Y111_CLUT (
.I0(CLBLM_L_X50Y107_SLICE_X76Y107_BQ),
.I1(CLBLM_R_X49Y108_SLICE_X74Y108_CQ),
.I2(CLBLL_R_X57Y102_SLICE_X86Y102_AQ),
.I3(CLBLL_R_X57Y102_SLICE_X86Y102_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y111_SLICE_X74Y111_CO5),
.O6(CLBLM_R_X49Y111_SLICE_X74Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccf0cccccccc)
  ) CLBLM_R_X49Y111_SLICE_X74Y111_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X49Y106_SLICE_X74Y106_AQ),
.I2(CLBLM_R_X49Y110_SLICE_X74Y110_A5Q),
.I3(CLBLL_R_X57Y102_SLICE_X86Y102_BQ),
.I4(1'b1),
.I5(CLBLL_R_X57Y102_SLICE_X86Y102_AQ),
.O5(CLBLM_R_X49Y111_SLICE_X74Y111_BO5),
.O6(CLBLM_R_X49Y111_SLICE_X74Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff3300cc0000)
  ) CLBLM_R_X49Y111_SLICE_X74Y111_ALUT (
.I0(1'b1),
.I1(CLBLL_R_X57Y102_SLICE_X86Y102_AQ),
.I2(1'b1),
.I3(CLBLL_R_X57Y102_SLICE_X86Y102_BQ),
.I4(CLBLM_R_X49Y110_SLICE_X74Y110_AQ),
.I5(CLBLM_R_X49Y105_SLICE_X75Y105_CQ),
.O5(CLBLM_R_X49Y111_SLICE_X74Y111_AO5),
.O6(CLBLM_R_X49Y111_SLICE_X74Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X49Y111_SLICE_X75Y111_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X49Y111_SLICE_X75Y111_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y111_SLICE_X75Y111_AO5),
.Q(CLBLM_R_X49Y111_SLICE_X75Y111_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X49Y111_SLICE_X75Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X49Y111_SLICE_X75Y111_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y111_SLICE_X75Y111_AO6),
.Q(CLBLM_R_X49Y111_SLICE_X75Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y111_SLICE_X75Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y111_SLICE_X75Y111_DO5),
.O6(CLBLM_R_X49Y111_SLICE_X75Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y111_SLICE_X75Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y111_SLICE_X75Y111_CO5),
.O6(CLBLM_R_X49Y111_SLICE_X75Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3333ffff3333)
  ) CLBLM_R_X49Y111_SLICE_X75Y111_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X49Y119_SLICE_X74Y119_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X49Y119_SLICE_X74Y119_AQ),
.I5(1'b1),
.O5(CLBLM_R_X49Y111_SLICE_X75Y111_BO5),
.O6(CLBLM_R_X49Y111_SLICE_X75Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff330000ffcc0000)
  ) CLBLM_R_X49Y111_SLICE_X75Y111_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X62Y105_SLICE_X92Y105_CQ),
.I2(1'b1),
.I3(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I4(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I5(1'b1),
.O5(CLBLM_R_X49Y111_SLICE_X75Y111_AO5),
.O6(CLBLM_R_X49Y111_SLICE_X75Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X49Y119_SLICE_X74Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y119_SLICE_X74Y119_AO6),
.Q(CLBLM_R_X49Y119_SLICE_X74Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X49Y119_SLICE_X74Y119_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y119_SLICE_X74Y119_BO6),
.Q(CLBLM_R_X49Y119_SLICE_X74Y119_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y119_SLICE_X74Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y119_SLICE_X74Y119_DO5),
.O6(CLBLM_R_X49Y119_SLICE_X74Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y119_SLICE_X74Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y119_SLICE_X74Y119_CO5),
.O6(CLBLM_R_X49Y119_SLICE_X74Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h010f010f010f000c)
  ) CLBLM_R_X49Y119_SLICE_X74Y119_BLUT (
.I0(LIOB33_X0Y121_IOB_X0Y121_I),
.I1(CLBLM_R_X49Y119_SLICE_X74Y119_BQ),
.I2(CLBLM_R_X49Y119_SLICE_X74Y119_AQ),
.I3(CLBLM_R_X47Y119_SLICE_X73Y119_BO6),
.I4(CLBLM_L_X56Y102_SLICE_X85Y102_A5Q),
.I5(CLBLM_R_X47Y119_SLICE_X73Y119_AO5),
.O5(CLBLM_R_X49Y119_SLICE_X74Y119_BO5),
.O6(CLBLM_R_X49Y119_SLICE_X74Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0e000f0f0e000e0c)
  ) CLBLM_R_X49Y119_SLICE_X74Y119_ALUT (
.I0(LIOB33_X0Y121_IOB_X0Y121_I),
.I1(CLBLM_R_X49Y119_SLICE_X74Y119_BQ),
.I2(CLBLM_R_X49Y119_SLICE_X74Y119_AQ),
.I3(CLBLM_R_X47Y119_SLICE_X73Y119_BO6),
.I4(CLBLM_R_X47Y119_SLICE_X73Y119_AO6),
.I5(LIOB33_X0Y119_IOB_X0Y120_I),
.O5(CLBLM_R_X49Y119_SLICE_X74Y119_AO5),
.O6(CLBLM_R_X49Y119_SLICE_X74Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y119_SLICE_X75Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y119_SLICE_X75Y119_DO5),
.O6(CLBLM_R_X49Y119_SLICE_X75Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y119_SLICE_X75Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y119_SLICE_X75Y119_CO5),
.O6(CLBLM_R_X49Y119_SLICE_X75Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y119_SLICE_X75Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y119_SLICE_X75Y119_BO5),
.O6(CLBLM_R_X49Y119_SLICE_X75Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y119_SLICE_X75Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y119_SLICE_X75Y119_AO5),
.O6(CLBLM_R_X49Y119_SLICE_X75Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X53Y98_SLICE_X80Y98_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X53Y98_SLICE_X80Y98_DO5),
.O6(CLBLM_R_X53Y98_SLICE_X80Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X53Y98_SLICE_X80Y98_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X53Y98_SLICE_X80Y98_CO5),
.O6(CLBLM_R_X53Y98_SLICE_X80Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X53Y98_SLICE_X80Y98_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X53Y98_SLICE_X80Y98_BO5),
.O6(CLBLM_R_X53Y98_SLICE_X80Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X53Y98_SLICE_X80Y98_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X53Y98_SLICE_X80Y98_AO5),
.O6(CLBLM_R_X53Y98_SLICE_X80Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X53Y98_SLICE_X81Y98_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X53Y98_SLICE_X81Y98_DO5),
.O6(CLBLM_R_X53Y98_SLICE_X81Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2226000122220000)
  ) CLBLM_R_X53Y98_SLICE_X81Y98_CLUT (
.I0(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I1(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.I2(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.I3(CLBLM_R_X53Y100_SLICE_X81Y100_AO5),
.I4(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.I5(CLBLM_R_X49Y107_SLICE_X75Y107_DQ),
.O5(CLBLM_R_X53Y98_SLICE_X81Y98_CO5),
.O6(CLBLM_R_X53Y98_SLICE_X81Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000221100000aee)
  ) CLBLM_R_X53Y98_SLICE_X81Y98_BLUT (
.I0(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.I1(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.I2(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.I3(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I4(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I5(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.O5(CLBLM_R_X53Y98_SLICE_X81Y98_BO5),
.O6(CLBLM_R_X53Y98_SLICE_X81Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffaaffba)
  ) CLBLM_R_X53Y98_SLICE_X81Y98_ALUT (
.I0(CLBLL_L_X52Y99_SLICE_X78Y99_AO6),
.I1(CLBLM_R_X53Y99_SLICE_X80Y99_AO5),
.I2(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.I3(CLBLM_R_X53Y98_SLICE_X81Y98_BO6),
.I4(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I5(CLBLM_R_X53Y98_SLICE_X81Y98_CO6),
.O5(CLBLM_R_X53Y98_SLICE_X81Y98_AO5),
.O6(CLBLM_R_X53Y98_SLICE_X81Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000c00000800)
  ) CLBLM_R_X53Y99_SLICE_X80Y99_DLUT (
.I0(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.I1(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I2(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I3(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.I4(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.I5(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.O5(CLBLM_R_X53Y99_SLICE_X80Y99_DO5),
.O6(CLBLM_R_X53Y99_SLICE_X80Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f4f0f0f0f8f0f8)
  ) CLBLM_R_X53Y99_SLICE_X80Y99_CLUT (
.I0(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I1(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.I2(CLBLM_R_X53Y100_SLICE_X81Y100_DO6),
.I3(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.I4(CLBLM_L_X56Y97_SLICE_X84Y97_AO6),
.I5(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.O5(CLBLM_R_X53Y99_SLICE_X80Y99_CO5),
.O6(CLBLM_R_X53Y99_SLICE_X80Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffb00500000)
  ) CLBLM_R_X53Y99_SLICE_X80Y99_BLUT (
.I0(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.I1(CLBLM_R_X49Y108_SLICE_X75Y108_DQ),
.I2(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.I3(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.I4(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I5(1'b1),
.O5(CLBLM_R_X53Y99_SLICE_X80Y99_BO5),
.O6(CLBLM_R_X53Y99_SLICE_X80Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffaffffffafff)
  ) CLBLM_R_X53Y99_SLICE_X80Y99_ALUT (
.I0(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.I1(1'b1),
.I2(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.I3(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.I4(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I5(1'b1),
.O5(CLBLM_R_X53Y99_SLICE_X80Y99_AO5),
.O6(CLBLM_R_X53Y99_SLICE_X80Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X53Y99_SLICE_X81Y99_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X0Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X53Y99_SLICE_X81Y99_BQ),
.Q(CLBLM_R_X53Y99_SLICE_X81Y99_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X53Y99_SLICE_X81Y99_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X0Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X53Y99_SLICE_X81Y99_BO6),
.Q(CLBLM_R_X53Y99_SLICE_X81Y99_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000100)
  ) CLBLM_R_X53Y99_SLICE_X81Y99_DLUT (
.I0(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I1(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.I2(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.I3(CLBLL_L_X54Y99_SLICE_X83Y99_BO5),
.I4(CLBLM_R_X49Y108_SLICE_X75Y108_DQ),
.I5(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.O5(CLBLM_R_X53Y99_SLICE_X81Y99_DO5),
.O6(CLBLM_R_X53Y99_SLICE_X81Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X53Y99_SLICE_X81Y99_CLUT (
.I0(CLBLM_R_X53Y99_SLICE_X81Y99_AO6),
.I1(CLBLL_L_X52Y99_SLICE_X78Y99_AO6),
.I2(CLBLM_R_X53Y99_SLICE_X80Y99_DO6),
.I3(CLBLM_R_X53Y99_SLICE_X81Y99_AO5),
.I4(CLBLM_R_X53Y99_SLICE_X81Y99_DO6),
.I5(CLBLM_R_X53Y99_SLICE_X80Y99_BO5),
.O5(CLBLM_R_X53Y99_SLICE_X81Y99_CO5),
.O6(CLBLM_R_X53Y99_SLICE_X81Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccdcccccffdcff)
  ) CLBLM_R_X53Y99_SLICE_X81Y99_BLUT (
.I0(CLBLM_R_X53Y99_SLICE_X80Y99_AO5),
.I1(CLBLL_L_X52Y99_SLICE_X79Y99_AO6),
.I2(CLBLM_R_X49Y107_SLICE_X75Y107_DQ),
.I3(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I4(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.I5(CLBLL_L_X54Y100_SLICE_X82Y100_AO5),
.O5(CLBLM_R_X53Y99_SLICE_X81Y99_BO5),
.O6(CLBLM_R_X53Y99_SLICE_X81Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0050000050000500)
  ) CLBLM_R_X53Y99_SLICE_X81Y99_ALUT (
.I0(CLBLM_R_X53Y99_SLICE_X80Y99_AO5),
.I1(1'b1),
.I2(CLBLM_R_X49Y107_SLICE_X75Y107_DQ),
.I3(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I4(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.I5(1'b1),
.O5(CLBLM_R_X53Y99_SLICE_X81Y99_AO5),
.O6(CLBLM_R_X53Y99_SLICE_X81Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X53Y100_SLICE_X80Y100_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X53Y100_SLICE_X80Y100_AO5),
.Q(CLBLM_R_X53Y100_SLICE_X80Y100_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X53Y100_SLICE_X80Y100_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X53Y100_SLICE_X80Y100_AO6),
.Q(CLBLM_R_X53Y100_SLICE_X80Y100_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaaafaaefaaafaaf)
  ) CLBLM_R_X53Y100_SLICE_X80Y100_DLUT (
.I0(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I1(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I2(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.I3(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.I4(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.I5(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.O5(CLBLM_R_X53Y100_SLICE_X80Y100_DO5),
.O6(CLBLM_R_X53Y100_SLICE_X80Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeeeeeeeeeeeeef)
  ) CLBLM_R_X53Y100_SLICE_X80Y100_CLUT (
.I0(CLBLM_L_X56Y99_SLICE_X84Y99_CO6),
.I1(CLBLL_R_X57Y102_SLICE_X86Y102_AO6),
.I2(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.I3(CLBLM_R_X53Y99_SLICE_X80Y99_BO6),
.I4(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I5(CLBLM_R_X49Y107_SLICE_X75Y107_DQ),
.O5(CLBLM_R_X53Y100_SLICE_X80Y100_CO5),
.O6(CLBLM_R_X53Y100_SLICE_X80Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdf000000200c0000)
  ) CLBLM_R_X53Y100_SLICE_X80Y100_BLUT (
.I0(CLBLM_R_X49Y108_SLICE_X75Y108_DQ),
.I1(CLBLM_R_X49Y107_SLICE_X75Y107_DQ),
.I2(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.I3(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I4(CLBLM_L_X56Y97_SLICE_X84Y97_CO5),
.I5(1'b1),
.O5(CLBLM_R_X53Y100_SLICE_X80Y100_BO5),
.O6(CLBLM_R_X53Y100_SLICE_X80Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffdcdcffddffdd)
  ) CLBLM_R_X53Y100_SLICE_X80Y100_ALUT (
.I0(CLBLM_R_X53Y100_SLICE_X80Y100_DO6),
.I1(CLBLM_R_X53Y99_SLICE_X80Y99_CO6),
.I2(CLBLM_R_X49Y107_SLICE_X75Y107_DQ),
.I3(CLBLM_R_X53Y100_SLICE_X80Y100_BO6),
.I4(CLBLM_R_X53Y100_SLICE_X80Y100_CO6),
.I5(1'b1),
.O5(CLBLM_R_X53Y100_SLICE_X80Y100_AO5),
.O6(CLBLM_R_X53Y100_SLICE_X80Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X53Y100_SLICE_X81Y100_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X53Y100_SLICE_X81Y100_AO6),
.Q(CLBLM_R_X53Y100_SLICE_X81Y100_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5400ffff00aa)
  ) CLBLM_R_X53Y100_SLICE_X81Y100_DLUT (
.I0(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I1(CLBLM_L_X56Y100_SLICE_X85Y100_AO5),
.I2(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.I3(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.I4(CLBLM_R_X53Y99_SLICE_X81Y99_AO5),
.I5(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.O5(CLBLM_R_X53Y100_SLICE_X81Y100_DO5),
.O6(CLBLM_R_X53Y100_SLICE_X81Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0100000000000000)
  ) CLBLM_R_X53Y100_SLICE_X81Y100_CLUT (
.I0(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I1(CLBLM_R_X49Y107_SLICE_X75Y107_DQ),
.I2(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.I3(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.I4(CLBLL_L_X54Y99_SLICE_X83Y99_BO5),
.I5(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.O5(CLBLM_R_X53Y100_SLICE_X81Y100_CO5),
.O6(CLBLM_R_X53Y100_SLICE_X81Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffff01)
  ) CLBLM_R_X53Y100_SLICE_X81Y100_BLUT (
.I0(CLBLM_R_X53Y100_SLICE_X81Y100_AO5),
.I1(CLBLM_R_X53Y99_SLICE_X80Y99_BO6),
.I2(CLBLM_R_X49Y107_SLICE_X75Y107_DQ),
.I3(CLBLL_R_X57Y102_SLICE_X86Y102_AO6),
.I4(CLBLM_L_X56Y99_SLICE_X84Y99_CO6),
.I5(CLBLM_R_X53Y100_SLICE_X81Y100_CO6),
.O5(CLBLM_R_X53Y100_SLICE_X81Y100_BO5),
.O6(CLBLM_R_X53Y100_SLICE_X81Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff11ff33fcfcfcfc)
  ) CLBLM_R_X53Y100_SLICE_X81Y100_ALUT (
.I0(CLBLL_L_X54Y100_SLICE_X82Y100_AO5),
.I1(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I2(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.I3(CLBLM_R_X53Y100_SLICE_X81Y100_BO6),
.I4(CLBLL_L_X54Y99_SLICE_X82Y99_BO6),
.I5(1'b1),
.O5(CLBLM_R_X53Y100_SLICE_X81Y100_AO5),
.O6(CLBLM_R_X53Y100_SLICE_X81Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X53Y101_SLICE_X80Y101_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X53Y101_SLICE_X80Y101_BO6),
.Q(CLBLM_R_X53Y101_SLICE_X80Y101_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0100000000000000)
  ) CLBLM_R_X53Y101_SLICE_X80Y101_DLUT (
.I0(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.I1(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I2(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.I3(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.I4(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.I5(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.O5(CLBLM_R_X53Y101_SLICE_X80Y101_DO5),
.O6(CLBLM_R_X53Y101_SLICE_X80Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0404101200001012)
  ) CLBLM_R_X53Y101_SLICE_X80Y101_CLUT (
.I0(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.I1(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.I2(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I3(CLBLM_R_X53Y100_SLICE_X81Y100_AO5),
.I4(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.I5(CLBLL_L_X54Y101_SLICE_X82Y101_AO5),
.O5(CLBLM_R_X53Y101_SLICE_X80Y101_CO5),
.O6(CLBLM_R_X53Y101_SLICE_X80Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X53Y101_SLICE_X80Y101_BLUT (
.I0(CLBLM_R_X53Y100_SLICE_X80Y100_BO5),
.I1(CLBLM_R_X53Y101_SLICE_X80Y101_DO6),
.I2(CLBLM_R_X53Y101_SLICE_X80Y101_CO6),
.I3(CLBLM_R_X53Y102_SLICE_X80Y102_AO6),
.I4(CLBLL_R_X57Y102_SLICE_X86Y102_AO6),
.I5(CLBLM_R_X53Y101_SLICE_X80Y101_AO5),
.O5(CLBLM_R_X53Y101_SLICE_X80Y101_BO5),
.O6(CLBLM_R_X53Y101_SLICE_X80Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h200020f001000100)
  ) CLBLM_R_X53Y101_SLICE_X80Y101_ALUT (
.I0(CLBLM_R_X49Y107_SLICE_X75Y107_DQ),
.I1(CLBLM_R_X53Y99_SLICE_X80Y99_BO6),
.I2(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.I3(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I4(CLBLM_R_X53Y99_SLICE_X80Y99_AO6),
.I5(1'b1),
.O5(CLBLM_R_X53Y101_SLICE_X80Y101_AO5),
.O6(CLBLM_R_X53Y101_SLICE_X80Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X53Y101_SLICE_X81Y101_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X53Y101_SLICE_X81Y101_AO6),
.Q(CLBLM_R_X53Y101_SLICE_X81Y101_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X53Y101_SLICE_X81Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X53Y101_SLICE_X81Y101_DO5),
.O6(CLBLM_R_X53Y101_SLICE_X81Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0002000800000000)
  ) CLBLM_R_X53Y101_SLICE_X81Y101_CLUT (
.I0(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.I1(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.I2(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I3(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.I4(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.I5(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.O5(CLBLM_R_X53Y101_SLICE_X81Y101_CO5),
.O6(CLBLM_R_X53Y101_SLICE_X81Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000100)
  ) CLBLM_R_X53Y101_SLICE_X81Y101_BLUT (
.I0(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I1(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.I2(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I3(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.I4(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.I5(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.O5(CLBLM_R_X53Y101_SLICE_X81Y101_BO5),
.O6(CLBLM_R_X53Y101_SLICE_X81Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X53Y101_SLICE_X81Y101_ALUT (
.I0(CLBLM_R_X53Y101_SLICE_X81Y101_BO6),
.I1(CLBLL_L_X52Y101_SLICE_X79Y101_AO6),
.I2(CLBLM_R_X53Y101_SLICE_X80Y101_AO6),
.I3(CLBLM_R_X53Y100_SLICE_X81Y100_BO6),
.I4(CLBLL_L_X54Y100_SLICE_X82Y100_DO6),
.I5(CLBLM_R_X53Y101_SLICE_X81Y101_CO6),
.O5(CLBLM_R_X53Y101_SLICE_X81Y101_AO5),
.O6(CLBLM_R_X53Y101_SLICE_X81Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X53Y102_SLICE_X80Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X53Y102_SLICE_X80Y102_DO5),
.O6(CLBLM_R_X53Y102_SLICE_X80Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X53Y102_SLICE_X80Y102_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X53Y102_SLICE_X80Y102_CO5),
.O6(CLBLM_R_X53Y102_SLICE_X80Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X53Y102_SLICE_X80Y102_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X53Y102_SLICE_X80Y102_BO5),
.O6(CLBLM_R_X53Y102_SLICE_X80Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0011044000010000)
  ) CLBLM_R_X53Y102_SLICE_X80Y102_ALUT (
.I0(CLBLM_R_X49Y106_SLICE_X75Y106_BQ),
.I1(CLBLM_R_X49Y104_SLICE_X74Y104_BQ),
.I2(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.I3(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I4(CLBLM_R_X49Y107_SLICE_X75Y107_BQ),
.I5(CLBLM_R_X49Y108_SLICE_X75Y108_CQ),
.O5(CLBLM_R_X53Y102_SLICE_X80Y102_AO5),
.O6(CLBLM_R_X53Y102_SLICE_X80Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X53Y102_SLICE_X81Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X53Y102_SLICE_X81Y102_DO5),
.O6(CLBLM_R_X53Y102_SLICE_X81Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X53Y102_SLICE_X81Y102_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X53Y102_SLICE_X81Y102_CO5),
.O6(CLBLM_R_X53Y102_SLICE_X81Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X53Y102_SLICE_X81Y102_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X53Y102_SLICE_X81Y102_BO5),
.O6(CLBLM_R_X53Y102_SLICE_X81Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X53Y102_SLICE_X81Y102_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X53Y102_SLICE_X81Y102_AO5),
.O6(CLBLM_R_X53Y102_SLICE_X81Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X53Y103_SLICE_X80Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X53Y103_SLICE_X80Y103_DO5),
.O6(CLBLM_R_X53Y103_SLICE_X80Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X53Y103_SLICE_X80Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X53Y103_SLICE_X80Y103_CO5),
.O6(CLBLM_R_X53Y103_SLICE_X80Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7888788878887888)
  ) CLBLM_R_X53Y103_SLICE_X80Y103_BLUT (
.I0(CLBLL_R_X57Y100_SLICE_X86Y100_AQ),
.I1(CLBLM_L_X56Y101_SLICE_X85Y101_CQ),
.I2(CLBLL_R_X57Y100_SLICE_X86Y100_CQ),
.I3(CLBLL_R_X57Y100_SLICE_X86Y100_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X53Y103_SLICE_X80Y103_BO5),
.O6(CLBLM_R_X53Y103_SLICE_X80Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h936c6c6c5fa0a0a0)
  ) CLBLM_R_X53Y103_SLICE_X80Y103_ALUT (
.I0(CLBLM_L_X56Y101_SLICE_X85Y101_AQ),
.I1(CLBLM_L_X56Y101_SLICE_X85Y101_CQ),
.I2(CLBLL_R_X57Y100_SLICE_X86Y100_CQ),
.I3(CLBLL_R_X57Y100_SLICE_X86Y100_DQ),
.I4(CLBLL_R_X57Y100_SLICE_X87Y100_AQ),
.I5(CLBLL_R_X57Y100_SLICE_X86Y100_BQ),
.O5(CLBLM_R_X53Y103_SLICE_X80Y103_AO5),
.O6(CLBLM_R_X53Y103_SLICE_X80Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X53Y103_SLICE_X81Y103_CARRY4 (
.CI(1'b0),
.CO({CLBLM_R_X53Y103_SLICE_X81Y103_D_CY, CLBLM_R_X53Y103_SLICE_X81Y103_C_CY, CLBLM_R_X53Y103_SLICE_X81Y103_B_CY, CLBLM_R_X53Y103_SLICE_X81Y103_A_CY}),
.CYINIT(1'b0),
.DI({CLBLM_R_X53Y103_SLICE_X80Y103_AO6, CLBLM_R_X53Y103_SLICE_X80Y103_BO6, CLBLM_R_X53Y103_SLICE_X81Y103_BO5, 1'b0}),
.O({CLBLM_R_X53Y103_SLICE_X81Y103_D_XOR, CLBLM_R_X53Y103_SLICE_X81Y103_C_XOR, CLBLM_R_X53Y103_SLICE_X81Y103_B_XOR, CLBLM_R_X53Y103_SLICE_X81Y103_A_XOR}),
.S({CLBLM_R_X53Y103_SLICE_X81Y103_DO6, CLBLM_R_X53Y103_SLICE_X81Y103_CO6, CLBLM_R_X53Y103_SLICE_X81Y103_BO6, CLBLM_R_X53Y103_SLICE_X81Y103_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h396c936cf5a05fa0)
  ) CLBLM_R_X53Y103_SLICE_X81Y103_DLUT (
.I0(CLBLL_R_X57Y100_SLICE_X86Y100_CQ),
.I1(CLBLL_R_X57Y100_SLICE_X87Y100_AQ),
.I2(CLBLM_L_X56Y101_SLICE_X85Y101_AQ),
.I3(CLBLL_L_X52Y105_SLICE_X78Y105_BO6),
.I4(CLBLL_R_X57Y100_SLICE_X86Y100_AQ),
.I5(CLBLL_R_X57Y100_SLICE_X86Y100_DQ),
.O5(CLBLM_R_X53Y103_SLICE_X81Y103_DO5),
.O6(CLBLM_R_X53Y103_SLICE_X81Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h953f6ac06ac06ac0)
  ) CLBLM_R_X53Y103_SLICE_X81Y103_CLUT (
.I0(CLBLL_R_X57Y100_SLICE_X86Y100_CQ),
.I1(CLBLL_R_X57Y100_SLICE_X86Y100_DQ),
.I2(CLBLM_L_X56Y101_SLICE_X85Y101_AQ),
.I3(CLBLL_R_X57Y100_SLICE_X86Y100_BQ),
.I4(CLBLL_R_X57Y100_SLICE_X86Y100_AQ),
.I5(CLBLM_L_X56Y101_SLICE_X85Y101_CQ),
.O5(CLBLM_R_X53Y103_SLICE_X81Y103_CO5),
.O6(CLBLM_R_X53Y103_SLICE_X81Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h66ccaa00cccc0000)
  ) CLBLM_R_X53Y103_SLICE_X81Y103_BLUT (
.I0(CLBLL_R_X57Y100_SLICE_X86Y100_BQ),
.I1(CLBLL_R_X57Y100_SLICE_X86Y100_AQ),
.I2(1'b1),
.I3(CLBLL_R_X57Y100_SLICE_X86Y100_DQ),
.I4(CLBLL_R_X57Y100_SLICE_X86Y100_CQ),
.I5(1'b1),
.O5(CLBLM_R_X53Y103_SLICE_X81Y103_BO5),
.O6(CLBLM_R_X53Y103_SLICE_X81Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00000000)
  ) CLBLM_R_X53Y103_SLICE_X81Y103_ALUT (
.I0(1'b1),
.I1(CLBLL_R_X57Y100_SLICE_X86Y100_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_R_X57Y100_SLICE_X86Y100_AQ),
.O5(CLBLM_R_X53Y103_SLICE_X81Y103_AO5),
.O6(CLBLM_R_X53Y103_SLICE_X81Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000a0a0a0a0)
  ) CLBLM_R_X53Y104_SLICE_X80Y104_DLUT (
.I0(CLBLM_L_X56Y101_SLICE_X85Y101_AQ),
.I1(1'b1),
.I2(CLBLM_L_X56Y101_SLICE_X85Y101_CQ),
.I3(CLBLL_R_X57Y100_SLICE_X86Y100_CQ),
.I4(CLBLL_R_X57Y100_SLICE_X87Y100_BQ),
.I5(1'b1),
.O5(CLBLM_R_X53Y104_SLICE_X80Y104_DO5),
.O6(CLBLM_R_X53Y104_SLICE_X80Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heac0800080008000)
  ) CLBLM_R_X53Y104_SLICE_X80Y104_CLUT (
.I0(CLBLM_L_X56Y101_SLICE_X85Y101_AQ),
.I1(CLBLL_R_X57Y100_SLICE_X87Y100_AQ),
.I2(CLBLL_R_X57Y100_SLICE_X86Y100_DQ),
.I3(CLBLL_R_X57Y100_SLICE_X86Y100_CQ),
.I4(CLBLM_L_X56Y101_SLICE_X85Y101_CQ),
.I5(CLBLL_R_X57Y100_SLICE_X86Y100_BQ),
.O5(CLBLM_R_X53Y104_SLICE_X80Y104_CO5),
.O6(CLBLM_R_X53Y104_SLICE_X80Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf880808088000000)
  ) CLBLM_R_X53Y104_SLICE_X80Y104_BLUT (
.I0(CLBLL_R_X57Y101_SLICE_X87Y101_AQ),
.I1(CLBLL_R_X57Y100_SLICE_X86Y100_DQ),
.I2(CLBLL_R_X57Y100_SLICE_X86Y100_CQ),
.I3(CLBLM_L_X56Y101_SLICE_X85Y101_CQ),
.I4(CLBLM_L_X56Y101_SLICE_X85Y101_AQ),
.I5(CLBLL_R_X57Y100_SLICE_X87Y100_AQ),
.O5(CLBLM_R_X53Y104_SLICE_X80Y104_BO5),
.O6(CLBLM_R_X53Y104_SLICE_X80Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00aa00aa00)
  ) CLBLM_R_X53Y104_SLICE_X80Y104_ALUT (
.I0(CLBLL_R_X57Y101_SLICE_X87Y101_AQ),
.I1(CLBLM_L_X56Y101_SLICE_X85Y101_BQ),
.I2(1'b1),
.I3(CLBLL_R_X57Y100_SLICE_X86Y100_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X53Y104_SLICE_X80Y104_AO5),
.O6(CLBLM_R_X53Y104_SLICE_X80Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X53Y104_SLICE_X81Y104_CARRY4 (
.CI(CLBLM_R_X53Y103_SLICE_X81Y103_COUT),
.CO({CLBLM_R_X53Y104_SLICE_X81Y104_D_CY, CLBLM_R_X53Y104_SLICE_X81Y104_C_CY, CLBLM_R_X53Y104_SLICE_X81Y104_B_CY, CLBLM_R_X53Y104_SLICE_X81Y104_A_CY}),
.CYINIT(1'b0),
.DI({CLBLL_L_X54Y104_SLICE_X82Y104_BO6, CLBLL_L_X54Y104_SLICE_X82Y104_AO6, CLBLM_R_X53Y104_SLICE_X80Y104_BO6, CLBLM_R_X53Y104_SLICE_X80Y104_CO6}),
.O({CLBLM_R_X53Y104_SLICE_X81Y104_D_XOR, CLBLM_R_X53Y104_SLICE_X81Y104_C_XOR, CLBLM_R_X53Y104_SLICE_X81Y104_B_XOR, CLBLM_R_X53Y104_SLICE_X81Y104_A_XOR}),
.S({CLBLM_R_X53Y104_SLICE_X81Y104_DO6, CLBLM_R_X53Y104_SLICE_X81Y104_CO6, CLBLM_R_X53Y104_SLICE_X81Y104_BO6, CLBLM_R_X53Y104_SLICE_X81Y104_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h69a5965ac30f3cf0)
  ) CLBLM_R_X53Y104_SLICE_X81Y104_DLUT (
.I0(CLBLL_R_X57Y100_SLICE_X86Y100_DQ),
.I1(CLBLM_L_X56Y101_SLICE_X85Y101_CQ),
.I2(CLBLM_R_X53Y104_SLICE_X80Y104_DO6),
.I3(CLBLM_L_X56Y101_SLICE_X85Y101_BQ),
.I4(CLBLL_L_X54Y104_SLICE_X82Y104_BO6),
.I5(CLBLL_R_X57Y99_SLICE_X86Y99_AQ),
.O5(CLBLM_R_X53Y104_SLICE_X81Y104_DO5),
.O6(CLBLM_R_X53Y104_SLICE_X81Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a95956ac03f3fc0)
  ) CLBLM_R_X53Y104_SLICE_X81Y104_CLUT (
.I0(CLBLL_R_X57Y100_SLICE_X86Y100_DQ),
.I1(CLBLM_L_X56Y101_SLICE_X85Y101_CQ),
.I2(CLBLL_R_X57Y101_SLICE_X87Y101_AQ),
.I3(CLBLL_L_X54Y104_SLICE_X82Y104_AO6),
.I4(CLBLM_R_X53Y104_SLICE_X80Y104_AO6),
.I5(CLBLL_R_X57Y100_SLICE_X87Y100_BQ),
.O5(CLBLM_R_X53Y104_SLICE_X81Y104_CO5),
.O6(CLBLM_R_X53Y104_SLICE_X81Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996c33c96963c3c)
  ) CLBLM_R_X53Y104_SLICE_X81Y104_BLUT (
.I0(CLBLM_L_X56Y101_SLICE_X85Y101_BQ),
.I1(CLBLM_R_X53Y104_SLICE_X80Y104_BO6),
.I2(CLBLM_R_X53Y104_SLICE_X80Y104_AO5),
.I3(CLBLM_L_X56Y101_SLICE_X85Y101_CQ),
.I4(CLBLL_R_X57Y100_SLICE_X86Y100_DQ),
.I5(CLBLL_R_X57Y100_SLICE_X87Y100_AQ),
.O5(CLBLM_R_X53Y104_SLICE_X81Y104_BO5),
.O6(CLBLM_R_X53Y104_SLICE_X81Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3963c963c963c)
  ) CLBLM_R_X53Y104_SLICE_X81Y104_ALUT (
.I0(CLBLL_R_X57Y101_SLICE_X87Y101_AQ),
.I1(CLBLM_R_X53Y104_SLICE_X80Y104_DO5),
.I2(CLBLM_R_X53Y104_SLICE_X80Y104_CO6),
.I3(CLBLL_R_X57Y100_SLICE_X86Y100_DQ),
.I4(CLBLL_R_X57Y100_SLICE_X86Y100_CQ),
.I5(CLBLL_R_X57Y100_SLICE_X87Y100_AQ),
.O5(CLBLM_R_X53Y104_SLICE_X81Y104_AO5),
.O6(CLBLM_R_X53Y104_SLICE_X81Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X53Y105_SLICE_X80Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X53Y105_SLICE_X80Y105_DO5),
.O6(CLBLM_R_X53Y105_SLICE_X80Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X53Y105_SLICE_X80Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X53Y105_SLICE_X80Y105_CO5),
.O6(CLBLM_R_X53Y105_SLICE_X80Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he8c0a00088000000)
  ) CLBLM_R_X53Y105_SLICE_X80Y105_BLUT (
.I0(CLBLM_L_X56Y101_SLICE_X85Y101_CQ),
.I1(CLBLL_R_X57Y100_SLICE_X86Y100_DQ),
.I2(CLBLL_R_X57Y100_SLICE_X86Y100_CQ),
.I3(CLBLM_L_X56Y101_SLICE_X85Y101_BQ),
.I4(CLBLL_R_X57Y99_SLICE_X86Y99_AQ),
.I5(CLBLL_R_X57Y100_SLICE_X87Y100_BQ),
.O5(CLBLM_R_X53Y105_SLICE_X80Y105_BO5),
.O6(CLBLM_R_X53Y105_SLICE_X80Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he800a000a000a000)
  ) CLBLM_R_X53Y105_SLICE_X80Y105_ALUT (
.I0(CLBLM_L_X56Y101_SLICE_X85Y101_AQ),
.I1(CLBLM_R_X53Y106_SLICE_X81Y106_D_XOR),
.I2(CLBLM_R_X53Y106_SLICE_X80Y106_AO5),
.I3(CLBLL_R_X57Y101_SLICE_X87Y101_DQ),
.I4(CLBLM_R_X53Y104_SLICE_X81Y104_C_XOR),
.I5(CLBLL_R_X57Y100_SLICE_X86Y100_BQ),
.O5(CLBLM_R_X53Y105_SLICE_X80Y105_AO5),
.O6(CLBLM_R_X53Y105_SLICE_X80Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X53Y105_SLICE_X81Y105_CARRY4 (
.CI(CLBLM_R_X53Y104_SLICE_X81Y104_COUT),
.CO({CLBLM_R_X53Y105_SLICE_X81Y105_D_CY, CLBLM_R_X53Y105_SLICE_X81Y105_C_CY, CLBLM_R_X53Y105_SLICE_X81Y105_B_CY, CLBLM_R_X53Y105_SLICE_X81Y105_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, CLBLM_R_X53Y105_SLICE_X81Y105_BO5, CLBLM_R_X53Y105_SLICE_X80Y105_BO6}),
.O({CLBLM_R_X53Y105_SLICE_X81Y105_D_XOR, CLBLM_R_X53Y105_SLICE_X81Y105_C_XOR, CLBLM_R_X53Y105_SLICE_X81Y105_B_XOR, CLBLM_R_X53Y105_SLICE_X81Y105_A_XOR}),
.S({CLBLM_R_X53Y105_SLICE_X81Y105_DO6, CLBLM_R_X53Y105_SLICE_X81Y105_CO6, CLBLM_R_X53Y105_SLICE_X81Y105_BO6, CLBLM_R_X53Y105_SLICE_X81Y105_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X53Y105_SLICE_X81Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X53Y105_SLICE_X81Y105_DO5),
.O6(CLBLM_R_X53Y105_SLICE_X81Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffff)
  ) CLBLM_R_X53Y105_SLICE_X81Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X53Y105_SLICE_X81Y105_CO5),
.O6(CLBLM_R_X53Y105_SLICE_X81Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h30f00000f0f00000)
  ) CLBLM_R_X53Y105_SLICE_X81Y105_BLUT (
.I0(1'b1),
.I1(CLBLL_R_X57Y100_SLICE_X87Y100_BQ),
.I2(CLBLL_R_X57Y99_SLICE_X86Y99_AQ),
.I3(CLBLL_R_X57Y100_SLICE_X86Y100_CQ),
.I4(CLBLM_L_X56Y101_SLICE_X85Y101_CQ),
.I5(1'b1),
.O5(CLBLM_R_X53Y105_SLICE_X81Y105_BO5),
.O6(CLBLM_R_X53Y105_SLICE_X81Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h90f02888b8788888)
  ) CLBLM_R_X53Y105_SLICE_X81Y105_ALUT (
.I0(CLBLM_L_X56Y101_SLICE_X85Y101_CQ),
.I1(CLBLL_R_X57Y100_SLICE_X87Y100_BQ),
.I2(CLBLL_R_X57Y99_SLICE_X86Y99_AQ),
.I3(CLBLL_R_X57Y100_SLICE_X86Y100_DQ),
.I4(CLBLL_R_X57Y100_SLICE_X86Y100_CQ),
.I5(CLBLM_L_X56Y101_SLICE_X85Y101_BQ),
.O5(CLBLM_R_X53Y105_SLICE_X81Y105_AO5),
.O6(CLBLM_R_X53Y105_SLICE_X81Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00aa00aa00)
  ) CLBLM_R_X53Y106_SLICE_X80Y106_DLUT (
.I0(CLBLL_R_X57Y100_SLICE_X86Y100_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X56Y101_SLICE_X85Y101_DQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X53Y106_SLICE_X80Y106_DO5),
.O6(CLBLM_R_X53Y106_SLICE_X80Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8777788878887888)
  ) CLBLM_R_X53Y106_SLICE_X80Y106_CLUT (
.I0(CLBLL_R_X57Y100_SLICE_X86Y100_BQ),
.I1(CLBLM_L_X56Y101_SLICE_X85Y101_DQ),
.I2(CLBLL_R_X57Y100_SLICE_X87Y100_AQ),
.I3(CLBLL_R_X57Y100_SLICE_X87Y100_CQ),
.I4(CLBLL_R_X57Y101_SLICE_X87Y101_CQ),
.I5(CLBLM_L_X56Y101_SLICE_X85Y101_AQ),
.O5(CLBLM_R_X53Y106_SLICE_X80Y106_CO5),
.O6(CLBLM_R_X53Y106_SLICE_X80Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h80ff7fff7f008000)
  ) CLBLM_R_X53Y106_SLICE_X80Y106_BLUT (
.I0(CLBLL_R_X57Y100_SLICE_X86Y100_BQ),
.I1(CLBLM_R_X53Y106_SLICE_X81Y106_D_XOR),
.I2(CLBLM_R_X53Y104_SLICE_X81Y104_C_XOR),
.I3(CLBLL_R_X57Y101_SLICE_X87Y101_DQ),
.I4(CLBLM_L_X56Y101_SLICE_X85Y101_AQ),
.I5(CLBLM_R_X53Y106_SLICE_X80Y106_AO5),
.O5(CLBLM_R_X53Y106_SLICE_X80Y106_BO5),
.O6(CLBLM_R_X53Y106_SLICE_X80Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h1777177796669666)
  ) CLBLM_R_X53Y106_SLICE_X80Y106_ALUT (
.I0(CLBLM_R_X53Y107_SLICE_X81Y107_B_XOR),
.I1(CLBLM_R_X53Y105_SLICE_X81Y105_A_XOR),
.I2(CLBLL_R_X57Y100_SLICE_X86Y100_BQ),
.I3(CLBLL_R_X57Y99_SLICE_X86Y99_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X53Y106_SLICE_X80Y106_AO5),
.O6(CLBLM_R_X53Y106_SLICE_X80Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X53Y106_SLICE_X81Y106_CARRY4 (
.CI(1'b0),
.CO({CLBLM_R_X53Y106_SLICE_X81Y106_D_CY, CLBLM_R_X53Y106_SLICE_X81Y106_C_CY, CLBLM_R_X53Y106_SLICE_X81Y106_B_CY, CLBLM_R_X53Y106_SLICE_X81Y106_A_CY}),
.CYINIT(1'b0),
.DI({CLBLM_R_X53Y106_SLICE_X80Y106_CO6, CLBLL_L_X52Y106_SLICE_X79Y106_BO6, CLBLM_R_X53Y106_SLICE_X81Y106_BO5, 1'b0}),
.O({CLBLM_R_X53Y106_SLICE_X81Y106_D_XOR, CLBLM_R_X53Y106_SLICE_X81Y106_C_XOR, CLBLM_R_X53Y106_SLICE_X81Y106_B_XOR, CLBLM_R_X53Y106_SLICE_X81Y106_A_XOR}),
.S({CLBLM_R_X53Y106_SLICE_X81Y106_DO6, CLBLM_R_X53Y106_SLICE_X81Y106_CO6, CLBLM_R_X53Y106_SLICE_X81Y106_BO6, CLBLM_R_X53Y106_SLICE_X81Y106_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7787787888787878)
  ) CLBLM_R_X53Y106_SLICE_X81Y106_DLUT (
.I0(CLBLL_R_X57Y100_SLICE_X87Y100_CQ),
.I1(CLBLL_R_X57Y100_SLICE_X87Y100_AQ),
.I2(CLBLM_R_X53Y106_SLICE_X80Y106_DO6),
.I3(CLBLL_R_X57Y100_SLICE_X86Y100_AQ),
.I4(CLBLL_R_X57Y101_SLICE_X87Y101_CQ),
.I5(CLBLM_L_X56Y101_SLICE_X85Y101_AQ),
.O5(CLBLM_R_X53Y106_SLICE_X81Y106_DO5),
.O6(CLBLM_R_X53Y106_SLICE_X81Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h936c6c6c5fa0a0a0)
  ) CLBLM_R_X53Y106_SLICE_X81Y106_CLUT (
.I0(CLBLL_R_X57Y100_SLICE_X86Y100_BQ),
.I1(CLBLL_R_X57Y100_SLICE_X87Y100_CQ),
.I2(CLBLL_R_X57Y101_SLICE_X87Y101_CQ),
.I3(CLBLM_L_X56Y101_SLICE_X85Y101_DQ),
.I4(CLBLL_R_X57Y100_SLICE_X86Y100_AQ),
.I5(CLBLM_L_X56Y101_SLICE_X85Y101_AQ),
.O5(CLBLM_R_X53Y106_SLICE_X81Y106_CO5),
.O6(CLBLM_R_X53Y106_SLICE_X81Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cccf000f000f000)
  ) CLBLM_R_X53Y106_SLICE_X81Y106_BLUT (
.I0(1'b1),
.I1(CLBLL_R_X57Y100_SLICE_X87Y100_CQ),
.I2(CLBLL_R_X57Y100_SLICE_X86Y100_AQ),
.I3(CLBLL_R_X57Y101_SLICE_X87Y101_CQ),
.I4(CLBLL_R_X57Y100_SLICE_X86Y100_BQ),
.I5(1'b1),
.O5(CLBLM_R_X53Y106_SLICE_X81Y106_BO5),
.O6(CLBLM_R_X53Y106_SLICE_X81Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0c0c0c0c0)
  ) CLBLM_R_X53Y106_SLICE_X81Y106_ALUT (
.I0(1'b1),
.I1(CLBLL_R_X57Y100_SLICE_X87Y100_CQ),
.I2(CLBLL_R_X57Y100_SLICE_X86Y100_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X53Y106_SLICE_X81Y106_AO5),
.O6(CLBLM_R_X53Y106_SLICE_X81Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he888c000a0000000)
  ) CLBLM_R_X53Y107_SLICE_X80Y107_DLUT (
.I0(CLBLL_R_X57Y100_SLICE_X87Y100_AQ),
.I1(CLBLL_R_X57Y100_SLICE_X87Y100_CQ),
.I2(CLBLL_R_X57Y101_SLICE_X87Y101_AQ),
.I3(CLBLL_R_X57Y101_SLICE_X87Y101_CQ),
.I4(CLBLM_L_X56Y101_SLICE_X85Y101_DQ),
.I5(CLBLM_L_X56Y101_SLICE_X85Y101_BQ),
.O5(CLBLM_R_X53Y107_SLICE_X80Y107_DO5),
.O6(CLBLM_R_X53Y107_SLICE_X80Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf880880080800000)
  ) CLBLM_R_X53Y107_SLICE_X80Y107_CLUT (
.I0(CLBLL_R_X57Y100_SLICE_X87Y100_BQ),
.I1(CLBLL_R_X57Y100_SLICE_X87Y100_CQ),
.I2(CLBLL_R_X57Y101_SLICE_X87Y101_AQ),
.I3(CLBLM_L_X56Y101_SLICE_X85Y101_BQ),
.I4(CLBLM_L_X56Y101_SLICE_X85Y101_DQ),
.I5(CLBLL_R_X57Y101_SLICE_X87Y101_CQ),
.O5(CLBLM_R_X53Y107_SLICE_X80Y107_CO5),
.O6(CLBLM_R_X53Y107_SLICE_X80Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h13137f7f93936c6c)
  ) CLBLM_R_X53Y107_SLICE_X80Y107_BLUT (
.I0(CLBLL_R_X57Y100_SLICE_X87Y100_AQ),
.I1(CLBLM_R_X53Y107_SLICE_X81Y107_D_XOR),
.I2(CLBLL_R_X57Y99_SLICE_X86Y99_BQ),
.I3(1'b1),
.I4(CLBLM_R_X53Y105_SLICE_X81Y105_C_CY),
.I5(1'b1),
.O5(CLBLM_R_X53Y107_SLICE_X80Y107_BO5),
.O6(CLBLM_R_X53Y107_SLICE_X80Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000f0f00000)
  ) CLBLM_R_X53Y107_SLICE_X80Y107_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_R_X57Y100_SLICE_X87Y100_AQ),
.I3(CLBLM_L_X56Y101_SLICE_X85Y101_BQ),
.I4(CLBLL_R_X57Y101_SLICE_X87Y101_CQ),
.I5(1'b1),
.O5(CLBLM_R_X53Y107_SLICE_X80Y107_AO5),
.O6(CLBLM_R_X53Y107_SLICE_X80Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X53Y107_SLICE_X81Y107_CARRY4 (
.CI(CLBLM_R_X53Y106_SLICE_X81Y106_COUT),
.CO({CLBLM_R_X53Y107_SLICE_X81Y107_D_CY, CLBLM_R_X53Y107_SLICE_X81Y107_C_CY, CLBLM_R_X53Y107_SLICE_X81Y107_B_CY, CLBLM_R_X53Y107_SLICE_X81Y107_A_CY}),
.CYINIT(1'b0),
.DI({CLBLM_R_X53Y107_SLICE_X80Y107_CO6, CLBLM_R_X53Y107_SLICE_X80Y107_DO6, CLBLM_R_X53Y108_SLICE_X80Y108_AO6, CLBLM_R_X53Y108_SLICE_X80Y108_BO6}),
.O({CLBLM_R_X53Y107_SLICE_X81Y107_D_XOR, CLBLM_R_X53Y107_SLICE_X81Y107_C_XOR, CLBLM_R_X53Y107_SLICE_X81Y107_B_XOR, CLBLM_R_X53Y107_SLICE_X81Y107_A_XOR}),
.S({CLBLM_R_X53Y107_SLICE_X81Y107_DO6, CLBLM_R_X53Y107_SLICE_X81Y107_CO6, CLBLM_R_X53Y107_SLICE_X81Y107_BO6, CLBLM_R_X53Y107_SLICE_X81Y107_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h69a5c30f965a3cf0)
  ) CLBLM_R_X53Y107_SLICE_X81Y107_DLUT (
.I0(CLBLL_R_X57Y100_SLICE_X87Y100_CQ),
.I1(CLBLL_R_X57Y101_SLICE_X87Y101_CQ),
.I2(CLBLM_R_X53Y107_SLICE_X80Y107_CO6),
.I3(CLBLL_R_X57Y100_SLICE_X87Y100_BQ),
.I4(CLBLL_R_X57Y99_SLICE_X86Y99_AQ),
.I5(CLBLL_L_X52Y107_SLICE_X78Y107_AO6),
.O5(CLBLM_R_X53Y107_SLICE_X81Y107_DO5),
.O6(CLBLM_R_X53Y107_SLICE_X81Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a95956ac03f3fc0)
  ) CLBLM_R_X53Y107_SLICE_X81Y107_CLUT (
.I0(CLBLL_R_X57Y100_SLICE_X87Y100_CQ),
.I1(CLBLM_L_X56Y101_SLICE_X85Y101_DQ),
.I2(CLBLL_R_X57Y101_SLICE_X87Y101_AQ),
.I3(CLBLM_R_X53Y107_SLICE_X80Y107_DO6),
.I4(CLBLM_R_X53Y107_SLICE_X80Y107_AO6),
.I5(CLBLL_R_X57Y100_SLICE_X87Y100_BQ),
.O5(CLBLM_R_X53Y107_SLICE_X81Y107_CO5),
.O6(CLBLM_R_X53Y107_SLICE_X81Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69969696c33c3c3c)
  ) CLBLM_R_X53Y107_SLICE_X81Y107_BLUT (
.I0(CLBLM_L_X56Y101_SLICE_X85Y101_BQ),
.I1(CLBLM_R_X53Y108_SLICE_X80Y108_AO6),
.I2(CLBLL_L_X52Y106_SLICE_X79Y106_AO6),
.I3(CLBLM_L_X56Y101_SLICE_X85Y101_DQ),
.I4(CLBLL_R_X57Y100_SLICE_X87Y100_AQ),
.I5(CLBLL_R_X57Y100_SLICE_X87Y100_CQ),
.O5(CLBLM_R_X53Y107_SLICE_X81Y107_BO5),
.O6(CLBLM_R_X53Y107_SLICE_X81Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3a50f963c5af0)
  ) CLBLM_R_X53Y107_SLICE_X81Y107_ALUT (
.I0(CLBLL_R_X57Y101_SLICE_X87Y101_AQ),
.I1(CLBLM_L_X56Y101_SLICE_X85Y101_DQ),
.I2(CLBLM_R_X53Y107_SLICE_X80Y107_AO5),
.I3(CLBLL_R_X57Y100_SLICE_X87Y100_CQ),
.I4(CLBLM_L_X56Y101_SLICE_X85Y101_AQ),
.I5(CLBLM_R_X53Y108_SLICE_X80Y108_BO6),
.O5(CLBLM_R_X53Y107_SLICE_X81Y107_AO5),
.O6(CLBLM_R_X53Y107_SLICE_X81Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X53Y108_SLICE_X80Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X53Y108_SLICE_X80Y108_DO5),
.O6(CLBLM_R_X53Y108_SLICE_X80Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heac0800080008000)
  ) CLBLM_R_X53Y108_SLICE_X80Y108_CLUT (
.I0(CLBLM_L_X56Y101_SLICE_X85Y101_DQ),
.I1(CLBLL_R_X57Y100_SLICE_X87Y100_BQ),
.I2(CLBLL_R_X57Y101_SLICE_X87Y101_CQ),
.I3(CLBLM_L_X56Y101_SLICE_X85Y101_BQ),
.I4(CLBLL_R_X57Y100_SLICE_X87Y100_CQ),
.I5(CLBLL_R_X57Y99_SLICE_X86Y99_AQ),
.O5(CLBLM_R_X53Y108_SLICE_X80Y108_CO5),
.O6(CLBLM_R_X53Y108_SLICE_X80Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he8c0a00088000000)
  ) CLBLM_R_X53Y108_SLICE_X80Y108_BLUT (
.I0(CLBLL_R_X57Y100_SLICE_X87Y100_AQ),
.I1(CLBLL_R_X57Y100_SLICE_X86Y100_BQ),
.I2(CLBLM_L_X56Y101_SLICE_X85Y101_AQ),
.I3(CLBLL_R_X57Y100_SLICE_X87Y100_CQ),
.I4(CLBLM_L_X56Y101_SLICE_X85Y101_DQ),
.I5(CLBLL_R_X57Y101_SLICE_X87Y101_CQ),
.O5(CLBLM_R_X53Y108_SLICE_X80Y108_BO5),
.O6(CLBLM_R_X53Y108_SLICE_X80Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hec80a00080800000)
  ) CLBLM_R_X53Y108_SLICE_X80Y108_ALUT (
.I0(CLBLM_L_X56Y101_SLICE_X85Y101_DQ),
.I1(CLBLL_R_X57Y101_SLICE_X87Y101_CQ),
.I2(CLBLM_L_X56Y101_SLICE_X85Y101_AQ),
.I3(CLBLL_R_X57Y101_SLICE_X87Y101_AQ),
.I4(CLBLL_R_X57Y100_SLICE_X87Y100_AQ),
.I5(CLBLL_R_X57Y100_SLICE_X87Y100_CQ),
.O5(CLBLM_R_X53Y108_SLICE_X80Y108_AO5),
.O6(CLBLM_R_X53Y108_SLICE_X80Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X53Y108_SLICE_X81Y108_CARRY4 (
.CI(CLBLM_R_X53Y107_SLICE_X81Y107_COUT),
.CO({CLBLM_R_X53Y108_SLICE_X81Y108_D_CY, CLBLM_R_X53Y108_SLICE_X81Y108_C_CY, CLBLM_R_X53Y108_SLICE_X81Y108_B_CY, CLBLM_R_X53Y108_SLICE_X81Y108_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, CLBLM_R_X53Y108_SLICE_X81Y108_BO5, CLBLM_R_X53Y108_SLICE_X80Y108_CO6}),
.O({CLBLM_R_X53Y108_SLICE_X81Y108_D_XOR, CLBLM_R_X53Y108_SLICE_X81Y108_C_XOR, CLBLM_R_X53Y108_SLICE_X81Y108_B_XOR, CLBLM_R_X53Y108_SLICE_X81Y108_A_XOR}),
.S({CLBLM_R_X53Y108_SLICE_X81Y108_DO6, CLBLM_R_X53Y108_SLICE_X81Y108_CO6, CLBLM_R_X53Y108_SLICE_X81Y108_BO6, CLBLM_R_X53Y108_SLICE_X81Y108_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X53Y108_SLICE_X81Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X53Y108_SLICE_X81Y108_DO5),
.O6(CLBLM_R_X53Y108_SLICE_X81Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffff)
  ) CLBLM_R_X53Y108_SLICE_X81Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X53Y108_SLICE_X81Y108_CO5),
.O6(CLBLM_R_X53Y108_SLICE_X81Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4040c0c0c0c0c0c0)
  ) CLBLM_R_X53Y108_SLICE_X81Y108_BLUT (
.I0(CLBLL_R_X57Y101_SLICE_X87Y101_CQ),
.I1(CLBLL_R_X57Y99_SLICE_X86Y99_AQ),
.I2(CLBLM_L_X56Y101_SLICE_X85Y101_DQ),
.I3(1'b1),
.I4(CLBLL_R_X57Y100_SLICE_X87Y100_BQ),
.I5(1'b1),
.O5(CLBLM_R_X53Y108_SLICE_X81Y108_BO5),
.O6(CLBLM_R_X53Y108_SLICE_X81Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc4704c80b4f0cc00)
  ) CLBLM_R_X53Y108_SLICE_X81Y108_ALUT (
.I0(CLBLL_R_X57Y100_SLICE_X87Y100_CQ),
.I1(CLBLL_R_X57Y99_SLICE_X86Y99_AQ),
.I2(CLBLM_L_X56Y101_SLICE_X85Y101_DQ),
.I3(CLBLL_R_X57Y101_SLICE_X87Y101_CQ),
.I4(CLBLL_R_X57Y100_SLICE_X87Y100_BQ),
.I5(CLBLM_L_X56Y101_SLICE_X85Y101_BQ),
.O5(CLBLM_R_X53Y108_SLICE_X81Y108_AO5),
.O6(CLBLM_R_X53Y108_SLICE_X81Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y96_SLICE_X88Y96_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y96_SLICE_X88Y96_AO6),
.Q(CLBLM_R_X59Y96_SLICE_X88Y96_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y96_SLICE_X88Y96_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y96_SLICE_X88Y96_BO6),
.Q(CLBLM_R_X59Y96_SLICE_X88Y96_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff10ff00ff02)
  ) CLBLM_R_X59Y96_SLICE_X88Y96_DLUT (
.I0(CLBLM_L_X50Y107_SLICE_X77Y107_AQ),
.I1(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I2(CLBLL_R_X57Y99_SLICE_X86Y99_AQ),
.I3(CLBLM_R_X59Y96_SLICE_X89Y96_BO6),
.I4(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I5(CLBLL_R_X57Y99_SLICE_X86Y99_BQ),
.O5(CLBLM_R_X59Y96_SLICE_X88Y96_DO5),
.O6(CLBLM_R_X59Y96_SLICE_X88Y96_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000faca00000aca)
  ) CLBLM_R_X59Y96_SLICE_X88Y96_CLUT (
.I0(CLBLM_L_X50Y107_SLICE_X77Y107_AQ),
.I1(CLBLM_R_X59Y96_SLICE_X88Y96_AQ),
.I2(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I3(CLBLL_R_X57Y97_SLICE_X86Y97_CO6),
.I4(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I5(CLBLM_R_X59Y97_SLICE_X89Y97_B5Q),
.O5(CLBLM_R_X59Y96_SLICE_X88Y96_CO5),
.O6(CLBLM_R_X59Y96_SLICE_X88Y96_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffe0ccccff40cccc)
  ) CLBLM_R_X59Y96_SLICE_X88Y96_BLUT (
.I0(CLBLM_L_X60Y99_SLICE_X91Y99_DO6),
.I1(CLBLM_R_X59Y96_SLICE_X88Y96_BQ),
.I2(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I3(CLBLM_R_X59Y96_SLICE_X88Y96_DO6),
.I4(CLBLL_R_X57Y98_SLICE_X86Y98_BO6),
.I5(CLBLM_R_X49Y106_SLICE_X74Y106_AQ),
.O5(CLBLM_R_X59Y96_SLICE_X88Y96_BO5),
.O6(CLBLM_R_X59Y96_SLICE_X88Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcfcfcb830b0b0)
  ) CLBLM_R_X59Y96_SLICE_X88Y96_ALUT (
.I0(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I1(CLBLL_R_X57Y98_SLICE_X86Y98_CO6),
.I2(CLBLM_R_X59Y96_SLICE_X88Y96_AQ),
.I3(CLBLM_L_X50Y106_SLICE_X76Y106_AQ),
.I4(CLBLM_L_X60Y99_SLICE_X91Y99_DO6),
.I5(CLBLM_R_X59Y96_SLICE_X88Y96_CO6),
.O5(CLBLM_R_X59Y96_SLICE_X88Y96_AO5),
.O6(CLBLM_R_X59Y96_SLICE_X88Y96_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y96_SLICE_X89Y96_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_R_X59Y98_SLICE_X89Y98_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y96_SLICE_X89Y96_AO5),
.Q(CLBLM_R_X59Y96_SLICE_X89Y96_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y96_SLICE_X89Y96_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_R_X59Y98_SLICE_X89Y98_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y96_SLICE_X89Y96_AO6),
.Q(CLBLM_R_X59Y96_SLICE_X89Y96_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X59Y96_SLICE_X89Y96_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y96_SLICE_X89Y96_DO5),
.O6(CLBLM_R_X59Y96_SLICE_X89Y96_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X59Y96_SLICE_X89Y96_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y96_SLICE_X89Y96_CO5),
.O6(CLBLM_R_X59Y96_SLICE_X89Y96_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aa2000008a00)
  ) CLBLM_R_X59Y96_SLICE_X89Y96_BLUT (
.I0(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I1(CLBLM_L_X56Y98_SLICE_X85Y98_CQ),
.I2(CLBLM_L_X56Y98_SLICE_X85Y98_BQ),
.I3(CLBLM_R_X59Y96_SLICE_X88Y96_BQ),
.I4(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I5(CLBLM_R_X59Y97_SLICE_X89Y97_A5Q),
.O5(CLBLM_R_X59Y96_SLICE_X89Y96_BO5),
.O6(CLBLM_R_X59Y96_SLICE_X89Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8d8d8ff55aa00)
  ) CLBLM_R_X59Y96_SLICE_X89Y96_ALUT (
.I0(CLBLM_L_X60Y98_SLICE_X90Y98_DO6),
.I1(CLBLM_L_X50Y107_SLICE_X76Y107_BQ),
.I2(CLBLM_L_X60Y96_SLICE_X90Y96_AQ),
.I3(CLBLM_L_X50Y107_SLICE_X77Y107_AQ),
.I4(CLBLM_L_X60Y96_SLICE_X90Y96_BQ),
.I5(1'b1),
.O5(CLBLM_R_X59Y96_SLICE_X89Y96_AO5),
.O6(CLBLM_R_X59Y96_SLICE_X89Y96_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y97_SLICE_X88Y97_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y97_SLICE_X88Y97_AO6),
.Q(CLBLM_R_X59Y97_SLICE_X88Y97_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y97_SLICE_X88Y97_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y97_SLICE_X88Y97_BO6),
.Q(CLBLM_R_X59Y97_SLICE_X88Y97_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0802000f0d0705)
  ) CLBLM_R_X59Y97_SLICE_X88Y97_DLUT (
.I0(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I1(CLBLL_R_X57Y97_SLICE_X86Y97_CO6),
.I2(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I3(CLBLM_R_X59Y97_SLICE_X88Y97_BQ),
.I4(CLBLM_R_X59Y97_SLICE_X89Y97_DQ),
.I5(CLBLM_L_X60Y97_SLICE_X90Y97_BO6),
.O5(CLBLM_R_X59Y97_SLICE_X88Y97_DO5),
.O6(CLBLM_R_X59Y97_SLICE_X88Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5410555554100000)
  ) CLBLM_R_X59Y97_SLICE_X88Y97_CLUT (
.I0(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I1(CLBLL_R_X57Y97_SLICE_X86Y97_CO6),
.I2(CLBLM_R_X59Y97_SLICE_X88Y97_AQ),
.I3(CLBLM_R_X59Y97_SLICE_X89Y97_CQ),
.I4(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I5(CLBLM_L_X50Y106_SLICE_X76Y106_AQ),
.O5(CLBLM_R_X59Y97_SLICE_X88Y97_CO5),
.O6(CLBLM_R_X59Y97_SLICE_X88Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaeeaaaacccccccc)
  ) CLBLM_R_X59Y97_SLICE_X88Y97_BLUT (
.I0(CLBLM_R_X59Y97_SLICE_X88Y97_DO6),
.I1(CLBLM_R_X59Y97_SLICE_X88Y97_BQ),
.I2(CLBLM_R_X49Y105_SLICE_X75Y105_CQ),
.I3(CLBLM_L_X60Y99_SLICE_X91Y99_DO6),
.I4(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I5(CLBLL_R_X57Y98_SLICE_X86Y98_DO6),
.O5(CLBLM_R_X59Y97_SLICE_X88Y97_BO5),
.O6(CLBLM_R_X59Y97_SLICE_X88Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcfcfcec4c0c0c)
  ) CLBLM_R_X59Y97_SLICE_X88Y97_ALUT (
.I0(CLBLM_L_X60Y99_SLICE_X91Y99_DO6),
.I1(CLBLM_R_X59Y97_SLICE_X88Y97_AQ),
.I2(CLBLL_R_X57Y98_SLICE_X86Y98_BO6),
.I3(CLBLM_L_X50Y105_SLICE_X77Y105_AQ),
.I4(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I5(CLBLM_R_X59Y97_SLICE_X88Y97_CO6),
.O5(CLBLM_R_X59Y97_SLICE_X88Y97_AO5),
.O6(CLBLM_R_X59Y97_SLICE_X88Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y97_SLICE_X89Y97_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_R_X57Y97_SLICE_X87Y97_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y96_SLICE_X88Y96_BQ),
.Q(CLBLM_R_X59Y97_SLICE_X89Y97_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y97_SLICE_X89Y97_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_R_X57Y97_SLICE_X87Y97_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y96_SLICE_X88Y96_AQ),
.Q(CLBLM_R_X59Y97_SLICE_X89Y97_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y97_SLICE_X89Y97_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_R_X57Y97_SLICE_X87Y97_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y98_SLICE_X89Y98_BQ),
.Q(CLBLM_R_X59Y97_SLICE_X89Y97_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y97_SLICE_X89Y97_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_R_X57Y97_SLICE_X87Y97_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y98_SLICE_X89Y98_B5Q),
.Q(CLBLM_R_X59Y97_SLICE_X89Y97_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y97_SLICE_X89Y97_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_R_X57Y97_SLICE_X87Y97_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y97_SLICE_X89Y97_AO6),
.Q(CLBLM_R_X59Y97_SLICE_X89Y97_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y97_SLICE_X89Y97_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_R_X57Y97_SLICE_X87Y97_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y97_SLICE_X89Y97_BO6),
.Q(CLBLM_R_X59Y97_SLICE_X89Y97_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y97_SLICE_X89Y97_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_R_X57Y97_SLICE_X87Y97_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y97_SLICE_X89Y97_CO6),
.Q(CLBLM_R_X59Y97_SLICE_X89Y97_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y97_SLICE_X89Y97_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_R_X57Y97_SLICE_X87Y97_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y97_SLICE_X89Y97_DO6),
.Q(CLBLM_R_X59Y97_SLICE_X89Y97_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X59Y97_SLICE_X89Y97_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X59Y97_SLICE_X88Y97_BQ),
.O5(CLBLM_R_X59Y97_SLICE_X89Y97_DO5),
.O6(CLBLM_R_X59Y97_SLICE_X89Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X59Y97_SLICE_X89Y97_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X59Y97_SLICE_X88Y97_AQ),
.O5(CLBLM_R_X59Y97_SLICE_X89Y97_CO5),
.O6(CLBLM_R_X59Y97_SLICE_X89Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X59Y97_SLICE_X89Y97_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X59Y98_SLICE_X88Y98_AQ),
.O5(CLBLM_R_X59Y97_SLICE_X89Y97_BO5),
.O6(CLBLM_R_X59Y97_SLICE_X89Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X59Y97_SLICE_X89Y97_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X59Y98_SLICE_X88Y98_DQ),
.O5(CLBLM_R_X59Y97_SLICE_X89Y97_AO5),
.O6(CLBLM_R_X59Y97_SLICE_X89Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y98_SLICE_X88Y98_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_R_X57Y101_SLICE_X86Y101_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y98_SLICE_X88Y98_AO6),
.Q(CLBLM_R_X59Y98_SLICE_X88Y98_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y98_SLICE_X88Y98_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_R_X57Y101_SLICE_X86Y101_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y98_SLICE_X88Y98_BO6),
.Q(CLBLM_R_X59Y98_SLICE_X88Y98_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y98_SLICE_X88Y98_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_R_X57Y101_SLICE_X86Y101_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y98_SLICE_X88Y98_CO6),
.Q(CLBLM_R_X59Y98_SLICE_X88Y98_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y98_SLICE_X88Y98_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_R_X57Y101_SLICE_X86Y101_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y98_SLICE_X88Y98_DO6),
.Q(CLBLM_R_X59Y98_SLICE_X88Y98_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfb08f80ff00ff00)
  ) CLBLM_R_X59Y98_SLICE_X88Y98_DLUT (
.I0(CLBLM_L_X50Y104_SLICE_X76Y104_AQ),
.I1(CLBLM_L_X60Y99_SLICE_X91Y99_AO5),
.I2(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I3(CLBLM_L_X62Y100_SLICE_X92Y100_AQ),
.I4(CLBLM_R_X59Y97_SLICE_X89Y97_AQ),
.I5(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.O5(CLBLM_R_X59Y98_SLICE_X88Y98_DO5),
.O6(CLBLM_R_X59Y98_SLICE_X88Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5dda088ffff0000)
  ) CLBLM_R_X59Y98_SLICE_X88Y98_CLUT (
.I0(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I1(CLBLM_R_X59Y100_SLICE_X88Y100_CQ),
.I2(CLBLM_L_X50Y106_SLICE_X76Y106_AQ),
.I3(CLBLM_L_X60Y99_SLICE_X91Y99_AO5),
.I4(CLBLM_L_X64Y100_SLICE_X97Y100_AQ),
.I5(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.O5(CLBLM_R_X59Y98_SLICE_X88Y98_CO5),
.O6(CLBLM_R_X59Y98_SLICE_X88Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heecce4cc4ecc44cc)
  ) CLBLM_R_X59Y98_SLICE_X88Y98_BLUT (
.I0(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I1(CLBLM_L_X62Y101_SLICE_X93Y101_AQ),
.I2(CLBLM_L_X60Y99_SLICE_X91Y99_AO5),
.I3(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I4(CLBLM_R_X59Y100_SLICE_X88Y100_AQ),
.I5(CLBLM_R_X49Y105_SLICE_X75Y105_CQ),
.O5(CLBLM_R_X59Y98_SLICE_X88Y98_BO5),
.O6(CLBLM_R_X59Y98_SLICE_X88Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafcccccca0cccccc)
  ) CLBLM_R_X59Y98_SLICE_X88Y98_ALUT (
.I0(CLBLM_L_X50Y105_SLICE_X77Y105_AQ),
.I1(CLBLM_L_X62Y100_SLICE_X92Y100_BQ),
.I2(CLBLM_L_X60Y99_SLICE_X91Y99_AO5),
.I3(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I4(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I5(CLBLM_R_X59Y97_SLICE_X89Y97_BQ),
.O5(CLBLM_R_X59Y98_SLICE_X88Y98_AO5),
.O6(CLBLM_R_X59Y98_SLICE_X88Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y98_SLICE_X89Y98_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_R_X59Y98_SLICE_X89Y98_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y98_SLICE_X89Y98_AO5),
.Q(CLBLM_R_X59Y98_SLICE_X89Y98_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y98_SLICE_X89Y98_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_R_X59Y98_SLICE_X89Y98_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y98_SLICE_X89Y98_BO5),
.Q(CLBLM_R_X59Y98_SLICE_X89Y98_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y98_SLICE_X89Y98_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_R_X59Y98_SLICE_X89Y98_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y98_SLICE_X89Y98_CO5),
.Q(CLBLM_R_X59Y98_SLICE_X89Y98_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y98_SLICE_X89Y98_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_R_X59Y98_SLICE_X89Y98_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y98_SLICE_X89Y98_AO6),
.Q(CLBLM_R_X59Y98_SLICE_X89Y98_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y98_SLICE_X89Y98_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_R_X59Y98_SLICE_X89Y98_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y98_SLICE_X89Y98_BO6),
.Q(CLBLM_R_X59Y98_SLICE_X89Y98_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y98_SLICE_X89Y98_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_R_X59Y98_SLICE_X89Y98_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y98_SLICE_X89Y98_CO6),
.Q(CLBLM_R_X59Y98_SLICE_X89Y98_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0000000f0a00000)
  ) CLBLM_R_X59Y98_SLICE_X89Y98_DLUT (
.I0(CLBLM_L_X56Y98_SLICE_X85Y98_BQ),
.I1(1'b1),
.I2(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.I3(CLBLM_L_X60Y98_SLICE_X90Y98_DO6),
.I4(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I5(CLBLM_L_X56Y98_SLICE_X85Y98_CQ),
.O5(CLBLM_R_X59Y98_SLICE_X89Y98_DO5),
.O6(CLBLM_R_X59Y98_SLICE_X89Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc00ccaaf0aaf0)
  ) CLBLM_R_X59Y98_SLICE_X89Y98_CLUT (
.I0(CLBLM_L_X50Y106_SLICE_X76Y106_CQ),
.I1(CLBLL_R_X57Y98_SLICE_X87Y98_CQ),
.I2(CLBLL_R_X57Y98_SLICE_X87Y98_DQ),
.I3(CLBLM_L_X60Y98_SLICE_X90Y98_DO6),
.I4(CLBLM_L_X50Y106_SLICE_X76Y106_AQ),
.I5(1'b1),
.O5(CLBLM_R_X59Y98_SLICE_X89Y98_CO5),
.O6(CLBLM_R_X59Y98_SLICE_X89Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88fafa5050)
  ) CLBLM_R_X59Y98_SLICE_X89Y98_BLUT (
.I0(CLBLM_L_X60Y98_SLICE_X90Y98_DO6),
.I1(CLBLM_R_X49Y105_SLICE_X75Y105_CQ),
.I2(CLBLM_R_X59Y97_SLICE_X89Y97_D5Q),
.I3(CLBLM_R_X59Y97_SLICE_X89Y97_C5Q),
.I4(CLBLM_R_X49Y106_SLICE_X74Y106_AQ),
.I5(1'b1),
.O5(CLBLM_R_X59Y98_SLICE_X89Y98_BO5),
.O6(CLBLM_R_X59Y98_SLICE_X89Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8d8d8ffaa5500)
  ) CLBLM_R_X59Y98_SLICE_X89Y98_ALUT (
.I0(CLBLM_L_X60Y98_SLICE_X90Y98_DO6),
.I1(CLBLM_L_X50Y104_SLICE_X76Y104_AQ),
.I2(CLBLL_R_X57Y98_SLICE_X87Y98_AQ),
.I3(CLBLL_R_X57Y98_SLICE_X87Y98_BQ),
.I4(CLBLM_L_X50Y105_SLICE_X77Y105_AQ),
.I5(1'b1),
.O5(CLBLM_R_X59Y98_SLICE_X89Y98_AO5),
.O6(CLBLM_R_X59Y98_SLICE_X89Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X59Y99_SLICE_X88Y99_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_R_X57Y99_SLICE_X87Y99_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y99_SLICE_X88Y99_BO5),
.Q(CLBLM_R_X59Y99_SLICE_X88Y99_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X59Y99_SLICE_X88Y99_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_R_X57Y99_SLICE_X87Y99_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y99_SLICE_X88Y99_AO6),
.Q(CLBLM_R_X59Y99_SLICE_X88Y99_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X59Y99_SLICE_X88Y99_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_R_X57Y99_SLICE_X87Y99_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y99_SLICE_X88Y99_BO6),
.Q(CLBLM_R_X59Y99_SLICE_X88Y99_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X59Y99_SLICE_X88Y99_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_R_X57Y99_SLICE_X87Y99_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y99_SLICE_X88Y99_CO6),
.Q(CLBLM_R_X59Y99_SLICE_X88Y99_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X59Y99_SLICE_X88Y99_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_R_X57Y99_SLICE_X87Y99_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y99_SLICE_X88Y99_DO6),
.Q(CLBLM_R_X59Y99_SLICE_X88Y99_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc00ccf0ccf0cc)
  ) CLBLM_R_X59Y99_SLICE_X88Y99_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X49Y107_SLICE_X75Y107_DQ),
.I2(CLBLM_R_X49Y107_SLICE_X75Y107_CQ),
.I3(CLBLM_L_X56Y99_SLICE_X84Y99_BQ),
.I4(CLBLM_R_X59Y98_SLICE_X88Y98_AQ),
.I5(CLBLM_L_X56Y99_SLICE_X84Y99_AQ),
.O5(CLBLM_R_X59Y99_SLICE_X88Y99_DO5),
.O6(CLBLM_R_X59Y99_SLICE_X88Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88bb88ffcc3300)
  ) CLBLM_R_X59Y99_SLICE_X88Y99_CLUT (
.I0(CLBLM_R_X59Y98_SLICE_X88Y98_DQ),
.I1(CLBLM_L_X56Y99_SLICE_X84Y99_BQ),
.I2(1'b1),
.I3(CLBLM_R_X49Y108_SLICE_X75Y108_DQ),
.I4(CLBLM_R_X49Y107_SLICE_X75Y107_CQ),
.I5(CLBLM_L_X56Y99_SLICE_X84Y99_AQ),
.O5(CLBLM_R_X59Y99_SLICE_X88Y99_CO5),
.O6(CLBLM_R_X59Y99_SLICE_X88Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaccaaccaa)
  ) CLBLM_R_X59Y99_SLICE_X88Y99_BLUT (
.I0(CLBLM_R_X49Y107_SLICE_X75Y107_CQ),
.I1(CLBLM_R_X59Y100_SLICE_X89Y100_BQ),
.I2(CLBLM_R_X59Y98_SLICE_X88Y98_CQ),
.I3(CLBLM_L_X56Y99_SLICE_X84Y99_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y99_SLICE_X88Y99_BO5),
.O6(CLBLM_R_X59Y99_SLICE_X88Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ee22f0f0f0f0)
  ) CLBLM_R_X59Y99_SLICE_X88Y99_ALUT (
.I0(CLBLM_R_X49Y107_SLICE_X75Y107_CQ),
.I1(CLBLM_L_X56Y99_SLICE_X84Y99_AQ),
.I2(CLBLM_R_X49Y108_SLICE_X75Y108_BQ),
.I3(CLBLM_R_X59Y100_SLICE_X89Y100_AQ),
.I4(1'b1),
.I5(CLBLM_L_X56Y99_SLICE_X84Y99_BQ),
.O5(CLBLM_R_X59Y99_SLICE_X88Y99_AO5),
.O6(CLBLM_R_X59Y99_SLICE_X88Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X59Y99_SLICE_X89Y99_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_R_X57Y99_SLICE_X87Y99_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y99_SLICE_X89Y99_AO5),
.Q(CLBLM_R_X59Y99_SLICE_X89Y99_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X59Y99_SLICE_X89Y99_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_R_X57Y99_SLICE_X87Y99_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y99_SLICE_X89Y99_AO6),
.Q(CLBLM_R_X59Y99_SLICE_X89Y99_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X59Y99_SLICE_X89Y99_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_R_X57Y99_SLICE_X87Y99_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y99_SLICE_X89Y99_BO6),
.Q(CLBLM_R_X59Y99_SLICE_X89Y99_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X59Y99_SLICE_X89Y99_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y99_SLICE_X89Y99_DO5),
.O6(CLBLM_R_X59Y99_SLICE_X89Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h020a020a02020202)
  ) CLBLM_R_X59Y99_SLICE_X89Y99_CLUT (
.I0(CLBLM_L_X62Y99_SLICE_X92Y99_AO6),
.I1(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I2(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I3(CLBLM_L_X56Y99_SLICE_X84Y99_BQ),
.I4(1'b1),
.I5(CLBLM_L_X56Y99_SLICE_X84Y99_AQ),
.O5(CLBLM_R_X59Y99_SLICE_X89Y99_CO5),
.O6(CLBLM_R_X59Y99_SLICE_X89Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000cccccccc)
  ) CLBLM_R_X59Y99_SLICE_X89Y99_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X49Y108_SLICE_X75Y108_AQ),
.I2(CLBLM_R_X59Y98_SLICE_X88Y98_BQ),
.I3(CLBLM_L_X56Y99_SLICE_X84Y99_AQ),
.I4(CLBLM_R_X49Y107_SLICE_X75Y107_CQ),
.I5(CLBLM_L_X56Y99_SLICE_X84Y99_BQ),
.O5(CLBLM_R_X59Y99_SLICE_X89Y99_BO5),
.O6(CLBLM_R_X59Y99_SLICE_X89Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00f0fff000)
  ) CLBLM_R_X59Y99_SLICE_X89Y99_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X59Y100_SLICE_X89Y100_CQ),
.I2(CLBLM_R_X59Y100_SLICE_X89Y100_DQ),
.I3(CLBLM_L_X56Y99_SLICE_X84Y99_AQ),
.I4(CLBLM_R_X49Y107_SLICE_X75Y107_CQ),
.I5(1'b1),
.O5(CLBLM_R_X59Y99_SLICE_X89Y99_AO5),
.O6(CLBLM_R_X59Y99_SLICE_X89Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y100_SLICE_X88Y100_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLL_R_X57Y97_SLICE_X87Y97_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y100_SLICE_X89Y100_CQ),
.Q(CLBLM_R_X59Y100_SLICE_X88Y100_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y100_SLICE_X88Y100_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLL_R_X57Y97_SLICE_X87Y97_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y100_SLICE_X89Y100_DQ),
.Q(CLBLM_R_X59Y100_SLICE_X88Y100_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y100_SLICE_X88Y100_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLL_R_X57Y97_SLICE_X87Y97_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y98_SLICE_X88Y98_BQ),
.Q(CLBLM_R_X59Y100_SLICE_X88Y100_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y100_SLICE_X88Y100_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLL_R_X57Y97_SLICE_X87Y97_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y100_SLICE_X88Y100_BO6),
.Q(CLBLM_R_X59Y100_SLICE_X88Y100_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y100_SLICE_X88Y100_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLL_R_X57Y97_SLICE_X87Y97_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y100_SLICE_X88Y100_CO6),
.Q(CLBLM_R_X59Y100_SLICE_X88Y100_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y100_SLICE_X88Y100_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLL_R_X57Y97_SLICE_X87Y97_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y100_SLICE_X89Y100_BQ),
.Q(CLBLM_R_X59Y100_SLICE_X88Y100_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffdf0000ffff0000)
  ) CLBLM_R_X59Y100_SLICE_X88Y100_DLUT (
.I0(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I1(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I2(CLBLL_L_X54Y101_SLICE_X83Y101_AO6),
.I3(CLBLM_L_X64Y100_SLICE_X97Y100_BQ),
.I4(CLBLM_R_X59Y101_SLICE_X88Y101_CO6),
.I5(CLBLM_L_X64Y100_SLICE_X97Y100_AQ),
.O5(CLBLM_R_X59Y100_SLICE_X88Y100_DO5),
.O6(CLBLM_R_X59Y100_SLICE_X88Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X59Y100_SLICE_X88Y100_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X59Y98_SLICE_X88Y98_CQ),
.O5(CLBLM_R_X59Y100_SLICE_X88Y100_CO5),
.O6(CLBLM_R_X59Y100_SLICE_X88Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X59Y100_SLICE_X88Y100_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X59Y100_SLICE_X89Y100_AQ),
.O5(CLBLM_R_X59Y100_SLICE_X88Y100_BO5),
.O6(CLBLM_R_X59Y100_SLICE_X88Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h05050505f353a303)
  ) CLBLM_R_X59Y100_SLICE_X88Y100_ALUT (
.I0(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I1(CLBLM_L_X60Y100_SLICE_X90Y100_AQ),
.I2(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I3(CLBLM_L_X50Y104_SLICE_X76Y104_AQ),
.I4(CLBLM_R_X49Y104_SLICE_X74Y104_AQ),
.I5(1'b1),
.O5(CLBLM_R_X59Y100_SLICE_X88Y100_AO5),
.O6(CLBLM_R_X59Y100_SLICE_X88Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y100_SLICE_X89Y100_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLL_R_X57Y101_SLICE_X86Y101_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y100_SLICE_X89Y100_AO6),
.Q(CLBLM_R_X59Y100_SLICE_X89Y100_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y100_SLICE_X89Y100_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLL_R_X57Y101_SLICE_X86Y101_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y100_SLICE_X89Y100_BO6),
.Q(CLBLM_R_X59Y100_SLICE_X89Y100_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y100_SLICE_X89Y100_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLL_R_X57Y101_SLICE_X86Y101_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y100_SLICE_X89Y100_CO6),
.Q(CLBLM_R_X59Y100_SLICE_X89Y100_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y100_SLICE_X89Y100_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLL_R_X57Y101_SLICE_X86Y101_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y100_SLICE_X89Y100_DO6),
.Q(CLBLM_R_X59Y100_SLICE_X89Y100_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7a2d580ff00ff00)
  ) CLBLM_R_X59Y100_SLICE_X89Y100_DLUT (
.I0(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I1(CLBLM_L_X60Y99_SLICE_X91Y99_AO5),
.I2(CLBLM_L_X50Y107_SLICE_X77Y107_AQ),
.I3(CLBLM_L_X62Y101_SLICE_X93Y101_CQ),
.I4(CLBLM_R_X59Y100_SLICE_X88Y100_C5Q),
.I5(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.O5(CLBLM_R_X59Y100_SLICE_X89Y100_DO5),
.O6(CLBLM_R_X59Y100_SLICE_X89Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfda8ff007520ff00)
  ) CLBLM_R_X59Y100_SLICE_X89Y100_CLUT (
.I0(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I1(CLBLM_L_X60Y99_SLICE_X91Y99_AO5),
.I2(CLBLM_R_X59Y100_SLICE_X88Y100_B5Q),
.I3(CLBLM_L_X62Y101_SLICE_X93Y101_BQ),
.I4(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I5(CLBLM_L_X50Y107_SLICE_X76Y107_BQ),
.O5(CLBLM_R_X59Y100_SLICE_X89Y100_CO5),
.O6(CLBLM_R_X59Y100_SLICE_X89Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7d5ffffa2800000)
  ) CLBLM_R_X59Y100_SLICE_X89Y100_BLUT (
.I0(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I1(CLBLM_L_X60Y99_SLICE_X91Y99_AO5),
.I2(CLBLM_L_X50Y106_SLICE_X76Y106_CQ),
.I3(CLBLM_R_X59Y100_SLICE_X88Y100_DQ),
.I4(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I5(CLBLM_L_X64Y100_SLICE_X97Y100_BQ),
.O5(CLBLM_R_X59Y100_SLICE_X89Y100_BO5),
.O6(CLBLM_R_X59Y100_SLICE_X89Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7d5ffffa2800000)
  ) CLBLM_R_X59Y100_SLICE_X89Y100_ALUT (
.I0(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I1(CLBLM_L_X60Y99_SLICE_X91Y99_AO5),
.I2(CLBLM_R_X49Y106_SLICE_X74Y106_AQ),
.I3(CLBLM_R_X59Y100_SLICE_X88Y100_BQ),
.I4(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I5(CLBLM_L_X62Y100_SLICE_X92Y100_CQ),
.O5(CLBLM_R_X59Y100_SLICE_X89Y100_AO5),
.O6(CLBLM_R_X59Y100_SLICE_X89Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h03034477cfcf4477)
  ) CLBLM_R_X59Y101_SLICE_X88Y101_DLUT (
.I0(CLBLM_R_X59Y111_SLICE_X89Y111_AQ),
.I1(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I2(CLBLM_R_X59Y106_SLICE_X89Y106_CQ),
.I3(CLBLM_R_X59Y98_SLICE_X89Y98_A5Q),
.I4(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I5(CLBLM_R_X59Y98_SLICE_X88Y98_AQ),
.O5(CLBLM_R_X59Y101_SLICE_X88Y101_DO5),
.O6(CLBLM_R_X59Y101_SLICE_X88Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff7ffcfffff)
  ) CLBLM_R_X59Y101_SLICE_X88Y101_CLUT (
.I0(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I1(CLBLM_R_X59Y103_SLICE_X89Y103_CQ),
.I2(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I3(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I4(CLBLM_R_X59Y103_SLICE_X89Y103_DQ),
.I5(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.O5(CLBLM_R_X59Y101_SLICE_X88Y101_CO5),
.O6(CLBLM_R_X59Y101_SLICE_X88Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000202000100)
  ) CLBLM_R_X59Y101_SLICE_X88Y101_BLUT (
.I0(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I1(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I2(CLBLM_R_X59Y103_SLICE_X89Y103_DQ),
.I3(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I4(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I5(CLBLM_R_X59Y103_SLICE_X89Y103_CQ),
.O5(CLBLM_R_X59Y101_SLICE_X88Y101_BO5),
.O6(CLBLM_R_X59Y101_SLICE_X88Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00fb00ff00ff)
  ) CLBLM_R_X59Y101_SLICE_X88Y101_ALUT (
.I0(CLBLM_L_X64Y100_SLICE_X97Y100_AQ),
.I1(CLBLL_L_X54Y101_SLICE_X83Y101_AO6),
.I2(CLBLM_L_X64Y100_SLICE_X97Y100_BQ),
.I3(CLBLM_R_X59Y101_SLICE_X88Y101_BO6),
.I4(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I5(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.O5(CLBLM_R_X59Y101_SLICE_X88Y101_AO5),
.O6(CLBLM_R_X59Y101_SLICE_X88Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X59Y101_SLICE_X89Y101_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y101_SLICE_X89Y101_AO6),
.Q(CLBLM_R_X59Y101_SLICE_X89Y101_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h555533330f0f00ff)
  ) CLBLM_R_X59Y101_SLICE_X89Y101_DLUT (
.I0(CLBLM_R_X59Y100_SLICE_X89Y100_AQ),
.I1(CLBLM_R_X59Y110_SLICE_X89Y110_AQ),
.I2(CLBLM_R_X59Y104_SLICE_X89Y104_CQ),
.I3(CLBLM_R_X59Y98_SLICE_X89Y98_B5Q),
.I4(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I5(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.O5(CLBLM_R_X59Y101_SLICE_X89Y101_DO5),
.O6(CLBLM_R_X59Y101_SLICE_X89Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h535300f053530fff)
  ) CLBLM_R_X59Y101_SLICE_X89Y101_CLUT (
.I0(CLBLM_R_X59Y98_SLICE_X88Y98_BQ),
.I1(CLBLM_R_X59Y111_SLICE_X89Y111_BQ),
.I2(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I3(CLBLM_R_X59Y105_SLICE_X89Y105_CQ),
.I4(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I5(CLBLM_R_X59Y98_SLICE_X89Y98_BQ),
.O5(CLBLM_R_X59Y101_SLICE_X89Y101_CO5),
.O6(CLBLM_R_X59Y101_SLICE_X89Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfff6ffffffffff)
  ) CLBLM_R_X59Y101_SLICE_X89Y101_BLUT (
.I0(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I1(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I2(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I3(CLBLM_R_X59Y103_SLICE_X89Y103_DQ),
.I4(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I5(CLBLM_R_X59Y103_SLICE_X89Y103_CQ),
.O5(CLBLM_R_X59Y101_SLICE_X89Y101_BO5),
.O6(CLBLM_R_X59Y101_SLICE_X89Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000001000)
  ) CLBLM_R_X59Y101_SLICE_X89Y101_ALUT (
.I0(CLBLM_R_X49Y107_SLICE_X75Y107_CQ),
.I1(CLBLM_R_X49Y106_SLICE_X75Y106_DQ),
.I2(CLBLM_L_X56Y102_SLICE_X85Y102_BO6),
.I3(CLBLM_R_X49Y104_SLICE_X75Y104_CQ),
.I4(CLBLM_R_X49Y106_SLICE_X75Y106_CQ),
.I5(CLBLM_R_X49Y104_SLICE_X75Y104_DQ),
.O5(CLBLM_R_X59Y101_SLICE_X89Y101_AO5),
.O6(CLBLM_R_X59Y101_SLICE_X89Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X59Y102_SLICE_X88Y102_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_R_X59Y99_SLICE_X89Y99_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y102_SLICE_X88Y102_AO6),
.Q(CLBLM_R_X59Y102_SLICE_X88Y102_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff330033f055f055)
  ) CLBLM_R_X59Y102_SLICE_X88Y102_DLUT (
.I0(CLBLM_R_X59Y101_SLICE_X88Y101_DO6),
.I1(CLBLM_R_X59Y102_SLICE_X89Y102_CO6),
.I2(CLBLM_R_X63Y103_SLICE_X94Y103_AO6),
.I3(CLBLM_L_X62Y103_SLICE_X93Y103_BO6),
.I4(CLBLL_R_X57Y105_SLICE_X86Y105_CO6),
.I5(CLBLM_L_X62Y106_SLICE_X93Y106_CO6),
.O5(CLBLM_R_X59Y102_SLICE_X88Y102_DO5),
.O6(CLBLM_R_X59Y102_SLICE_X88Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h555500ff0f0f3333)
  ) CLBLM_R_X59Y102_SLICE_X88Y102_CLUT (
.I0(CLBLM_R_X63Y100_SLICE_X94Y100_AQ),
.I1(CLBLM_L_X60Y101_SLICE_X90Y101_AQ),
.I2(CLBLL_R_X57Y97_SLICE_X86Y97_AQ),
.I3(CLBLM_L_X62Y102_SLICE_X92Y102_BQ),
.I4(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I5(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.O5(CLBLM_R_X59Y102_SLICE_X88Y102_CO5),
.O6(CLBLM_R_X59Y102_SLICE_X88Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h333333333535c0cf)
  ) CLBLM_R_X59Y102_SLICE_X88Y102_BLUT (
.I0(CLBLL_R_X57Y109_SLICE_X87Y109_A_XOR),
.I1(CLBLL_R_X57Y101_SLICE_X86Y101_AQ),
.I2(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I3(CLBLM_R_X59Y103_SLICE_X88Y103_BQ),
.I4(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I5(CLBLM_R_X59Y103_SLICE_X89Y103_CQ),
.O5(CLBLM_R_X59Y102_SLICE_X88Y102_BO5),
.O6(CLBLM_R_X59Y102_SLICE_X88Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfcfcfc0c0c0c5)
  ) CLBLM_R_X59Y102_SLICE_X88Y102_ALUT (
.I0(CLBLM_R_X59Y103_SLICE_X89Y103_DQ),
.I1(CLBLM_R_X49Y104_SLICE_X74Y104_AQ),
.I2(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I3(CLBLM_R_X59Y102_SLICE_X88Y102_BO6),
.I4(CLBLM_L_X62Y106_SLICE_X92Y106_AO5),
.I5(CLBLM_R_X59Y103_SLICE_X88Y103_F7AMUX_O),
.O5(CLBLM_R_X59Y102_SLICE_X88Y102_AO5),
.O6(CLBLM_R_X59Y102_SLICE_X88Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X59Y102_SLICE_X89Y102_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_R_X59Y99_SLICE_X89Y99_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y102_SLICE_X89Y102_AO6),
.Q(CLBLM_R_X59Y102_SLICE_X89Y102_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ff550f000fff)
  ) CLBLM_R_X59Y102_SLICE_X89Y102_DLUT (
.I0(CLBLM_L_X60Y102_SLICE_X90Y102_AQ),
.I1(1'b1),
.I2(CLBLM_R_X59Y96_SLICE_X88Y96_BQ),
.I3(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I4(CLBLM_L_X60Y109_SLICE_X91Y109_BQ),
.I5(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.O5(CLBLM_R_X59Y102_SLICE_X89Y102_DO5),
.O6(CLBLM_R_X59Y102_SLICE_X89Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ffff53535353)
  ) CLBLM_R_X59Y102_SLICE_X89Y102_CLUT (
.I0(CLBLM_R_X59Y97_SLICE_X88Y97_AQ),
.I1(CLBLM_L_X60Y109_SLICE_X91Y109_AQ),
.I2(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I3(1'b1),
.I4(CLBLM_L_X60Y102_SLICE_X90Y102_CQ),
.I5(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.O5(CLBLM_R_X59Y102_SLICE_X89Y102_CO5),
.O6(CLBLM_R_X59Y102_SLICE_X89Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h505003f35f5f03f3)
  ) CLBLM_R_X59Y102_SLICE_X89Y102_BLUT (
.I0(CLBLL_R_X57Y105_SLICE_X86Y105_DO6),
.I1(CLBLM_R_X59Y101_SLICE_X89Y101_DO6),
.I2(CLBLM_L_X62Y106_SLICE_X93Y106_CO6),
.I3(CLBLM_R_X59Y102_SLICE_X89Y102_DO6),
.I4(CLBLM_L_X62Y103_SLICE_X93Y103_BO6),
.I5(CLBLM_L_X62Y107_SLICE_X93Y107_CO6),
.O5(CLBLM_R_X59Y102_SLICE_X89Y102_BO5),
.O6(CLBLM_R_X59Y102_SLICE_X89Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfaccfacc50cc50)
  ) CLBLM_R_X59Y102_SLICE_X89Y102_ALUT (
.I0(CLBLM_R_X59Y103_SLICE_X89Y103_DQ),
.I1(CLBLM_R_X49Y104_SLICE_X75Y104_CQ),
.I2(CLBLM_R_X59Y106_SLICE_X89Y106_DO6),
.I3(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I4(1'b1),
.I5(CLBLM_L_X60Y102_SLICE_X90Y102_DO6),
.O5(CLBLM_R_X59Y102_SLICE_X89Y102_AO5),
.O6(CLBLM_R_X59Y102_SLICE_X89Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X59Y103_SLICE_X88Y103_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLL_R_X57Y99_SLICE_X87Y99_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y104_SLICE_X74Y104_AQ),
.Q(CLBLM_R_X59Y103_SLICE_X88Y103_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X59Y103_SLICE_X88Y103_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLL_R_X57Y99_SLICE_X87Y99_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y104_SLICE_X75Y104_AQ),
.Q(CLBLM_R_X59Y103_SLICE_X88Y103_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X59Y103_SLICE_X88Y103_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLL_R_X57Y99_SLICE_X87Y99_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y104_SLICE_X75Y104_BQ),
.Q(CLBLM_R_X59Y103_SLICE_X88Y103_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h110cdd0c113fdd3f)
  ) CLBLM_R_X59Y103_SLICE_X88Y103_DLUT (
.I0(CLBLM_L_X60Y100_SLICE_X90Y100_AQ),
.I1(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I2(CLBLM_R_X59Y111_SLICE_X89Y111_CQ),
.I3(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I4(CLBLM_R_X59Y98_SLICE_X88Y98_DQ),
.I5(CLBLM_R_X59Y98_SLICE_X89Y98_AQ),
.O5(CLBLM_R_X59Y103_SLICE_X88Y103_DO5),
.O6(CLBLM_R_X59Y103_SLICE_X88Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a5f0a5f22227777)
  ) CLBLM_R_X59Y103_SLICE_X88Y103_CLUT (
.I0(CLBLM_L_X62Y106_SLICE_X93Y106_CO6),
.I1(CLBLM_R_X59Y102_SLICE_X88Y102_CO6),
.I2(CLBLL_R_X57Y104_SLICE_X86Y104_DO6),
.I3(CLBLM_R_X59Y104_SLICE_X88Y104_DO6),
.I4(CLBLM_R_X59Y103_SLICE_X88Y103_DO6),
.I5(CLBLM_L_X62Y103_SLICE_X93Y103_BO6),
.O5(CLBLM_R_X59Y103_SLICE_X88Y103_CO5),
.O6(CLBLM_R_X59Y103_SLICE_X88Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f00aa0000000000)
  ) CLBLM_R_X59Y103_SLICE_X88Y103_BLUT (
.I0(CLBLM_R_X59Y108_SLICE_X88Y108_A_XOR),
.I1(1'b1),
.I2(CLBLM_L_X60Y100_SLICE_X90Y100_AQ),
.I3(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I4(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I5(CLBLM_R_X59Y103_SLICE_X89Y103_CQ),
.O5(CLBLM_R_X59Y103_SLICE_X88Y103_BO5),
.O6(CLBLM_R_X59Y103_SLICE_X88Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccc33aaf0f0f0)
  ) CLBLM_R_X59Y103_SLICE_X88Y103_ALUT (
.I0(CLBLM_L_X60Y105_SLICE_X90Y105_A_XOR),
.I1(CLBLM_L_X62Y102_SLICE_X92Y102_BQ),
.I2(CLBLM_L_X60Y100_SLICE_X90Y100_AQ),
.I3(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I4(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I5(CLBLM_R_X59Y103_SLICE_X89Y103_CQ),
.O5(CLBLM_R_X59Y103_SLICE_X88Y103_AO5),
.O6(CLBLM_R_X59Y103_SLICE_X88Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X59Y103_SLICE_X88Y103_MUXF7A (
.I0(CLBLM_R_X59Y103_SLICE_X88Y103_BO6),
.I1(CLBLM_R_X59Y103_SLICE_X88Y103_AO6),
.O(CLBLM_R_X59Y103_SLICE_X88Y103_F7AMUX_O),
.S(CLBLM_R_X59Y103_SLICE_X89Y103_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X59Y103_SLICE_X89Y103_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLL_R_X57Y102_SLICE_X86Y102_AO5),
.Q(CLBLM_R_X59Y103_SLICE_X89Y103_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X59Y103_SLICE_X89Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y103_SLICE_X89Y103_AO6),
.Q(CLBLM_R_X59Y103_SLICE_X89Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X59Y103_SLICE_X89Y103_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y103_SLICE_X89Y103_BO6),
.Q(CLBLM_R_X59Y103_SLICE_X89Y103_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X59Y103_SLICE_X89Y103_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y103_SLICE_X89Y103_CO6),
.Q(CLBLM_R_X59Y103_SLICE_X89Y103_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X59Y103_SLICE_X89Y103_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y103_SLICE_X89Y103_DO6),
.Q(CLBLM_R_X59Y103_SLICE_X89Y103_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777550077550000)
  ) CLBLM_R_X59Y103_SLICE_X89Y103_DLUT (
.I0(CLBLM_R_X59Y104_SLICE_X88Y104_AO6),
.I1(CLBLM_R_X59Y104_SLICE_X88Y104_AO5),
.I2(1'b1),
.I3(CLBLM_R_X59Y103_SLICE_X88Y103_CQ),
.I4(CLBLM_R_X59Y103_SLICE_X88Y103_DQ),
.I5(CLBLM_R_X59Y103_SLICE_X88Y103_BQ),
.O5(CLBLM_R_X59Y103_SLICE_X89Y103_DO5),
.O6(CLBLM_R_X59Y103_SLICE_X89Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4f5533005f770000)
  ) CLBLM_R_X59Y103_SLICE_X89Y103_CLUT (
.I0(CLBLM_R_X59Y104_SLICE_X88Y104_AO6),
.I1(CLBLM_R_X59Y104_SLICE_X88Y104_AO5),
.I2(CLBLM_R_X59Y104_SLICE_X89Y104_DO6),
.I3(CLBLM_R_X59Y103_SLICE_X88Y103_CQ),
.I4(CLBLM_R_X59Y103_SLICE_X88Y103_DQ),
.I5(CLBLM_R_X59Y103_SLICE_X88Y103_BQ),
.O5(CLBLM_R_X59Y103_SLICE_X89Y103_CO5),
.O6(CLBLM_R_X59Y103_SLICE_X89Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c082222cc0822aa)
  ) CLBLM_R_X59Y103_SLICE_X89Y103_BLUT (
.I0(CLBLM_R_X59Y103_SLICE_X88Y103_DQ),
.I1(CLBLM_R_X59Y104_SLICE_X89Y104_DO6),
.I2(CLBLM_R_X59Y104_SLICE_X88Y104_AO6),
.I3(CLBLM_R_X59Y103_SLICE_X88Y103_BQ),
.I4(CLBLM_R_X59Y103_SLICE_X88Y103_CQ),
.I5(CLBLM_R_X59Y104_SLICE_X88Y104_AO5),
.O5(CLBLM_R_X59Y103_SLICE_X89Y103_BO5),
.O6(CLBLM_R_X59Y103_SLICE_X89Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3020f0a03a2afaaa)
  ) CLBLM_R_X59Y103_SLICE_X89Y103_ALUT (
.I0(CLBLM_R_X59Y103_SLICE_X88Y103_DQ),
.I1(CLBLM_R_X59Y104_SLICE_X89Y104_DO6),
.I2(CLBLM_R_X59Y103_SLICE_X88Y103_BQ),
.I3(CLBLM_R_X59Y103_SLICE_X88Y103_CQ),
.I4(CLBLM_R_X59Y104_SLICE_X88Y104_AO6),
.I5(CLBLM_R_X59Y104_SLICE_X88Y104_AO5),
.O5(CLBLM_R_X59Y103_SLICE_X89Y103_AO5),
.O6(CLBLM_R_X59Y103_SLICE_X89Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X59Y104_SLICE_X88Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLL_R_X57Y99_SLICE_X87Y99_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y104_SLICE_X75Y104_CQ),
.Q(CLBLM_R_X59Y104_SLICE_X88Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X59Y104_SLICE_X88Y104_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLL_R_X57Y99_SLICE_X87Y99_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y106_SLICE_X75Y106_CQ),
.Q(CLBLM_R_X59Y104_SLICE_X88Y104_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0f3300ff0f33ff)
  ) CLBLM_R_X59Y104_SLICE_X88Y104_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X62Y105_SLICE_X92Y105_CQ),
.I2(CLBLM_R_X49Y109_SLICE_X74Y109_DQ),
.I3(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I4(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I5(CLBLM_L_X64Y107_SLICE_X97Y107_BQ),
.O5(CLBLM_R_X59Y104_SLICE_X88Y104_DO5),
.O6(CLBLM_R_X59Y104_SLICE_X88Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5ffffffffffa)
  ) CLBLM_R_X59Y104_SLICE_X88Y104_CLUT (
.I0(CLBLM_R_X59Y99_SLICE_X88Y99_BQ),
.I1(1'b1),
.I2(CLBLM_R_X59Y99_SLICE_X89Y99_A5Q),
.I3(CLBLM_R_X59Y99_SLICE_X88Y99_B5Q),
.I4(CLBLM_R_X59Y106_SLICE_X88Y106_DO6),
.I5(CLBLM_R_X59Y99_SLICE_X89Y99_AQ),
.O5(CLBLM_R_X59Y104_SLICE_X88Y104_CO5),
.O6(CLBLM_R_X59Y104_SLICE_X88Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfffffffffffffef)
  ) CLBLM_R_X59Y104_SLICE_X88Y104_BLUT (
.I0(CLBLM_R_X59Y106_SLICE_X88Y106_DO6),
.I1(CLBLM_R_X59Y99_SLICE_X89Y99_AQ),
.I2(CLBLM_R_X59Y104_SLICE_X88Y104_AQ),
.I3(CLBLM_R_X59Y99_SLICE_X89Y99_A5Q),
.I4(CLBLM_R_X59Y99_SLICE_X88Y99_BQ),
.I5(CLBLM_R_X59Y99_SLICE_X88Y99_B5Q),
.O5(CLBLM_R_X59Y104_SLICE_X88Y104_BO5),
.O6(CLBLM_R_X59Y104_SLICE_X88Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffddffddfffffbfb)
  ) CLBLM_R_X59Y104_SLICE_X88Y104_ALUT (
.I0(CLBLM_R_X59Y107_SLICE_X89Y107_BQ),
.I1(CLBLM_R_X59Y104_SLICE_X88Y104_BQ),
.I2(CLBLM_R_X59Y104_SLICE_X88Y104_AQ),
.I3(CLBLM_R_X59Y104_SLICE_X88Y104_BO6),
.I4(CLBLM_R_X59Y104_SLICE_X88Y104_CO6),
.I5(1'b1),
.O5(CLBLM_R_X59Y104_SLICE_X88Y104_AO5),
.O6(CLBLM_R_X59Y104_SLICE_X88Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y104_SLICE_X89Y104_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y99_SLICE_X90Y99_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y104_SLICE_X89Y104_CO6),
.Q(CLBLM_R_X59Y104_SLICE_X89Y104_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcfcfcffffffff)
  ) CLBLM_R_X59Y104_SLICE_X89Y104_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X59Y107_SLICE_X89Y107_BQ),
.I2(CLBLM_R_X59Y104_SLICE_X88Y104_BO6),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X59Y104_SLICE_X88Y104_BQ),
.O5(CLBLM_R_X59Y104_SLICE_X89Y104_DO5),
.O6(CLBLM_R_X59Y104_SLICE_X89Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccefeeccccecee)
  ) CLBLM_R_X59Y104_SLICE_X89Y104_CLUT (
.I0(CLBLM_L_X60Y108_SLICE_X90Y108_C_XOR),
.I1(CLBLM_L_X62Y98_SLICE_X92Y98_AO6),
.I2(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I3(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I4(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I5(CLBLM_R_X59Y107_SLICE_X89Y107_C_XOR),
.O5(CLBLM_R_X59Y104_SLICE_X89Y104_CO5),
.O6(CLBLM_R_X59Y104_SLICE_X89Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33bb338800bb0088)
  ) CLBLM_R_X59Y104_SLICE_X89Y104_BLUT (
.I0(CLBLM_L_X64Y106_SLICE_X96Y106_BQ),
.I1(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I2(1'b1),
.I3(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I4(CLBLM_L_X64Y108_SLICE_X96Y108_BQ),
.I5(CLBLM_R_X49Y109_SLICE_X74Y109_CQ),
.O5(CLBLM_R_X59Y104_SLICE_X89Y104_BO5),
.O6(CLBLM_R_X59Y104_SLICE_X89Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7e6b3a2d5c49180)
  ) CLBLM_R_X59Y104_SLICE_X89Y104_ALUT (
.I0(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I1(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I2(CLBLM_R_X59Y106_SLICE_X88Y106_AQ),
.I3(CLBLL_R_X57Y104_SLICE_X87Y104_BQ),
.I4(CLBLM_L_X60Y107_SLICE_X90Y107_AQ),
.I5(CLBLM_L_X56Y104_SLICE_X85Y104_AQ),
.O5(CLBLM_R_X59Y104_SLICE_X89Y104_AO5),
.O6(CLBLM_R_X59Y104_SLICE_X89Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X59Y104_SLICE_X89Y104_MUXF7A (
.I0(CLBLM_R_X59Y104_SLICE_X89Y104_BO6),
.I1(CLBLM_R_X59Y104_SLICE_X89Y104_AO6),
.O(CLBLM_R_X59Y104_SLICE_X89Y104_F7AMUX_O),
.S(CLBLM_L_X62Y106_SLICE_X93Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y105_SLICE_X88Y105_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y100_SLICE_X90Y100_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y106_SLICE_X93Y106_BO6),
.Q(CLBLM_R_X59Y105_SLICE_X88Y105_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X59Y105_SLICE_X88Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y105_SLICE_X88Y105_DO5),
.O6(CLBLM_R_X59Y105_SLICE_X88Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcf6fffefcf7ffff)
  ) CLBLM_R_X59Y105_SLICE_X88Y105_CLUT (
.I0(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I1(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I2(CLBLM_R_X59Y103_SLICE_X89Y103_DQ),
.I3(CLBLM_R_X59Y103_SLICE_X89Y103_CQ),
.I4(CLBLM_R_X59Y105_SLICE_X88Y105_BQ),
.I5(CLBLM_R_X59Y99_SLICE_X88Y99_B5Q),
.O5(CLBLM_R_X59Y105_SLICE_X88Y105_CO5),
.O6(CLBLM_R_X59Y105_SLICE_X88Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha2f2a2f2a7f7a7f7)
  ) CLBLM_R_X59Y105_SLICE_X88Y105_BLUT (
.I0(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I1(CLBLM_R_X49Y109_SLICE_X74Y109_BQ),
.I2(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I3(CLBLM_L_X62Y105_SLICE_X93Y105_BQ),
.I4(1'b1),
.I5(CLBLM_L_X64Y108_SLICE_X97Y108_AQ),
.O5(CLBLM_R_X59Y105_SLICE_X88Y105_BO5),
.O6(CLBLM_R_X59Y105_SLICE_X88Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h05af222205af7777)
  ) CLBLM_R_X59Y105_SLICE_X88Y105_ALUT (
.I0(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I1(CLBLM_R_X59Y105_SLICE_X88Y105_BQ),
.I2(CLBLM_L_X56Y105_SLICE_X85Y105_BQ),
.I3(CLBLL_R_X57Y108_SLICE_X87Y108_AQ),
.I4(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I5(CLBLM_L_X56Y105_SLICE_X84Y105_BQ),
.O5(CLBLM_R_X59Y105_SLICE_X88Y105_AO5),
.O6(CLBLM_R_X59Y105_SLICE_X88Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X59Y105_SLICE_X88Y105_MUXF7A (
.I0(CLBLM_R_X59Y105_SLICE_X88Y105_BO6),
.I1(CLBLM_R_X59Y105_SLICE_X88Y105_AO6),
.O(CLBLM_R_X59Y105_SLICE_X88Y105_F7AMUX_O),
.S(CLBLM_L_X62Y106_SLICE_X93Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y105_SLICE_X89Y105_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y99_SLICE_X90Y99_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y105_SLICE_X89Y105_CO6),
.Q(CLBLM_R_X59Y105_SLICE_X89Y105_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55d8d8aa00d8d8)
  ) CLBLM_R_X59Y105_SLICE_X89Y105_DLUT (
.I0(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I1(CLBLM_R_X59Y108_SLICE_X89Y108_AQ),
.I2(CLBLM_R_X59Y96_SLICE_X89Y96_AQ),
.I3(CLBLM_R_X59Y100_SLICE_X89Y100_CQ),
.I4(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I5(CLBLM_R_X59Y112_SLICE_X89Y112_BQ),
.O5(CLBLM_R_X59Y105_SLICE_X89Y105_DO5),
.O6(CLBLM_R_X59Y105_SLICE_X89Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff22223022)
  ) CLBLM_R_X59Y105_SLICE_X89Y105_CLUT (
.I0(CLBLM_L_X60Y108_SLICE_X90Y108_B_XOR),
.I1(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I2(CLBLM_R_X59Y107_SLICE_X89Y107_B_XOR),
.I3(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I4(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I5(CLBLM_L_X62Y105_SLICE_X92Y105_AO6),
.O5(CLBLM_R_X59Y105_SLICE_X89Y105_CO5),
.O6(CLBLM_R_X59Y105_SLICE_X89Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aaaaff00f0f0)
  ) CLBLM_R_X59Y105_SLICE_X89Y105_BLUT (
.I0(CLBLM_R_X49Y111_SLICE_X74Y111_CQ),
.I1(1'b1),
.I2(CLBLM_R_X63Y110_SLICE_X94Y110_AQ),
.I3(CLBLM_L_X64Y106_SLICE_X96Y106_AQ),
.I4(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I5(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.O5(CLBLM_R_X59Y105_SLICE_X89Y105_BO5),
.O6(CLBLM_R_X59Y105_SLICE_X89Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000aaccaacc)
  ) CLBLM_R_X59Y105_SLICE_X89Y105_ALUT (
.I0(CLBLM_L_X56Y105_SLICE_X85Y105_CQ),
.I1(CLBLM_L_X56Y105_SLICE_X84Y105_CQ),
.I2(CLBLL_R_X57Y108_SLICE_X87Y108_BQ),
.I3(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I4(CLBLM_R_X59Y108_SLICE_X88Y108_AQ),
.I5(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.O5(CLBLM_R_X59Y105_SLICE_X89Y105_AO5),
.O6(CLBLM_R_X59Y105_SLICE_X89Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X59Y105_SLICE_X89Y105_MUXF7A (
.I0(CLBLM_R_X59Y105_SLICE_X89Y105_BO6),
.I1(CLBLM_R_X59Y105_SLICE_X89Y105_AO6),
.O(CLBLM_R_X59Y105_SLICE_X89Y105_F7AMUX_O),
.S(CLBLM_L_X62Y106_SLICE_X93Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y106_SLICE_X88Y106_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y100_SLICE_X90Y100_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y106_SLICE_X88Y106_AO6),
.Q(CLBLM_R_X59Y106_SLICE_X88Y106_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y106_SLICE_X88Y106_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y100_SLICE_X90Y100_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y106_SLICE_X88Y106_BO6),
.Q(CLBLM_R_X59Y106_SLICE_X88Y106_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffffffffffffff)
  ) CLBLM_R_X59Y106_SLICE_X88Y106_DLUT (
.I0(CLBLL_R_X57Y106_SLICE_X87Y106_AQ),
.I1(CLBLM_R_X59Y107_SLICE_X88Y107_AQ),
.I2(CLBLM_R_X59Y99_SLICE_X89Y99_BQ),
.I3(CLBLM_R_X59Y99_SLICE_X88Y99_CQ),
.I4(CLBLM_R_X59Y99_SLICE_X88Y99_AQ),
.I5(CLBLM_R_X59Y99_SLICE_X88Y99_DQ),
.O5(CLBLM_R_X59Y106_SLICE_X88Y106_DO5),
.O6(CLBLM_R_X59Y106_SLICE_X88Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33e2e2cc00e2e2)
  ) CLBLM_R_X59Y106_SLICE_X88Y106_CLUT (
.I0(CLBLM_R_X59Y104_SLICE_X88Y104_AQ),
.I1(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I2(CLBLL_R_X57Y106_SLICE_X86Y106_C_XOR),
.I3(CLBLL_R_X57Y105_SLICE_X86Y105_BQ),
.I4(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I5(CLBLL_R_X57Y109_SLICE_X87Y109_D_XOR),
.O5(CLBLM_R_X59Y106_SLICE_X88Y106_CO5),
.O6(CLBLM_R_X59Y106_SLICE_X88Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff23ff33ff20ff00)
  ) CLBLM_R_X59Y106_SLICE_X88Y106_BLUT (
.I0(CLBLL_R_X57Y105_SLICE_X87Y105_A_XOR),
.I1(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I2(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I3(CLBLM_L_X62Y103_SLICE_X93Y103_AO6),
.I4(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I5(CLBLL_R_X57Y106_SLICE_X86Y106_A_XOR),
.O5(CLBLM_R_X59Y106_SLICE_X88Y106_BO5),
.O6(CLBLM_R_X59Y106_SLICE_X88Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff33201300)
  ) CLBLM_R_X59Y106_SLICE_X88Y106_ALUT (
.I0(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I1(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I2(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I3(CLBLL_R_X57Y107_SLICE_X86Y107_C_XOR),
.I4(CLBLL_R_X57Y106_SLICE_X87Y106_C_XOR),
.I5(CLBLM_L_X62Y107_SLICE_X92Y107_BO5),
.O5(CLBLM_R_X59Y106_SLICE_X88Y106_AO5),
.O6(CLBLM_R_X59Y106_SLICE_X88Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y106_SLICE_X89Y106_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y99_SLICE_X90Y99_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y106_SLICE_X89Y106_BO6),
.Q(CLBLM_R_X59Y106_SLICE_X89Y106_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y106_SLICE_X89Y106_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y99_SLICE_X90Y99_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y106_SLICE_X89Y106_CO6),
.Q(CLBLM_R_X59Y106_SLICE_X89Y106_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafaee445050ee44)
  ) CLBLM_R_X59Y106_SLICE_X89Y106_DLUT (
.I0(CLBLM_R_X59Y106_SLICE_X89Y106_AO6),
.I1(CLBLM_R_X59Y106_SLICE_X88Y106_CO6),
.I2(CLBLM_L_X60Y108_SLICE_X90Y108_C_XOR),
.I3(CLBLL_R_X57Y105_SLICE_X86Y105_BQ),
.I4(CLBLM_L_X62Y106_SLICE_X92Y106_AO5),
.I5(CLBLM_R_X59Y108_SLICE_X88Y108_D_XOR),
.O5(CLBLM_R_X59Y106_SLICE_X89Y106_DO5),
.O6(CLBLM_R_X59Y106_SLICE_X89Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff54ff04ff55ff00)
  ) CLBLM_R_X59Y106_SLICE_X89Y106_CLUT (
.I0(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I1(CLBLM_R_X59Y107_SLICE_X89Y107_A_XOR),
.I2(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I3(CLBLM_L_X62Y103_SLICE_X93Y103_AO6),
.I4(CLBLM_L_X60Y108_SLICE_X90Y108_A_XOR),
.I5(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.O5(CLBLM_R_X59Y106_SLICE_X89Y106_CO5),
.O6(CLBLM_R_X59Y106_SLICE_X89Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff44544404)
  ) CLBLM_R_X59Y106_SLICE_X89Y106_BLUT (
.I0(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I1(CLBLM_L_X60Y109_SLICE_X90Y109_C_XOR),
.I2(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I3(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I4(CLBLM_R_X59Y108_SLICE_X89Y108_C_XOR),
.I5(CLBLM_L_X62Y107_SLICE_X92Y107_BO5),
.O5(CLBLM_R_X59Y106_SLICE_X89Y106_BO5),
.O6(CLBLM_R_X59Y106_SLICE_X89Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f00ff00acaccccc)
  ) CLBLM_R_X59Y106_SLICE_X89Y106_ALUT (
.I0(CLBLM_L_X60Y106_SLICE_X90Y106_A_XOR),
.I1(CLBLM_L_X60Y104_SLICE_X90Y104_AQ),
.I2(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I3(CLBLM_R_X59Y103_SLICE_X89Y103_CQ),
.I4(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I5(1'b1),
.O5(CLBLM_R_X59Y106_SLICE_X89Y106_AO5),
.O6(CLBLM_R_X59Y106_SLICE_X89Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X59Y107_SLICE_X88Y107_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLL_R_X57Y99_SLICE_X87Y99_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X49Y107_SLICE_X75Y107_CQ),
.Q(CLBLM_R_X59Y107_SLICE_X88Y107_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaf0ffccaaf000)
  ) CLBLM_R_X59Y107_SLICE_X88Y107_DLUT (
.I0(CLBLL_R_X57Y107_SLICE_X86Y107_C_XOR),
.I1(CLBLM_R_X59Y106_SLICE_X88Y106_AQ),
.I2(CLBLL_R_X57Y110_SLICE_X87Y110_D_XOR),
.I3(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I4(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I5(CLBLM_R_X59Y107_SLICE_X88Y107_AQ),
.O5(CLBLM_R_X59Y107_SLICE_X88Y107_DO5),
.O6(CLBLM_R_X59Y107_SLICE_X88Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcaffcaf0ca0fca00)
  ) CLBLM_R_X59Y107_SLICE_X88Y107_CLUT (
.I0(CLBLM_R_X59Y106_SLICE_X88Y106_AQ),
.I1(CLBLM_R_X59Y109_SLICE_X88Y109_D_XOR),
.I2(CLBLM_L_X62Y106_SLICE_X92Y106_AO5),
.I3(CLBLM_R_X59Y106_SLICE_X89Y106_AO6),
.I4(CLBLM_R_X59Y107_SLICE_X88Y107_DO6),
.I5(CLBLM_L_X60Y109_SLICE_X90Y109_C_XOR),
.O5(CLBLM_R_X59Y107_SLICE_X88Y107_CO5),
.O6(CLBLM_R_X59Y107_SLICE_X88Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa00aaccf0ccf0)
  ) CLBLM_R_X59Y107_SLICE_X88Y107_BLUT (
.I0(CLBLL_R_X57Y109_SLICE_X87Y109_B_XOR),
.I1(CLBLL_R_X57Y106_SLICE_X86Y106_A_XOR),
.I2(CLBLM_R_X59Y103_SLICE_X88Y103_CQ),
.I3(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I4(CLBLM_R_X59Y106_SLICE_X88Y106_BQ),
.I5(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.O5(CLBLM_R_X59Y107_SLICE_X88Y107_BO5),
.O6(CLBLM_R_X59Y107_SLICE_X88Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b8b8b8ffcc3300)
  ) CLBLM_R_X59Y107_SLICE_X88Y107_ALUT (
.I0(CLBLM_R_X59Y108_SLICE_X88Y108_B_XOR),
.I1(CLBLM_L_X62Y106_SLICE_X92Y106_AO5),
.I2(CLBLM_R_X59Y106_SLICE_X88Y106_BQ),
.I3(CLBLM_R_X59Y107_SLICE_X88Y107_BO6),
.I4(CLBLM_L_X60Y108_SLICE_X90Y108_A_XOR),
.I5(CLBLM_R_X59Y106_SLICE_X89Y106_AO6),
.O5(CLBLM_R_X59Y107_SLICE_X88Y107_AO5),
.O6(CLBLM_R_X59Y107_SLICE_X88Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X59Y107_SLICE_X89Y107_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLL_R_X57Y99_SLICE_X87Y99_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y107_SLICE_X89Y107_BO5),
.Q(CLBLM_R_X59Y107_SLICE_X89Y107_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X59Y107_SLICE_X89Y107_CARRY4 (
.CI(1'b0),
.CO({CLBLM_R_X59Y107_SLICE_X89Y107_D_CY, CLBLM_R_X59Y107_SLICE_X89Y107_C_CY, CLBLM_R_X59Y107_SLICE_X89Y107_B_CY, CLBLM_R_X59Y107_SLICE_X89Y107_A_CY}),
.CYINIT(CLBLM_L_X60Y100_SLICE_X90Y100_AQ),
.DI({CLBLM_L_X60Y104_SLICE_X90Y104_AQ, CLBLM_R_X59Y104_SLICE_X89Y104_CQ, CLBLM_R_X59Y105_SLICE_X89Y105_CQ, CLBLM_R_X59Y107_SLICE_X89Y107_AO5}),
.O({CLBLM_R_X59Y107_SLICE_X89Y107_D_XOR, CLBLM_R_X59Y107_SLICE_X89Y107_C_XOR, CLBLM_R_X59Y107_SLICE_X89Y107_B_XOR, CLBLM_R_X59Y107_SLICE_X89Y107_A_XOR}),
.S({CLBLM_R_X59Y107_SLICE_X89Y107_DO6, CLBLM_R_X59Y107_SLICE_X89Y107_CO6, CLBLM_R_X59Y107_SLICE_X89Y107_BO6, CLBLM_R_X59Y107_SLICE_X89Y107_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00ff00ff)
  ) CLBLM_R_X59Y107_SLICE_X89Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X60Y104_SLICE_X90Y104_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y107_SLICE_X89Y107_DO5),
.O6(CLBLM_R_X59Y107_SLICE_X89Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333333333333)
  ) CLBLM_R_X59Y107_SLICE_X89Y107_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X59Y104_SLICE_X89Y104_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y107_SLICE_X89Y107_CO5),
.O6(CLBLM_R_X59Y107_SLICE_X89Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffffcccccccc)
  ) CLBLM_R_X59Y107_SLICE_X89Y107_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X49Y104_SLICE_X75Y104_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X59Y105_SLICE_X89Y105_CQ),
.I5(1'b1),
.O5(CLBLM_R_X59Y107_SLICE_X89Y107_BO5),
.O6(CLBLM_R_X59Y107_SLICE_X89Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ffff00ff00)
  ) CLBLM_R_X59Y107_SLICE_X89Y107_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X59Y106_SLICE_X89Y106_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y107_SLICE_X89Y107_AO5),
.O6(CLBLM_R_X59Y107_SLICE_X89Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y108_SLICE_X88Y108_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y100_SLICE_X90Y100_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y108_SLICE_X88Y108_AO5),
.Q(CLBLM_R_X59Y108_SLICE_X88Y108_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X59Y108_SLICE_X88Y108_CARRY4 (
.CI(1'b0),
.CO({CLBLM_R_X59Y108_SLICE_X88Y108_D_CY, CLBLM_R_X59Y108_SLICE_X88Y108_C_CY, CLBLM_R_X59Y108_SLICE_X88Y108_B_CY, CLBLM_R_X59Y108_SLICE_X88Y108_A_CY}),
.CYINIT(1'b0),
.DI({CLBLM_R_X59Y104_SLICE_X89Y104_CQ, CLBLM_R_X59Y105_SLICE_X89Y105_CQ, CLBLM_R_X59Y106_SLICE_X89Y106_CQ, CLBLM_L_X60Y100_SLICE_X90Y100_AQ}),
.O({CLBLM_R_X59Y108_SLICE_X88Y108_D_XOR, CLBLM_R_X59Y108_SLICE_X88Y108_C_XOR, CLBLM_R_X59Y108_SLICE_X88Y108_B_XOR, CLBLM_R_X59Y108_SLICE_X88Y108_A_XOR}),
.S({CLBLM_R_X59Y108_SLICE_X88Y108_DO6, CLBLM_R_X59Y108_SLICE_X88Y108_CO6, CLBLM_R_X59Y108_SLICE_X88Y108_BO6, CLBLM_R_X59Y108_SLICE_X88Y108_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555555aaaaaaaa)
  ) CLBLM_R_X59Y108_SLICE_X88Y108_DLUT (
.I0(CLBLM_R_X59Y104_SLICE_X89Y104_CQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X59Y98_SLICE_X89Y98_B5Q),
.O5(CLBLM_R_X59Y108_SLICE_X88Y108_DO5),
.O6(CLBLM_R_X59Y108_SLICE_X88Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa55aa55aa55aa)
  ) CLBLM_R_X59Y108_SLICE_X88Y108_CLUT (
.I0(CLBLM_R_X59Y98_SLICE_X89Y98_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X59Y105_SLICE_X89Y105_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y108_SLICE_X88Y108_CO5),
.O6(CLBLM_R_X59Y108_SLICE_X88Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333333cccccccc)
  ) CLBLM_R_X59Y108_SLICE_X88Y108_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X59Y106_SLICE_X89Y106_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X59Y98_SLICE_X89Y98_A5Q),
.O5(CLBLM_R_X59Y108_SLICE_X88Y108_BO5),
.O6(CLBLM_R_X59Y108_SLICE_X88Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ccccf0f0f0f0)
  ) CLBLM_R_X59Y108_SLICE_X88Y108_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X59Y98_SLICE_X89Y98_AQ),
.I2(CLBLM_L_X62Y108_SLICE_X92Y108_BO6),
.I3(1'b1),
.I4(CLBLM_L_X60Y100_SLICE_X90Y100_AQ),
.I5(1'b1),
.O5(CLBLM_R_X59Y108_SLICE_X88Y108_AO5),
.O6(CLBLM_R_X59Y108_SLICE_X88Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y108_SLICE_X89Y108_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y100_SLICE_X90Y100_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y108_SLICE_X89Y108_AO5),
.Q(CLBLM_R_X59Y108_SLICE_X89Y108_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X59Y108_SLICE_X89Y108_CARRY4 (
.CI(CLBLM_R_X59Y107_SLICE_X89Y107_COUT),
.CO({CLBLM_R_X59Y108_SLICE_X89Y108_D_CY, CLBLM_R_X59Y108_SLICE_X89Y108_C_CY, CLBLM_R_X59Y108_SLICE_X89Y108_B_CY, CLBLM_R_X59Y108_SLICE_X89Y108_A_CY}),
.CYINIT(1'b0),
.DI({CLBLM_R_X59Y111_SLICE_X89Y111_CQ, CLBLM_R_X59Y106_SLICE_X89Y106_BQ, CLBLM_R_X59Y112_SLICE_X89Y112_BQ, CLBLM_R_X59Y112_SLICE_X89Y112_AQ}),
.O({CLBLM_R_X59Y108_SLICE_X89Y108_D_XOR, CLBLM_R_X59Y108_SLICE_X89Y108_C_XOR, CLBLM_R_X59Y108_SLICE_X89Y108_B_XOR, CLBLM_R_X59Y108_SLICE_X89Y108_A_XOR}),
.S({CLBLM_R_X59Y108_SLICE_X89Y108_DO6, CLBLM_R_X59Y108_SLICE_X89Y108_CO6, CLBLM_R_X59Y108_SLICE_X89Y108_BO6, CLBLM_R_X59Y108_SLICE_X89Y108_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333333333333)
  ) CLBLM_R_X59Y108_SLICE_X89Y108_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X59Y111_SLICE_X89Y111_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y108_SLICE_X89Y108_DO5),
.O6(CLBLM_R_X59Y108_SLICE_X89Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555555)
  ) CLBLM_R_X59Y108_SLICE_X89Y108_CLUT (
.I0(CLBLM_R_X59Y106_SLICE_X89Y106_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y108_SLICE_X89Y108_CO5),
.O6(CLBLM_R_X59Y108_SLICE_X89Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333333333333)
  ) CLBLM_R_X59Y108_SLICE_X89Y108_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X59Y112_SLICE_X89Y112_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y108_SLICE_X89Y108_BO5),
.O6(CLBLM_R_X59Y108_SLICE_X89Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0fff00ff00)
  ) CLBLM_R_X59Y108_SLICE_X89Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X59Y112_SLICE_X89Y112_AQ),
.I3(CLBLM_L_X62Y108_SLICE_X92Y108_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y108_SLICE_X89Y108_AO5),
.O6(CLBLM_R_X59Y108_SLICE_X89Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X59Y109_SLICE_X88Y109_CARRY4 (
.CI(CLBLM_R_X59Y108_SLICE_X88Y108_COUT),
.CO({CLBLM_R_X59Y109_SLICE_X88Y109_D_CY, CLBLM_R_X59Y109_SLICE_X88Y109_C_CY, CLBLM_R_X59Y109_SLICE_X88Y109_B_CY, CLBLM_R_X59Y109_SLICE_X88Y109_A_CY}),
.CYINIT(1'b0),
.DI({CLBLM_R_X59Y106_SLICE_X89Y106_BQ, CLBLM_R_X59Y112_SLICE_X89Y112_BQ, CLBLM_R_X59Y112_SLICE_X89Y112_AQ, CLBLM_L_X60Y104_SLICE_X90Y104_AQ}),
.O({CLBLM_R_X59Y109_SLICE_X88Y109_D_XOR, CLBLM_R_X59Y109_SLICE_X88Y109_C_XOR, CLBLM_R_X59Y109_SLICE_X88Y109_B_XOR, CLBLM_R_X59Y109_SLICE_X88Y109_A_XOR}),
.S({CLBLM_R_X59Y109_SLICE_X88Y109_DO6, CLBLM_R_X59Y109_SLICE_X88Y109_CO6, CLBLM_R_X59Y109_SLICE_X88Y109_BO6, CLBLM_R_X59Y109_SLICE_X88Y109_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5a5a5a5a5a)
  ) CLBLM_R_X59Y109_SLICE_X88Y109_DLUT (
.I0(CLBLM_R_X59Y106_SLICE_X89Y106_BQ),
.I1(1'b1),
.I2(CLBLM_R_X59Y96_SLICE_X89Y96_A5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y109_SLICE_X88Y109_DO5),
.O6(CLBLM_R_X59Y109_SLICE_X88Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0ff0f0f0f0)
  ) CLBLM_R_X59Y109_SLICE_X88Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X59Y96_SLICE_X89Y96_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X59Y112_SLICE_X89Y112_BQ),
.O5(CLBLM_R_X59Y109_SLICE_X88Y109_CO5),
.O6(CLBLM_R_X59Y109_SLICE_X88Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0ff0f00f0ff0f0)
  ) CLBLM_R_X59Y109_SLICE_X88Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X59Y98_SLICE_X89Y98_C5Q),
.I3(1'b1),
.I4(CLBLM_R_X59Y112_SLICE_X89Y112_AQ),
.I5(1'b1),
.O5(CLBLM_R_X59Y109_SLICE_X88Y109_BO5),
.O6(CLBLM_R_X59Y109_SLICE_X88Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333cccc3333cccc)
  ) CLBLM_R_X59Y109_SLICE_X88Y109_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X59Y98_SLICE_X89Y98_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X60Y104_SLICE_X90Y104_AQ),
.I5(1'b1),
.O5(CLBLM_R_X59Y109_SLICE_X88Y109_AO5),
.O6(CLBLM_R_X59Y109_SLICE_X88Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X59Y109_SLICE_X89Y109_CARRY4 (
.CI(CLBLM_R_X59Y108_SLICE_X89Y108_COUT),
.CO({CLBLM_R_X59Y109_SLICE_X89Y109_D_CY, CLBLM_R_X59Y109_SLICE_X89Y109_C_CY, CLBLM_R_X59Y109_SLICE_X89Y109_B_CY, CLBLM_R_X59Y109_SLICE_X89Y109_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, CLBLM_R_X59Y111_SLICE_X89Y111_BQ, CLBLM_R_X59Y111_SLICE_X89Y111_AQ}),
.O({CLBLM_R_X59Y109_SLICE_X89Y109_D_XOR, CLBLM_R_X59Y109_SLICE_X89Y109_C_XOR, CLBLM_R_X59Y109_SLICE_X89Y109_B_XOR, CLBLM_R_X59Y109_SLICE_X89Y109_A_XOR}),
.S({CLBLM_R_X59Y109_SLICE_X89Y109_DO6, CLBLM_R_X59Y109_SLICE_X89Y109_CO6, CLBLM_R_X59Y109_SLICE_X89Y109_BO6, CLBLM_R_X59Y109_SLICE_X89Y109_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X59Y109_SLICE_X89Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y109_SLICE_X89Y109_DO5),
.O6(CLBLM_R_X59Y109_SLICE_X89Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333333333333)
  ) CLBLM_R_X59Y109_SLICE_X89Y109_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X59Y110_SLICE_X89Y110_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y109_SLICE_X89Y109_CO5),
.O6(CLBLM_R_X59Y109_SLICE_X89Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffffffff)
  ) CLBLM_R_X59Y109_SLICE_X89Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X59Y111_SLICE_X89Y111_BQ),
.O5(CLBLM_R_X59Y109_SLICE_X89Y109_BO5),
.O6(CLBLM_R_X59Y109_SLICE_X89Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00ff00ff)
  ) CLBLM_R_X59Y109_SLICE_X89Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X59Y111_SLICE_X89Y111_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y109_SLICE_X89Y109_AO5),
.O6(CLBLM_R_X59Y109_SLICE_X89Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X59Y110_SLICE_X88Y110_CARRY4 (
.CI(CLBLM_R_X59Y109_SLICE_X88Y109_COUT),
.CO({CLBLM_R_X59Y110_SLICE_X88Y110_D_CY, CLBLM_R_X59Y110_SLICE_X88Y110_C_CY, CLBLM_R_X59Y110_SLICE_X88Y110_B_CY, CLBLM_R_X59Y110_SLICE_X88Y110_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X59Y110_SLICE_X88Y110_D_XOR, CLBLM_R_X59Y110_SLICE_X88Y110_C_XOR, CLBLM_R_X59Y110_SLICE_X88Y110_B_XOR, CLBLM_R_X59Y110_SLICE_X88Y110_A_XOR}),
.S({CLBLM_R_X59Y110_SLICE_X88Y110_DO6, CLBLM_R_X59Y110_SLICE_X88Y110_CO6, CLBLM_R_X59Y110_SLICE_X88Y110_BO6, CLBLM_R_X59Y110_SLICE_X88Y110_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X59Y110_SLICE_X88Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X59Y110_SLICE_X89Y110_AQ),
.O5(CLBLM_R_X59Y110_SLICE_X88Y110_DO5),
.O6(CLBLM_R_X59Y110_SLICE_X88Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X59Y110_SLICE_X88Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X59Y111_SLICE_X89Y111_BQ),
.O5(CLBLM_R_X59Y110_SLICE_X88Y110_CO5),
.O6(CLBLM_R_X59Y110_SLICE_X88Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X59Y110_SLICE_X88Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X59Y111_SLICE_X89Y111_AQ),
.O5(CLBLM_R_X59Y110_SLICE_X88Y110_BO5),
.O6(CLBLM_R_X59Y110_SLICE_X88Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X59Y110_SLICE_X88Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X59Y111_SLICE_X89Y111_CQ),
.O5(CLBLM_R_X59Y110_SLICE_X88Y110_AO5),
.O6(CLBLM_R_X59Y110_SLICE_X88Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y110_SLICE_X89Y110_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y100_SLICE_X90Y100_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y110_SLICE_X89Y110_AO6),
.Q(CLBLM_R_X59Y110_SLICE_X89Y110_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0ccffaaf0cc00)
  ) CLBLM_R_X59Y110_SLICE_X89Y110_DLUT (
.I0(CLBLL_R_X57Y108_SLICE_X87Y108_AQ),
.I1(CLBLL_R_X57Y107_SLICE_X86Y107_A_XOR),
.I2(CLBLL_R_X57Y110_SLICE_X87Y110_B_XOR),
.I3(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I4(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I5(CLBLM_R_X59Y104_SLICE_X88Y104_BQ),
.O5(CLBLM_R_X59Y110_SLICE_X89Y110_DO5),
.O6(CLBLM_R_X59Y110_SLICE_X89Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcaf0caffca00ca0)
  ) CLBLM_R_X59Y110_SLICE_X89Y110_CLUT (
.I0(CLBLL_R_X57Y108_SLICE_X87Y108_AQ),
.I1(CLBLM_L_X60Y109_SLICE_X90Y109_A_XOR),
.I2(CLBLM_R_X59Y106_SLICE_X89Y106_AO6),
.I3(CLBLM_L_X62Y106_SLICE_X92Y106_AO5),
.I4(CLBLM_R_X59Y109_SLICE_X88Y109_B_XOR),
.I5(CLBLM_R_X59Y110_SLICE_X89Y110_DO6),
.O5(CLBLM_R_X59Y110_SLICE_X89Y110_CO5),
.O6(CLBLM_R_X59Y110_SLICE_X89Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7e6d5c4b3a29180)
  ) CLBLM_R_X59Y110_SLICE_X89Y110_BLUT (
.I0(CLBLM_R_X59Y106_SLICE_X89Y106_AO6),
.I1(CLBLM_L_X62Y106_SLICE_X92Y106_AO5),
.I2(CLBLM_R_X59Y110_SLICE_X88Y110_C_XOR),
.I3(CLBLL_R_X57Y109_SLICE_X86Y109_DO6),
.I4(CLBLL_R_X57Y109_SLICE_X86Y109_BQ),
.I5(CLBLM_L_X60Y110_SLICE_X90Y110_B_XOR),
.O5(CLBLM_R_X59Y110_SLICE_X89Y110_BO5),
.O6(CLBLM_R_X59Y110_SLICE_X89Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffcce40000cce4)
  ) CLBLM_R_X59Y110_SLICE_X89Y110_ALUT (
.I0(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I1(CLBLM_L_X60Y110_SLICE_X90Y110_C_XOR),
.I2(CLBLM_R_X59Y109_SLICE_X89Y109_C_XOR),
.I3(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I4(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I5(CLBLM_L_X62Y100_SLICE_X93Y100_BO6),
.O5(CLBLM_R_X59Y110_SLICE_X89Y110_AO5),
.O6(CLBLM_R_X59Y110_SLICE_X89Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0f0ff00cccc)
  ) CLBLM_R_X59Y111_SLICE_X88Y111_DLUT (
.I0(CLBLL_R_X57Y109_SLICE_X86Y109_AQ),
.I1(CLBLM_R_X59Y99_SLICE_X88Y99_DQ),
.I2(CLBLL_R_X57Y111_SLICE_X87Y111_B_XOR),
.I3(CLBLL_R_X57Y108_SLICE_X86Y108_A_XOR),
.I4(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I5(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.O5(CLBLM_R_X59Y111_SLICE_X88Y111_DO5),
.O6(CLBLM_R_X59Y111_SLICE_X88Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he2ffe2cce233e200)
  ) CLBLM_R_X59Y111_SLICE_X88Y111_CLUT (
.I0(CLBLL_R_X57Y109_SLICE_X86Y109_AQ),
.I1(CLBLM_L_X62Y106_SLICE_X92Y106_AO5),
.I2(CLBLM_R_X59Y110_SLICE_X88Y110_B_XOR),
.I3(CLBLM_R_X59Y106_SLICE_X89Y106_AO6),
.I4(CLBLM_R_X59Y111_SLICE_X88Y111_DO6),
.I5(CLBLM_L_X60Y110_SLICE_X90Y110_A_XOR),
.O5(CLBLM_R_X59Y111_SLICE_X88Y111_CO5),
.O6(CLBLM_R_X59Y111_SLICE_X88Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffe233e2cce200e2)
  ) CLBLM_R_X59Y111_SLICE_X88Y111_BLUT (
.I0(CLBLM_R_X59Y99_SLICE_X88Y99_CQ),
.I1(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I2(CLBLL_R_X57Y107_SLICE_X86Y107_D_XOR),
.I3(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I4(CLBLM_L_X60Y108_SLICE_X91Y108_AQ),
.I5(CLBLL_R_X57Y111_SLICE_X87Y111_A_XOR),
.O5(CLBLM_R_X59Y111_SLICE_X88Y111_BO5),
.O6(CLBLM_R_X59Y111_SLICE_X88Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ee22f3f3c0c0)
  ) CLBLM_R_X59Y111_SLICE_X88Y111_ALUT (
.I0(CLBLL_R_X57Y111_SLICE_X87Y111_D_XOR),
.I1(CLBLM_R_X59Y103_SLICE_X89Y103_BQ),
.I2(CLBLL_R_X57Y108_SLICE_X86Y108_C_XOR),
.I3(CLBLL_R_X57Y109_SLICE_X86Y109_CQ),
.I4(CLBLM_R_X59Y99_SLICE_X88Y99_AQ),
.I5(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.O5(CLBLM_R_X59Y111_SLICE_X88Y111_AO5),
.O6(CLBLM_R_X59Y111_SLICE_X88Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y111_SLICE_X89Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y100_SLICE_X90Y100_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y111_SLICE_X89Y111_AO6),
.Q(CLBLM_R_X59Y111_SLICE_X89Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y111_SLICE_X89Y111_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y100_SLICE_X90Y100_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y111_SLICE_X89Y111_BO6),
.Q(CLBLM_R_X59Y111_SLICE_X89Y111_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y111_SLICE_X89Y111_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y100_SLICE_X90Y100_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y111_SLICE_X89Y111_CO6),
.Q(CLBLM_R_X59Y111_SLICE_X89Y111_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0aacc00f0aacc)
  ) CLBLM_R_X59Y111_SLICE_X89Y111_DLUT (
.I0(CLBLM_L_X60Y110_SLICE_X90Y110_C_XOR),
.I1(CLBLM_R_X59Y111_SLICE_X88Y111_AO6),
.I2(CLBLL_R_X57Y109_SLICE_X86Y109_CQ),
.I3(CLBLM_L_X62Y106_SLICE_X92Y106_AO5),
.I4(CLBLM_R_X59Y106_SLICE_X89Y106_AO6),
.I5(CLBLM_R_X59Y110_SLICE_X88Y110_D_XOR),
.O5(CLBLM_R_X59Y111_SLICE_X89Y111_DO5),
.O6(CLBLM_R_X59Y111_SLICE_X89Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ee22f0f0ff00)
  ) CLBLM_R_X59Y111_SLICE_X89Y111_CLUT (
.I0(CLBLM_R_X59Y108_SLICE_X89Y108_D_XOR),
.I1(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I2(CLBLM_L_X62Y97_SLICE_X92Y97_AO6),
.I3(CLBLM_L_X60Y109_SLICE_X90Y109_D_XOR),
.I4(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I5(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.O5(CLBLM_R_X59Y111_SLICE_X89Y111_CO5),
.O6(CLBLM_R_X59Y111_SLICE_X89Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffb00fbff080008)
  ) CLBLM_R_X59Y111_SLICE_X89Y111_BLUT (
.I0(CLBLM_R_X59Y109_SLICE_X89Y109_B_XOR),
.I1(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I2(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I3(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I4(CLBLM_L_X62Y100_SLICE_X93Y100_AO6),
.I5(CLBLM_L_X60Y110_SLICE_X90Y110_B_XOR),
.O5(CLBLM_R_X59Y111_SLICE_X89Y111_BO5),
.O6(CLBLM_R_X59Y111_SLICE_X89Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hefee4544eaee4044)
  ) CLBLM_R_X59Y111_SLICE_X89Y111_ALUT (
.I0(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I1(CLBLM_L_X60Y110_SLICE_X90Y110_A_XOR),
.I2(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I3(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I4(CLBLM_L_X62Y97_SLICE_X92Y97_BO6),
.I5(CLBLM_R_X59Y109_SLICE_X89Y109_A_XOR),
.O5(CLBLM_R_X59Y111_SLICE_X89Y111_AO5),
.O6(CLBLM_R_X59Y111_SLICE_X89Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X59Y112_SLICE_X88Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y112_SLICE_X88Y112_DO5),
.O6(CLBLM_R_X59Y112_SLICE_X88Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X59Y112_SLICE_X88Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y112_SLICE_X88Y112_CO5),
.O6(CLBLM_R_X59Y112_SLICE_X88Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X59Y112_SLICE_X88Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y112_SLICE_X88Y112_BO5),
.O6(CLBLM_R_X59Y112_SLICE_X88Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X59Y112_SLICE_X88Y112_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y112_SLICE_X88Y112_AO5),
.O6(CLBLM_R_X59Y112_SLICE_X88Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y112_SLICE_X89Y112_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y99_SLICE_X90Y99_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y112_SLICE_X89Y112_AO6),
.Q(CLBLM_R_X59Y112_SLICE_X89Y112_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y112_SLICE_X89Y112_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y99_SLICE_X90Y99_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X59Y112_SLICE_X89Y112_BO6),
.Q(CLBLM_R_X59Y112_SLICE_X89Y112_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X59Y112_SLICE_X89Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y112_SLICE_X89Y112_DO5),
.O6(CLBLM_R_X59Y112_SLICE_X89Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbfcbb3088fc8830)
  ) CLBLM_R_X59Y112_SLICE_X89Y112_CLUT (
.I0(CLBLM_R_X59Y109_SLICE_X88Y109_C_XOR),
.I1(CLBLM_L_X62Y106_SLICE_X92Y106_AO5),
.I2(CLBLL_R_X57Y108_SLICE_X87Y108_DO6),
.I3(CLBLM_R_X59Y106_SLICE_X89Y106_AO6),
.I4(CLBLM_L_X60Y109_SLICE_X90Y109_B_XOR),
.I5(CLBLL_R_X57Y108_SLICE_X87Y108_BQ),
.O5(CLBLM_R_X59Y112_SLICE_X89Y112_CO5),
.O6(CLBLM_R_X59Y112_SLICE_X89Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fbfaf0f0f8fa)
  ) CLBLM_R_X59Y112_SLICE_X89Y112_BLUT (
.I0(CLBLM_L_X60Y109_SLICE_X90Y109_B_XOR),
.I1(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I2(CLBLM_L_X62Y108_SLICE_X92Y108_BO5),
.I3(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I4(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I5(CLBLM_R_X59Y108_SLICE_X89Y108_B_XOR),
.O5(CLBLM_R_X59Y112_SLICE_X89Y112_BO5),
.O6(CLBLM_R_X59Y112_SLICE_X89Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafbfaaaaaeafa)
  ) CLBLM_R_X59Y112_SLICE_X89Y112_ALUT (
.I0(CLBLM_L_X62Y106_SLICE_X93Y106_BO5),
.I1(CLBLM_R_X59Y103_SLICE_X89Y103_AQ),
.I2(CLBLM_L_X60Y109_SLICE_X90Y109_A_XOR),
.I3(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I4(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I5(CLBLM_R_X59Y108_SLICE_X89Y108_A_XOR),
.O5(CLBLM_R_X59Y112_SLICE_X89Y112_AO5),
.O6(CLBLM_R_X59Y112_SLICE_X89Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y94_SLICE_X94Y94_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y99_SLICE_X93Y99_AO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y94_SLICE_X94Y94_AO6),
.Q(CLBLM_R_X63Y94_SLICE_X94Y94_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y94_SLICE_X94Y94_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y94_SLICE_X94Y94_DO5),
.O6(CLBLM_R_X63Y94_SLICE_X94Y94_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y94_SLICE_X94Y94_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y94_SLICE_X94Y94_CO5),
.O6(CLBLM_R_X63Y94_SLICE_X94Y94_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y94_SLICE_X94Y94_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y94_SLICE_X94Y94_BO5),
.O6(CLBLM_R_X63Y94_SLICE_X94Y94_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc5cfc5cac0cac0)
  ) CLBLM_R_X63Y94_SLICE_X94Y94_ALUT (
.I0(CLBLM_L_X56Y98_SLICE_X85Y98_DQ),
.I1(CLBLM_L_X50Y107_SLICE_X77Y107_AQ),
.I2(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I3(CLBLM_R_X63Y99_SLICE_X95Y99_A5Q),
.I4(1'b1),
.I5(CLBLM_R_X63Y96_SLICE_X94Y96_BO6),
.O5(CLBLM_R_X63Y94_SLICE_X94Y94_AO5),
.O6(CLBLM_R_X63Y94_SLICE_X94Y94_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y94_SLICE_X95Y94_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y99_SLICE_X93Y99_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y94_SLICE_X95Y94_AO6),
.Q(CLBLM_R_X63Y94_SLICE_X95Y94_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y94_SLICE_X95Y94_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y94_SLICE_X95Y94_DO5),
.O6(CLBLM_R_X63Y94_SLICE_X95Y94_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y94_SLICE_X95Y94_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y94_SLICE_X95Y94_CO5),
.O6(CLBLM_R_X63Y94_SLICE_X95Y94_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y94_SLICE_X95Y94_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y94_SLICE_X95Y94_BO5),
.O6(CLBLM_R_X63Y94_SLICE_X95Y94_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf505f505f000f000)
  ) CLBLM_R_X63Y94_SLICE_X95Y94_ALUT (
.I0(CLBLM_L_X56Y98_SLICE_X85Y98_DQ),
.I1(1'b1),
.I2(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I3(CLBLM_L_X50Y104_SLICE_X76Y104_AQ),
.I4(1'b1),
.I5(CLBLM_L_X64Y95_SLICE_X96Y95_AO5),
.O5(CLBLM_R_X63Y94_SLICE_X95Y94_AO5),
.O6(CLBLM_R_X63Y94_SLICE_X95Y94_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y95_SLICE_X95Y95_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y99_SLICE_X93Y99_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y95_SLICE_X95Y95_AO5),
.Q(CLBLM_R_X63Y95_SLICE_X95Y95_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y95_SLICE_X95Y95_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y99_SLICE_X93Y99_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y97_SLICE_X93Y97_CO5),
.Q(CLBLM_R_X63Y95_SLICE_X95Y95_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y95_SLICE_X95Y95_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y99_SLICE_X93Y99_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y96_SLICE_X95Y96_AO5),
.Q(CLBLM_R_X63Y95_SLICE_X95Y95_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y95_SLICE_X95Y95_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y99_SLICE_X93Y99_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y97_SLICE_X94Y97_CO5),
.Q(CLBLM_R_X63Y95_SLICE_X95Y95_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y95_SLICE_X95Y95_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y99_SLICE_X93Y99_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y95_SLICE_X95Y95_BO6),
.Q(CLBLM_R_X63Y95_SLICE_X95Y95_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y95_SLICE_X95Y95_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y99_SLICE_X93Y99_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y95_SLICE_X95Y95_CO6),
.Q(CLBLM_R_X63Y95_SLICE_X95Y95_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y95_SLICE_X95Y95_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y99_SLICE_X93Y99_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y95_SLICE_X95Y95_DO6),
.Q(CLBLM_R_X63Y95_SLICE_X95Y95_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ff55ee44aa00)
  ) CLBLM_R_X63Y95_SLICE_X95Y95_DLUT (
.I0(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I1(CLBLM_R_X63Y99_SLICE_X95Y99_B5Q),
.I2(1'b1),
.I3(CLBLM_L_X50Y105_SLICE_X77Y105_AQ),
.I4(CLBLM_L_X56Y98_SLICE_X85Y98_DQ),
.I5(CLBLM_L_X64Y95_SLICE_X96Y95_AO6),
.O5(CLBLM_R_X63Y95_SLICE_X95Y95_DO5),
.O6(CLBLM_R_X63Y95_SLICE_X95Y95_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfcacac0c0caca)
  ) CLBLM_R_X63Y95_SLICE_X95Y95_CLUT (
.I0(CLBLM_L_X64Y95_SLICE_X96Y95_BO6),
.I1(CLBLM_R_X49Y106_SLICE_X74Y106_AQ),
.I2(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I3(1'b1),
.I4(CLBLM_L_X56Y98_SLICE_X85Y98_DQ),
.I5(CLBLM_R_X63Y99_SLICE_X95Y99_C5Q),
.O5(CLBLM_R_X63Y95_SLICE_X95Y95_CO5),
.O6(CLBLM_R_X63Y95_SLICE_X95Y95_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffaff5000fa0050)
  ) CLBLM_R_X63Y95_SLICE_X95Y95_BLUT (
.I0(CLBLM_L_X56Y98_SLICE_X85Y98_DQ),
.I1(1'b1),
.I2(CLBLM_L_X64Y95_SLICE_X96Y95_BO5),
.I3(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I4(CLBLM_R_X63Y99_SLICE_X95Y99_CQ),
.I5(CLBLM_R_X49Y105_SLICE_X75Y105_CQ),
.O5(CLBLM_R_X63Y95_SLICE_X95Y95_BO5),
.O6(CLBLM_R_X63Y95_SLICE_X95Y95_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000f0eef044)
  ) CLBLM_R_X63Y95_SLICE_X95Y95_ALUT (
.I0(CLBLM_L_X56Y98_SLICE_X85Y98_DQ),
.I1(CLBLM_L_X64Y95_SLICE_X96Y95_CO6),
.I2(CLBLM_L_X50Y106_SLICE_X76Y106_CQ),
.I3(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I4(CLBLM_R_X63Y98_SLICE_X95Y98_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X63Y95_SLICE_X95Y95_AO5),
.O6(CLBLM_R_X63Y95_SLICE_X95Y95_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y96_SLICE_X95Y96_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y99_SLICE_X93Y99_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y95_SLICE_X95Y95_AO6),
.Q(CLBLM_R_X63Y96_SLICE_X95Y96_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y96_SLICE_X95Y96_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y99_SLICE_X93Y99_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y96_SLICE_X95Y96_BO6),
.Q(CLBLM_R_X63Y96_SLICE_X95Y96_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y96_SLICE_X95Y96_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y96_SLICE_X95Y96_DO5),
.O6(CLBLM_R_X63Y96_SLICE_X95Y96_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h270027aa275527ff)
  ) CLBLM_R_X63Y96_SLICE_X95Y96_CLUT (
.I0(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I1(CLBLM_L_X62Y98_SLICE_X92Y98_AQ),
.I2(CLBLM_L_X62Y96_SLICE_X93Y96_CQ),
.I3(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I4(CLBLM_L_X64Y96_SLICE_X97Y96_CQ),
.I5(CLBLM_R_X63Y95_SLICE_X95Y95_CQ),
.O5(CLBLM_R_X63Y96_SLICE_X95Y96_CO5),
.O6(CLBLM_R_X63Y96_SLICE_X95Y96_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0fafa0f000a0a)
  ) CLBLM_R_X63Y96_SLICE_X95Y96_BLUT (
.I0(CLBLM_R_X63Y96_SLICE_X94Y96_CO6),
.I1(1'b1),
.I2(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I3(CLBLM_L_X64Y97_SLICE_X96Y97_B5Q),
.I4(CLBLM_L_X56Y98_SLICE_X85Y98_DQ),
.I5(CLBLM_L_X50Y105_SLICE_X77Y105_AQ),
.O5(CLBLM_R_X63Y96_SLICE_X95Y96_BO5),
.O6(CLBLM_R_X63Y96_SLICE_X95Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0e4e4f5a0)
  ) CLBLM_R_X63Y96_SLICE_X95Y96_ALUT (
.I0(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I1(CLBLM_R_X63Y98_SLICE_X95Y98_D5Q),
.I2(CLBLM_L_X50Y107_SLICE_X77Y107_AQ),
.I3(CLBLM_L_X64Y96_SLICE_X96Y96_AO6),
.I4(CLBLM_L_X56Y98_SLICE_X85Y98_DQ),
.I5(1'b1),
.O5(CLBLM_R_X63Y96_SLICE_X95Y96_AO5),
.O6(CLBLM_R_X63Y96_SLICE_X95Y96_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y97_SLICE_X94Y97_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y99_SLICE_X93Y99_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y97_SLICE_X94Y97_CO6),
.Q(CLBLM_R_X63Y97_SLICE_X94Y97_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y97_SLICE_X94Y97_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y99_SLICE_X93Y99_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_L_X62Y97_SLICE_X93Y97_CO6),
.Q(CLBLM_R_X63Y97_SLICE_X94Y97_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y97_SLICE_X94Y97_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X62Y99_SLICE_X93Y99_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y97_SLICE_X94Y97_DO6),
.Q(CLBLM_R_X63Y97_SLICE_X94Y97_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffaa5500)
  ) CLBLM_R_X63Y97_SLICE_X94Y97_DLUT (
.I0(CLBLM_L_X56Y98_SLICE_X85Y98_DQ),
.I1(CLBLM_R_X49Y105_SLICE_X75Y105_CQ),
.I2(1'b1),
.I3(CLBLM_R_X63Y95_SLICE_X94Y95_AO5),
.I4(CLBLM_R_X63Y100_SLICE_X95Y100_AQ),
.I5(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.O5(CLBLM_R_X63Y97_SLICE_X94Y97_DO5),
.O6(CLBLM_R_X63Y97_SLICE_X94Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0f3d1e2c0)
  ) CLBLM_R_X63Y97_SLICE_X94Y97_CLUT (
.I0(CLBLM_L_X56Y98_SLICE_X85Y98_DQ),
.I1(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I2(CLBLM_L_X50Y106_SLICE_X76Y106_AQ),
.I3(CLBLM_R_X63Y98_SLICE_X95Y98_CQ),
.I4(CLBLM_L_X64Y95_SLICE_X96Y95_CO5),
.I5(1'b1),
.O5(CLBLM_R_X63Y97_SLICE_X94Y97_CO5),
.O6(CLBLM_R_X63Y97_SLICE_X94Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44fafa5050)
  ) CLBLM_R_X63Y97_SLICE_X94Y97_BLUT (
.I0(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I1(CLBLM_R_X63Y97_SLICE_X94Y97_BQ),
.I2(CLBLM_R_X63Y95_SLICE_X95Y95_AQ),
.I3(CLBLM_L_X62Y95_SLICE_X92Y95_A5Q),
.I4(CLBLM_L_X64Y97_SLICE_X97Y97_AQ),
.I5(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.O5(CLBLM_R_X63Y97_SLICE_X94Y97_BO5),
.O6(CLBLM_R_X63Y97_SLICE_X94Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffe233e2cce200e2)
  ) CLBLM_R_X63Y97_SLICE_X94Y97_ALUT (
.I0(CLBLM_L_X62Y97_SLICE_X92Y97_CQ),
.I1(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I2(CLBLM_R_X63Y98_SLICE_X94Y98_CQ),
.I3(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I4(CLBLM_L_X62Y97_SLICE_X93Y97_BQ),
.I5(CLBLM_R_X63Y98_SLICE_X95Y98_CQ),
.O5(CLBLM_R_X63Y97_SLICE_X94Y97_AO5),
.O6(CLBLM_R_X63Y97_SLICE_X94Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X63Y97_SLICE_X94Y97_MUXF7A (
.I0(CLBLM_R_X63Y97_SLICE_X94Y97_BO6),
.I1(CLBLM_R_X63Y97_SLICE_X94Y97_AO6),
.O(CLBLM_R_X63Y97_SLICE_X94Y97_F7AMUX_O),
.S(CLBLM_L_X62Y106_SLICE_X93Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y97_SLICE_X95Y97_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_R_X63Y100_SLICE_X94Y100_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y97_SLICE_X95Y97_CO5),
.Q(CLBLM_R_X63Y97_SLICE_X95Y97_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y97_SLICE_X95Y97_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_R_X63Y100_SLICE_X94Y100_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y97_SLICE_X95Y97_DO5),
.Q(CLBLM_R_X63Y97_SLICE_X95Y97_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y97_SLICE_X95Y97_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_R_X63Y100_SLICE_X94Y100_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y97_SLICE_X95Y97_CO6),
.Q(CLBLM_R_X63Y97_SLICE_X95Y97_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y97_SLICE_X95Y97_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_R_X63Y100_SLICE_X94Y100_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y97_SLICE_X95Y97_DO6),
.Q(CLBLM_R_X63Y97_SLICE_X95Y97_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0afa0fcfc0c0c)
  ) CLBLM_R_X63Y97_SLICE_X95Y97_DLUT (
.I0(CLBLM_L_X64Y97_SLICE_X96Y97_AQ),
.I1(CLBLM_R_X49Y106_SLICE_X74Y106_AQ),
.I2(CLBLM_R_X63Y99_SLICE_X94Y99_DO6),
.I3(CLBLM_R_X49Y105_SLICE_X75Y105_CQ),
.I4(CLBLM_L_X64Y97_SLICE_X96Y97_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X63Y97_SLICE_X95Y97_DO5),
.O6(CLBLM_R_X63Y97_SLICE_X95Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaaaaf0f0ff00)
  ) CLBLM_R_X63Y97_SLICE_X95Y97_CLUT (
.I0(CLBLM_L_X50Y104_SLICE_X76Y104_AQ),
.I1(CLBLM_R_X63Y98_SLICE_X95Y98_AQ),
.I2(CLBLM_R_X63Y98_SLICE_X95Y98_A5Q),
.I3(CLBLM_L_X50Y105_SLICE_X77Y105_AQ),
.I4(CLBLM_R_X63Y99_SLICE_X94Y99_DO6),
.I5(1'b1),
.O5(CLBLM_R_X63Y97_SLICE_X95Y97_CO5),
.O6(CLBLM_R_X63Y97_SLICE_X95Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfceefc2230ee3022)
  ) CLBLM_R_X63Y97_SLICE_X95Y97_BLUT (
.I0(CLBLM_R_X63Y95_SLICE_X95Y95_DQ),
.I1(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I2(CLBLM_L_X64Y96_SLICE_X97Y96_AQ),
.I3(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I4(CLBLM_R_X63Y96_SLICE_X95Y96_BQ),
.I5(CLBLM_L_X62Y98_SLICE_X92Y98_CQ),
.O5(CLBLM_R_X63Y97_SLICE_X95Y97_BO5),
.O6(CLBLM_R_X63Y97_SLICE_X95Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7b3d591e6a2c480)
  ) CLBLM_R_X63Y97_SLICE_X95Y97_ALUT (
.I0(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I1(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I2(CLBLM_L_X62Y103_SLICE_X93Y103_AQ),
.I3(CLBLM_R_X63Y99_SLICE_X95Y99_B5Q),
.I4(CLBLM_R_X63Y97_SLICE_X95Y97_C5Q),
.I5(CLBLM_L_X62Y97_SLICE_X92Y97_BQ),
.O5(CLBLM_R_X63Y97_SLICE_X95Y97_AO5),
.O6(CLBLM_R_X63Y97_SLICE_X95Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X63Y97_SLICE_X95Y97_MUXF7A (
.I0(CLBLM_R_X63Y97_SLICE_X95Y97_BO6),
.I1(CLBLM_R_X63Y97_SLICE_X95Y97_AO6),
.O(CLBLM_R_X63Y97_SLICE_X95Y97_F7AMUX_O),
.S(CLBLM_L_X62Y106_SLICE_X93Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y98_SLICE_X94Y98_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_R_X63Y100_SLICE_X94Y100_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y98_SLICE_X94Y98_CO5),
.Q(CLBLM_R_X63Y98_SLICE_X94Y98_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y98_SLICE_X94Y98_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_R_X63Y100_SLICE_X94Y100_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y98_SLICE_X94Y98_CO6),
.Q(CLBLM_R_X63Y98_SLICE_X94Y98_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2202220222002200)
  ) CLBLM_R_X63Y98_SLICE_X94Y98_DLUT (
.I0(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I1(CLBLM_L_X56Y97_SLICE_X85Y97_AQ),
.I2(CLBLM_R_X63Y94_SLICE_X94Y94_AQ),
.I3(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I4(1'b1),
.I5(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.O5(CLBLM_R_X63Y98_SLICE_X94Y98_DO5),
.O6(CLBLM_R_X63Y98_SLICE_X94Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccff00f0f0aaaa)
  ) CLBLM_R_X63Y98_SLICE_X94Y98_CLUT (
.I0(CLBLM_L_X50Y106_SLICE_X76Y106_CQ),
.I1(CLBLM_R_X63Y98_SLICE_X95Y98_BQ),
.I2(CLBLM_R_X63Y98_SLICE_X95Y98_B5Q),
.I3(CLBLM_L_X50Y106_SLICE_X76Y106_AQ),
.I4(CLBLM_R_X63Y99_SLICE_X94Y99_DO6),
.I5(1'b1),
.O5(CLBLM_R_X63Y98_SLICE_X94Y98_CO5),
.O6(CLBLM_R_X63Y98_SLICE_X94Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfedc7654ba983210)
  ) CLBLM_R_X63Y98_SLICE_X94Y98_BLUT (
.I0(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I1(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I2(CLBLM_R_X63Y94_SLICE_X95Y94_AQ),
.I3(CLBLM_L_X64Y96_SLICE_X97Y96_DQ),
.I4(CLBLM_L_X62Y95_SLICE_X92Y95_AQ),
.I5(CLBLM_L_X62Y96_SLICE_X93Y96_DQ),
.O5(CLBLM_R_X63Y98_SLICE_X94Y98_BO5),
.O6(CLBLM_R_X63Y98_SLICE_X94Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdb97531eca86420)
  ) CLBLM_R_X63Y98_SLICE_X94Y98_ALUT (
.I0(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I1(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I2(CLBLM_R_X63Y97_SLICE_X95Y97_CQ),
.I3(CLBLM_R_X63Y99_SLICE_X95Y99_BQ),
.I4(CLBLM_L_X64Y109_SLICE_X96Y109_AQ),
.I5(CLBLM_L_X62Y97_SLICE_X92Y97_AQ),
.O5(CLBLM_R_X63Y98_SLICE_X94Y98_AO5),
.O6(CLBLM_R_X63Y98_SLICE_X94Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X63Y98_SLICE_X94Y98_MUXF7A (
.I0(CLBLM_R_X63Y98_SLICE_X94Y98_BO6),
.I1(CLBLM_R_X63Y98_SLICE_X94Y98_AO6),
.O(CLBLM_R_X63Y98_SLICE_X94Y98_F7AMUX_O),
.S(CLBLM_L_X62Y106_SLICE_X93Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X63Y98_SLICE_X95Y98_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y98_SLICE_X95Y98_AO5),
.Q(CLBLM_R_X63Y98_SLICE_X95Y98_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X63Y98_SLICE_X95Y98_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y98_SLICE_X95Y98_BO5),
.Q(CLBLM_R_X63Y98_SLICE_X95Y98_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X63Y98_SLICE_X95Y98_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y98_SLICE_X95Y98_CO5),
.Q(CLBLM_R_X63Y98_SLICE_X95Y98_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X63Y98_SLICE_X95Y98_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y98_SLICE_X95Y98_DO5),
.Q(CLBLM_R_X63Y98_SLICE_X95Y98_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X63Y98_SLICE_X95Y98_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y98_SLICE_X95Y98_AO6),
.Q(CLBLM_R_X63Y98_SLICE_X95Y98_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X63Y98_SLICE_X95Y98_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y98_SLICE_X95Y98_BO6),
.Q(CLBLM_R_X63Y98_SLICE_X95Y98_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X63Y98_SLICE_X95Y98_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y98_SLICE_X95Y98_CO6),
.Q(CLBLM_R_X63Y98_SLICE_X95Y98_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X63Y98_SLICE_X95Y98_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y98_SLICE_X95Y98_DO6),
.Q(CLBLM_R_X63Y98_SLICE_X95Y98_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaf0ffcc00cc)
  ) CLBLM_R_X63Y98_SLICE_X95Y98_DLUT (
.I0(CLBLM_L_X50Y107_SLICE_X76Y107_BQ),
.I1(CLBLM_L_X64Y99_SLICE_X96Y99_BQ),
.I2(CLBLM_R_X65Y101_SLICE_X99Y101_AQ),
.I3(CLBLM_R_X63Y99_SLICE_X94Y99_DO5),
.I4(CLBLM_L_X50Y107_SLICE_X77Y107_AQ),
.I5(1'b1),
.O5(CLBLM_R_X63Y98_SLICE_X95Y98_DO5),
.O6(CLBLM_R_X63Y98_SLICE_X95Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0f0aaaaff00)
  ) CLBLM_R_X63Y98_SLICE_X95Y98_CLUT (
.I0(CLBLM_L_X50Y106_SLICE_X76Y106_CQ),
.I1(CLBLM_L_X50Y106_SLICE_X76Y106_AQ),
.I2(CLBLM_L_X64Y99_SLICE_X97Y99_AQ),
.I3(CLBLM_R_X65Y98_SLICE_X99Y98_AQ),
.I4(CLBLM_R_X63Y99_SLICE_X94Y99_DO5),
.I5(1'b1),
.O5(CLBLM_R_X63Y98_SLICE_X95Y98_CO5),
.O6(CLBLM_R_X63Y98_SLICE_X95Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88f5f5a0a0)
  ) CLBLM_R_X63Y98_SLICE_X95Y98_BLUT (
.I0(CLBLM_R_X63Y99_SLICE_X94Y99_DO5),
.I1(CLBLM_R_X63Y98_SLICE_X94Y98_CQ),
.I2(CLBLM_R_X63Y98_SLICE_X94Y98_C5Q),
.I3(CLBLM_R_X65Y98_SLICE_X98Y98_AQ),
.I4(CLBLM_R_X65Y104_SLICE_X99Y104_AQ),
.I5(1'b1),
.O5(CLBLM_R_X63Y98_SLICE_X95Y98_BO5),
.O6(CLBLM_R_X63Y98_SLICE_X95Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50fa50eeee4444)
  ) CLBLM_R_X63Y98_SLICE_X95Y98_ALUT (
.I0(CLBLM_R_X63Y99_SLICE_X94Y99_DO5),
.I1(CLBLM_L_X64Y98_SLICE_X96Y98_AQ),
.I2(CLBLM_L_X64Y98_SLICE_X97Y98_AQ),
.I3(CLBLM_R_X63Y97_SLICE_X95Y97_CQ),
.I4(CLBLM_R_X63Y97_SLICE_X95Y97_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X63Y98_SLICE_X95Y98_AO5),
.O6(CLBLM_R_X63Y98_SLICE_X95Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y99_SLICE_X94Y99_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_R_X63Y100_SLICE_X94Y100_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y99_SLICE_X94Y99_CO5),
.Q(CLBLM_R_X63Y99_SLICE_X94Y99_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y99_SLICE_X94Y99_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_R_X63Y100_SLICE_X94Y100_BO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y99_SLICE_X94Y99_CO6),
.Q(CLBLM_R_X63Y99_SLICE_X94Y99_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff7f00400000)
  ) CLBLM_R_X63Y99_SLICE_X94Y99_DLUT (
.I0(CLBLM_L_X62Y104_SLICE_X93Y104_AQ),
.I1(CLBLM_L_X60Y98_SLICE_X90Y98_BQ),
.I2(CLBLM_R_X59Y102_SLICE_X89Y102_AQ),
.I3(CLBLM_L_X62Y102_SLICE_X93Y102_AO5),
.I4(CLBLM_R_X59Y102_SLICE_X88Y102_AQ),
.I5(1'b1),
.O5(CLBLM_R_X63Y99_SLICE_X94Y99_DO5),
.O6(CLBLM_R_X63Y99_SLICE_X94Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0f0ccccff00)
  ) CLBLM_R_X63Y99_SLICE_X94Y99_CLUT (
.I0(CLBLM_R_X63Y99_SLICE_X95Y99_AQ),
.I1(CLBLM_R_X63Y99_SLICE_X95Y99_A5Q),
.I2(CLBLM_L_X50Y107_SLICE_X76Y107_BQ),
.I3(CLBLM_L_X50Y107_SLICE_X77Y107_AQ),
.I4(CLBLM_R_X63Y99_SLICE_X94Y99_DO6),
.I5(1'b1),
.O5(CLBLM_R_X63Y99_SLICE_X94Y99_CO5),
.O6(CLBLM_R_X63Y99_SLICE_X94Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5ee44a0a0ee44)
  ) CLBLM_R_X63Y99_SLICE_X94Y99_BLUT (
.I0(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I1(CLBLM_R_X63Y95_SLICE_X95Y95_BQ),
.I2(CLBLM_L_X62Y98_SLICE_X92Y98_DQ),
.I3(CLBLM_L_X64Y96_SLICE_X97Y96_BQ),
.I4(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I5(CLBLM_R_X63Y97_SLICE_X94Y97_DQ),
.O5(CLBLM_R_X63Y99_SLICE_X94Y99_BO5),
.O6(CLBLM_R_X63Y99_SLICE_X94Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddfadd5088fa8850)
  ) CLBLM_R_X63Y99_SLICE_X94Y99_ALUT (
.I0(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I1(CLBLM_R_X63Y105_SLICE_X94Y105_AQ),
.I2(CLBLM_L_X62Y100_SLICE_X93Y100_AQ),
.I3(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I4(CLBLM_R_X63Y97_SLICE_X95Y97_DQ),
.I5(CLBLM_R_X63Y99_SLICE_X95Y99_CQ),
.O5(CLBLM_R_X63Y99_SLICE_X94Y99_AO5),
.O6(CLBLM_R_X63Y99_SLICE_X94Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X63Y99_SLICE_X94Y99_MUXF7A (
.I0(CLBLM_R_X63Y99_SLICE_X94Y99_BO6),
.I1(CLBLM_R_X63Y99_SLICE_X94Y99_AO6),
.O(CLBLM_R_X63Y99_SLICE_X94Y99_F7AMUX_O),
.S(CLBLM_L_X62Y106_SLICE_X93Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X63Y99_SLICE_X95Y99_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y99_SLICE_X95Y99_AO5),
.Q(CLBLM_R_X63Y99_SLICE_X95Y99_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X63Y99_SLICE_X95Y99_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y99_SLICE_X95Y99_BO5),
.Q(CLBLM_R_X63Y99_SLICE_X95Y99_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X63Y99_SLICE_X95Y99_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y99_SLICE_X95Y99_CO5),
.Q(CLBLM_R_X63Y99_SLICE_X95Y99_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X63Y99_SLICE_X95Y99_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y99_SLICE_X95Y99_AO6),
.Q(CLBLM_R_X63Y99_SLICE_X95Y99_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X63Y99_SLICE_X95Y99_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y99_SLICE_X95Y99_BO6),
.Q(CLBLM_R_X63Y99_SLICE_X95Y99_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X63Y99_SLICE_X95Y99_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y99_SLICE_X95Y99_CO6),
.Q(CLBLM_R_X63Y99_SLICE_X95Y99_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y99_SLICE_X95Y99_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y99_SLICE_X95Y99_DO5),
.O6(CLBLM_R_X63Y99_SLICE_X95Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ff000cacacaca)
  ) CLBLM_R_X63Y99_SLICE_X95Y99_CLUT (
.I0(CLBLM_R_X65Y99_SLICE_X98Y99_AQ),
.I1(CLBLM_R_X49Y106_SLICE_X74Y106_AQ),
.I2(CLBLM_R_X63Y99_SLICE_X94Y99_DO5),
.I3(CLBLM_R_X49Y105_SLICE_X75Y105_CQ),
.I4(CLBLM_R_X65Y99_SLICE_X99Y99_AQ),
.I5(1'b1),
.O5(CLBLM_R_X63Y99_SLICE_X95Y99_CO5),
.O6(CLBLM_R_X63Y99_SLICE_X95Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0bbbb8888)
  ) CLBLM_R_X63Y99_SLICE_X95Y99_BLUT (
.I0(CLBLM_L_X50Y105_SLICE_X77Y105_AQ),
.I1(CLBLM_R_X63Y99_SLICE_X94Y99_DO5),
.I2(CLBLM_L_X50Y104_SLICE_X76Y104_AQ),
.I3(1'b1),
.I4(CLBLM_R_X65Y98_SLICE_X98Y98_BQ),
.I5(1'b1),
.O5(CLBLM_R_X63Y99_SLICE_X95Y99_BO5),
.O6(CLBLM_R_X63Y99_SLICE_X95Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee2222f3c0f3c0)
  ) CLBLM_R_X63Y99_SLICE_X95Y99_ALUT (
.I0(CLBLM_R_X65Y105_SLICE_X98Y105_AQ),
.I1(CLBLM_R_X63Y99_SLICE_X94Y99_DO5),
.I2(CLBLM_R_X63Y99_SLICE_X94Y99_C5Q),
.I3(CLBLM_R_X65Y103_SLICE_X99Y103_AQ),
.I4(CLBLM_R_X63Y99_SLICE_X94Y99_CQ),
.I5(1'b1),
.O5(CLBLM_R_X63Y99_SLICE_X95Y99_AO5),
.O6(CLBLM_R_X63Y99_SLICE_X95Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y100_SLICE_X94Y100_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLM_R_X63Y100_SLICE_X94Y100_AO6),
.PRE(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.Q(CLBLM_R_X63Y100_SLICE_X94Y100_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000ff000000ff)
  ) CLBLM_R_X63Y100_SLICE_X94Y100_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X62Y104_SLICE_X93Y104_AQ),
.I4(CLBLM_R_X59Y102_SLICE_X89Y102_AQ),
.I5(1'b1),
.O5(CLBLM_R_X63Y100_SLICE_X94Y100_DO5),
.O6(CLBLM_R_X63Y100_SLICE_X94Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000400cccccccc)
  ) CLBLM_R_X63Y100_SLICE_X94Y100_CLUT (
.I0(CLBLM_L_X60Y99_SLICE_X91Y99_AO6),
.I1(CLBLM_L_X62Y99_SLICE_X92Y99_AO6),
.I2(CLBLM_R_X59Y102_SLICE_X89Y102_AQ),
.I3(CLBLM_L_X62Y104_SLICE_X93Y104_AQ),
.I4(CLBLM_L_X60Y99_SLICE_X91Y99_BO6),
.I5(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.O5(CLBLM_R_X63Y100_SLICE_X94Y100_CO5),
.O6(CLBLM_R_X63Y100_SLICE_X94Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0400000000004000)
  ) CLBLM_R_X63Y100_SLICE_X94Y100_BLUT (
.I0(CLBLM_L_X62Y102_SLICE_X93Y102_AO5),
.I1(CLBLM_R_X59Y102_SLICE_X89Y102_AQ),
.I2(CLBLM_R_X59Y102_SLICE_X88Y102_AQ),
.I3(CLBLM_L_X56Y103_SLICE_X85Y103_CO6),
.I4(CLBLM_L_X60Y98_SLICE_X90Y98_BQ),
.I5(CLBLM_L_X62Y104_SLICE_X93Y104_AQ),
.O5(CLBLM_R_X63Y100_SLICE_X94Y100_BO5),
.O6(CLBLM_R_X63Y100_SLICE_X94Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f2d0f0f0f0f0)
  ) CLBLM_R_X63Y100_SLICE_X94Y100_ALUT (
.I0(CLBLM_R_X63Y100_SLICE_X94Y100_DO6),
.I1(CLBLM_L_X60Y100_SLICE_X91Y100_CO6),
.I2(CLBLM_R_X63Y100_SLICE_X94Y100_AQ),
.I3(CLBLM_L_X50Y104_SLICE_X76Y104_AQ),
.I4(CLBLM_L_X60Y99_SLICE_X91Y99_AO6),
.I5(CLBLM_L_X56Y103_SLICE_X85Y103_CO6),
.O5(CLBLM_R_X63Y100_SLICE_X94Y100_AO5),
.O6(CLBLM_R_X63Y100_SLICE_X94Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X63Y100_SLICE_X95Y100_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y100_SLICE_X95Y100_AO5),
.Q(CLBLM_R_X63Y100_SLICE_X95Y100_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X63Y100_SLICE_X95Y100_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_DQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y100_SLICE_X95Y100_AO6),
.Q(CLBLM_R_X63Y100_SLICE_X95Y100_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y100_SLICE_X95Y100_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y100_SLICE_X95Y100_DO5),
.O6(CLBLM_R_X63Y100_SLICE_X95Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h303f303f303f303f)
  ) CLBLM_R_X63Y100_SLICE_X95Y100_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X63Y97_SLICE_X95Y97_D5Q),
.I2(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I3(CLBLM_L_X62Y100_SLICE_X93Y100_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y100_SLICE_X95Y100_CO5),
.O6(CLBLM_R_X63Y100_SLICE_X95Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3ffff33f33fff)
  ) CLBLM_R_X63Y100_SLICE_X95Y100_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I2(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I3(CLBLM_L_X62Y100_SLICE_X92Y100_CQ),
.I4(CLBLM_L_X64Y100_SLICE_X97Y100_D_XOR),
.I5(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.O5(CLBLM_R_X63Y100_SLICE_X95Y100_BO5),
.O6(CLBLM_R_X63Y100_SLICE_X95Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cfc0afafa0a0)
  ) CLBLM_R_X63Y100_SLICE_X95Y100_ALUT (
.I0(CLBLM_L_X62Y100_SLICE_X93Y100_BQ),
.I1(CLBLM_L_X62Y100_SLICE_X93Y100_AQ),
.I2(CLBLM_R_X63Y99_SLICE_X94Y99_DO5),
.I3(CLBLM_R_X65Y105_SLICE_X98Y105_BQ),
.I4(CLBLM_R_X65Y105_SLICE_X99Y105_AQ),
.I5(1'b1),
.O5(CLBLM_R_X63Y100_SLICE_X95Y100_AO5),
.O6(CLBLM_R_X63Y100_SLICE_X95Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y101_SLICE_X94Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y101_SLICE_X94Y101_DO5),
.O6(CLBLM_R_X63Y101_SLICE_X94Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y101_SLICE_X94Y101_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y101_SLICE_X94Y101_CO5),
.O6(CLBLM_R_X63Y101_SLICE_X94Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y101_SLICE_X94Y101_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y101_SLICE_X94Y101_BO5),
.O6(CLBLM_R_X63Y101_SLICE_X94Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y101_SLICE_X94Y101_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y101_SLICE_X94Y101_AO5),
.O6(CLBLM_R_X63Y101_SLICE_X94Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X63Y101_SLICE_X95Y101_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y105_SLICE_X93Y105_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y101_SLICE_X95Y101_AO6),
.Q(CLBLM_R_X63Y101_SLICE_X95Y101_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffddddff55ff55)
  ) CLBLM_R_X63Y101_SLICE_X95Y101_DLUT (
.I0(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I1(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I2(1'b1),
.I3(CLBLM_L_X64Y102_SLICE_X97Y102_A_XOR),
.I4(CLBLM_R_X49Y104_SLICE_X74Y104_AQ),
.I5(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.O5(CLBLM_R_X63Y101_SLICE_X95Y101_DO5),
.O6(CLBLM_R_X63Y101_SLICE_X95Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffddffddffff5555)
  ) CLBLM_R_X63Y101_SLICE_X95Y101_CLUT (
.I0(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I1(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I2(1'b1),
.I3(CLBLM_R_X49Y104_SLICE_X75Y104_BQ),
.I4(CLBLM_L_X64Y102_SLICE_X97Y102_C_XOR),
.I5(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.O5(CLBLM_R_X63Y101_SLICE_X95Y101_CO5),
.O6(CLBLM_R_X63Y101_SLICE_X95Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88c0bbf300000000)
  ) CLBLM_R_X63Y101_SLICE_X95Y101_BLUT (
.I0(CLBLM_L_X64Y109_SLICE_X96Y109_A5Q),
.I1(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I2(CLBLM_R_X63Y99_SLICE_X95Y99_C5Q),
.I3(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.I4(CLBLM_R_X63Y100_SLICE_X95Y100_CO6),
.I5(CLBLM_L_X62Y106_SLICE_X93Y106_CO6),
.O5(CLBLM_R_X63Y101_SLICE_X95Y101_BO5),
.O6(CLBLM_R_X63Y101_SLICE_X95Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf555a00055f500a0)
  ) CLBLM_R_X63Y101_SLICE_X95Y101_ALUT (
.I0(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I1(1'b1),
.I2(CLBLM_L_X64Y98_SLICE_X97Y98_AQ),
.I3(CLBLL_R_X57Y103_SLICE_X86Y103_AQ),
.I4(CLBLM_L_X64Y107_SLICE_X97Y107_BQ),
.I5(CLBLL_R_X57Y103_SLICE_X86Y103_A5Q),
.O5(CLBLM_R_X63Y101_SLICE_X95Y101_AO5),
.O6(CLBLM_R_X63Y101_SLICE_X95Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y102_SLICE_X94Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y102_SLICE_X94Y102_DO5),
.O6(CLBLM_R_X63Y102_SLICE_X94Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y102_SLICE_X94Y102_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y102_SLICE_X94Y102_CO5),
.O6(CLBLM_R_X63Y102_SLICE_X94Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y102_SLICE_X94Y102_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y102_SLICE_X94Y102_BO5),
.O6(CLBLM_R_X63Y102_SLICE_X94Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y102_SLICE_X94Y102_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y102_SLICE_X94Y102_AO5),
.O6(CLBLM_R_X63Y102_SLICE_X94Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y102_SLICE_X95Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y102_SLICE_X95Y102_DO5),
.O6(CLBLM_R_X63Y102_SLICE_X95Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y102_SLICE_X95Y102_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y102_SLICE_X95Y102_CO5),
.O6(CLBLM_R_X63Y102_SLICE_X95Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y102_SLICE_X95Y102_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y102_SLICE_X95Y102_BO5),
.O6(CLBLM_R_X63Y102_SLICE_X95Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbfffbff3b3f3b3)
  ) CLBLM_R_X63Y102_SLICE_X95Y102_ALUT (
.I0(CLBLM_R_X49Y104_SLICE_X75Y104_AQ),
.I1(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I2(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I3(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I4(1'b1),
.I5(CLBLM_L_X64Y102_SLICE_X97Y102_B_XOR),
.O5(CLBLM_R_X63Y102_SLICE_X95Y102_AO5),
.O6(CLBLM_R_X63Y102_SLICE_X95Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y103_SLICE_X94Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y103_SLICE_X94Y103_DO5),
.O6(CLBLM_R_X63Y103_SLICE_X94Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y103_SLICE_X94Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y103_SLICE_X94Y103_CO5),
.O6(CLBLM_R_X63Y103_SLICE_X94Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y103_SLICE_X94Y103_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y103_SLICE_X94Y103_BO5),
.O6(CLBLM_R_X63Y103_SLICE_X94Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0000cfc0cfc0)
  ) CLBLM_R_X63Y103_SLICE_X94Y103_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X49Y107_SLICE_X74Y107_AQ),
.I2(CLBLM_L_X62Y107_SLICE_X93Y107_BO6),
.I3(CLBLM_L_X64Y107_SLICE_X96Y107_AQ),
.I4(CLBLM_R_X63Y104_SLICE_X94Y104_AQ),
.I5(CLBLM_L_X62Y107_SLICE_X93Y107_AO6),
.O5(CLBLM_R_X63Y103_SLICE_X94Y103_AO5),
.O6(CLBLM_R_X63Y103_SLICE_X94Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X63Y103_SLICE_X95Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y105_SLICE_X93Y105_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y103_SLICE_X95Y103_AO6),
.Q(CLBLM_R_X63Y103_SLICE_X95Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X63Y103_SLICE_X95Y103_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y105_SLICE_X93Y105_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y103_SLICE_X95Y103_BO6),
.Q(CLBLM_R_X63Y103_SLICE_X95Y103_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X63Y103_SLICE_X95Y103_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y105_SLICE_X93Y105_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y103_SLICE_X95Y103_CO6),
.Q(CLBLM_R_X63Y103_SLICE_X95Y103_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffcfcfafafcfcf)
  ) CLBLM_R_X63Y103_SLICE_X95Y103_DLUT (
.I0(CLBLM_R_X49Y107_SLICE_X75Y107_CQ),
.I1(CLBLM_L_X64Y103_SLICE_X97Y103_D_XOR),
.I2(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I3(1'b1),
.I4(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I5(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.O5(CLBLM_R_X63Y103_SLICE_X95Y103_DO5),
.O6(CLBLM_R_X63Y103_SLICE_X95Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9090ffff90900000)
  ) CLBLM_R_X63Y103_SLICE_X95Y103_CLUT (
.I0(CLBLL_R_X57Y103_SLICE_X86Y103_AQ),
.I1(CLBLL_R_X57Y103_SLICE_X86Y103_A5Q),
.I2(CLBLM_L_X64Y98_SLICE_X96Y98_AQ),
.I3(1'b1),
.I4(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I5(CLBLM_L_X64Y107_SLICE_X96Y107_AQ),
.O5(CLBLM_R_X63Y103_SLICE_X95Y103_CO5),
.O6(CLBLM_R_X63Y103_SLICE_X95Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a055005500f5a0)
  ) CLBLM_R_X63Y103_SLICE_X95Y103_BLUT (
.I0(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I1(1'b1),
.I2(CLBLM_L_X64Y99_SLICE_X96Y99_BQ),
.I3(CLBLM_L_X64Y106_SLICE_X96Y106_BQ),
.I4(CLBLL_R_X57Y103_SLICE_X86Y103_AQ),
.I5(CLBLL_R_X57Y103_SLICE_X86Y103_A5Q),
.O5(CLBLM_R_X63Y103_SLICE_X95Y103_BO5),
.O6(CLBLM_R_X63Y103_SLICE_X95Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d850505050d8d8)
  ) CLBLM_R_X63Y103_SLICE_X95Y103_ALUT (
.I0(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I1(CLBLM_R_X65Y103_SLICE_X99Y103_BQ),
.I2(CLBLM_L_X64Y109_SLICE_X96Y109_AQ),
.I3(1'b1),
.I4(CLBLL_R_X57Y103_SLICE_X86Y103_AQ),
.I5(CLBLL_R_X57Y103_SLICE_X86Y103_A5Q),
.O5(CLBLM_R_X63Y103_SLICE_X95Y103_AO5),
.O6(CLBLM_R_X63Y103_SLICE_X95Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y104_SLICE_X94Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y100_SLICE_X92Y100_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y104_SLICE_X94Y104_AO6),
.Q(CLBLM_R_X63Y104_SLICE_X94Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y104_SLICE_X94Y104_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y100_SLICE_X92Y100_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y104_SLICE_X94Y104_BO6),
.Q(CLBLM_R_X63Y104_SLICE_X94Y104_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0bb88f0f00000)
  ) CLBLM_R_X63Y104_SLICE_X94Y104_DLUT (
.I0(CLBLM_R_X63Y105_SLICE_X95Y105_D_XOR),
.I1(CLBLM_L_X62Y105_SLICE_X93Y105_AO6),
.I2(CLBLM_L_X50Y106_SLICE_X76Y106_AQ),
.I3(CLBLM_R_X63Y106_SLICE_X94Y106_A_XOR),
.I4(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I5(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.O5(CLBLM_R_X63Y104_SLICE_X94Y104_DO5),
.O6(CLBLM_R_X63Y104_SLICE_X94Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5b1e4a0a0a0a0a0)
  ) CLBLM_R_X63Y104_SLICE_X94Y104_CLUT (
.I0(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I1(CLBLM_L_X62Y105_SLICE_X93Y105_AO6),
.I2(CLBLM_L_X50Y105_SLICE_X77Y105_AQ),
.I3(CLBLM_R_X63Y105_SLICE_X95Y105_A_XOR),
.I4(CLBLM_R_X63Y105_SLICE_X94Y105_B_XOR),
.I5(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.O5(CLBLM_R_X63Y104_SLICE_X94Y104_CO5),
.O6(CLBLM_R_X63Y104_SLICE_X94Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaafaaaaaaaee)
  ) CLBLM_R_X63Y104_SLICE_X94Y104_BLUT (
.I0(CLBLM_R_X63Y104_SLICE_X94Y104_DO6),
.I1(CLBLM_R_X63Y104_SLICE_X94Y104_BQ),
.I2(CLBLM_R_X63Y105_SLICE_X95Y105_D_XOR),
.I3(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I4(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I5(CLBLM_L_X62Y105_SLICE_X92Y105_BO5),
.O5(CLBLM_R_X63Y104_SLICE_X94Y104_BO5),
.O6(CLBLM_R_X63Y104_SLICE_X94Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0054ffff0010)
  ) CLBLM_R_X63Y104_SLICE_X94Y104_ALUT (
.I0(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I1(CLBLM_L_X62Y105_SLICE_X92Y105_BO5),
.I2(CLBLM_R_X63Y104_SLICE_X94Y104_AQ),
.I3(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I4(CLBLM_R_X63Y104_SLICE_X94Y104_CO6),
.I5(CLBLM_R_X63Y105_SLICE_X95Y105_A_XOR),
.O5(CLBLM_R_X63Y104_SLICE_X94Y104_AO5),
.O6(CLBLM_R_X63Y104_SLICE_X94Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y104_SLICE_X95Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y104_SLICE_X95Y104_DO5),
.O6(CLBLM_R_X63Y104_SLICE_X95Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y104_SLICE_X95Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y104_SLICE_X95Y104_CO5),
.O6(CLBLM_R_X63Y104_SLICE_X95Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y104_SLICE_X95Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y104_SLICE_X95Y104_BO5),
.O6(CLBLM_R_X63Y104_SLICE_X95Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hefefef2fefefef2f)
  ) CLBLM_R_X63Y104_SLICE_X95Y104_ALUT (
.I0(CLBLM_L_X64Y104_SLICE_X97Y104_A_XOR),
.I1(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I2(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I3(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I4(CLBLM_R_X49Y108_SLICE_X75Y108_DQ),
.I5(1'b1),
.O5(CLBLM_R_X63Y104_SLICE_X95Y104_AO5),
.O6(CLBLM_R_X63Y104_SLICE_X95Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y105_SLICE_X94Y105_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y100_SLICE_X92Y100_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y105_SLICE_X94Y105_AO5),
.Q(CLBLM_R_X63Y105_SLICE_X94Y105_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X63Y105_SLICE_X94Y105_CARRY4 (
.CI(1'b0),
.CO({CLBLM_R_X63Y105_SLICE_X94Y105_D_CY, CLBLM_R_X63Y105_SLICE_X94Y105_C_CY, CLBLM_R_X63Y105_SLICE_X94Y105_B_CY, CLBLM_R_X63Y105_SLICE_X94Y105_A_CY}),
.CYINIT(1'b1),
.DI({CLBLM_L_X64Y105_SLICE_X97Y105_AQ, CLBLM_L_X64Y105_SLICE_X96Y105_AQ, CLBLM_R_X63Y104_SLICE_X94Y104_AQ, CLBLM_L_X62Y105_SLICE_X92Y105_CQ}),
.O({CLBLM_R_X63Y105_SLICE_X94Y105_D_XOR, CLBLM_R_X63Y105_SLICE_X94Y105_C_XOR, CLBLM_R_X63Y105_SLICE_X94Y105_B_XOR, CLBLM_R_X63Y105_SLICE_X94Y105_A_XOR}),
.S({CLBLM_R_X63Y105_SLICE_X94Y105_DO6, CLBLM_R_X63Y105_SLICE_X94Y105_CO6, CLBLM_R_X63Y105_SLICE_X94Y105_BO6, CLBLM_R_X63Y105_SLICE_X94Y105_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333333333333)
  ) CLBLM_R_X63Y105_SLICE_X94Y105_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X64Y105_SLICE_X97Y105_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y105_SLICE_X94Y105_DO5),
.O6(CLBLM_R_X63Y105_SLICE_X94Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffff0000ffff)
  ) CLBLM_R_X63Y105_SLICE_X94Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X64Y105_SLICE_X96Y105_AQ),
.I5(1'b1),
.O5(CLBLM_R_X63Y105_SLICE_X94Y105_CO5),
.O6(CLBLM_R_X63Y105_SLICE_X94Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0f0f0f)
  ) CLBLM_R_X63Y105_SLICE_X94Y105_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X63Y104_SLICE_X94Y104_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y105_SLICE_X94Y105_BO5),
.O6(CLBLM_R_X63Y105_SLICE_X94Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c333333aaaaaaaa)
  ) CLBLM_R_X63Y105_SLICE_X94Y105_ALUT (
.I0(CLBLM_L_X62Y105_SLICE_X92Y105_AO5),
.I1(CLBLM_L_X62Y105_SLICE_X92Y105_CQ),
.I2(CLBLM_R_X59Y101_SLICE_X89Y101_AQ),
.I3(CLBLM_R_X59Y103_SLICE_X89Y103_A5Q),
.I4(CLBLL_R_X57Y102_SLICE_X86Y102_AQ),
.I5(1'b1),
.O5(CLBLM_R_X63Y105_SLICE_X94Y105_AO5),
.O6(CLBLM_R_X63Y105_SLICE_X94Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X63Y105_SLICE_X95Y105_CARRY4 (
.CI(1'b0),
.CO({CLBLM_R_X63Y105_SLICE_X95Y105_D_CY, CLBLM_R_X63Y105_SLICE_X95Y105_C_CY, CLBLM_R_X63Y105_SLICE_X95Y105_B_CY, CLBLM_R_X63Y105_SLICE_X95Y105_A_CY}),
.CYINIT(CLBLM_L_X62Y105_SLICE_X92Y105_CQ),
.DI({1'b0, 1'b0, 1'b0, CLBLM_R_X63Y105_SLICE_X95Y105_AO5}),
.O({CLBLM_R_X63Y105_SLICE_X95Y105_D_XOR, CLBLM_R_X63Y105_SLICE_X95Y105_C_XOR, CLBLM_R_X63Y105_SLICE_X95Y105_B_XOR, CLBLM_R_X63Y105_SLICE_X95Y105_A_XOR}),
.S({CLBLM_R_X63Y105_SLICE_X95Y105_DO6, CLBLM_R_X63Y105_SLICE_X95Y105_CO6, CLBLM_R_X63Y105_SLICE_X95Y105_BO6, CLBLM_R_X63Y105_SLICE_X95Y105_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X63Y105_SLICE_X95Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X63Y104_SLICE_X94Y104_BQ),
.O5(CLBLM_R_X63Y105_SLICE_X95Y105_DO5),
.O6(CLBLM_R_X63Y105_SLICE_X95Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X63Y105_SLICE_X95Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X64Y105_SLICE_X97Y105_AQ),
.O5(CLBLM_R_X63Y105_SLICE_X95Y105_CO5),
.O6(CLBLM_R_X63Y105_SLICE_X95Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X63Y105_SLICE_X95Y105_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X64Y105_SLICE_X96Y105_AQ),
.O5(CLBLM_R_X63Y105_SLICE_X95Y105_BO5),
.O6(CLBLM_R_X63Y105_SLICE_X95Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000000000)
  ) CLBLM_R_X63Y105_SLICE_X95Y105_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X63Y104_SLICE_X94Y104_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y105_SLICE_X95Y105_AO5),
.O6(CLBLM_R_X63Y105_SLICE_X95Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X63Y106_SLICE_X94Y106_CARRY4 (
.CI(CLBLM_R_X63Y105_SLICE_X94Y105_COUT),
.CO({CLBLM_R_X63Y106_SLICE_X94Y106_D_CY, CLBLM_R_X63Y106_SLICE_X94Y106_C_CY, CLBLM_R_X63Y106_SLICE_X94Y106_B_CY, CLBLM_R_X63Y106_SLICE_X94Y106_A_CY}),
.CYINIT(1'b0),
.DI({CLBLM_L_X64Y106_SLICE_X96Y106_BQ, CLBLM_L_X64Y106_SLICE_X96Y106_AQ, CLBLM_L_X62Y105_SLICE_X93Y105_BQ, CLBLM_R_X63Y104_SLICE_X94Y104_BQ}),
.O({CLBLM_R_X63Y106_SLICE_X94Y106_D_XOR, CLBLM_R_X63Y106_SLICE_X94Y106_C_XOR, CLBLM_R_X63Y106_SLICE_X94Y106_B_XOR, CLBLM_R_X63Y106_SLICE_X94Y106_A_XOR}),
.S({CLBLM_R_X63Y106_SLICE_X94Y106_DO6, CLBLM_R_X63Y106_SLICE_X94Y106_CO6, CLBLM_R_X63Y106_SLICE_X94Y106_BO6, CLBLM_R_X63Y106_SLICE_X94Y106_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555555)
  ) CLBLM_R_X63Y106_SLICE_X94Y106_DLUT (
.I0(CLBLM_L_X64Y106_SLICE_X96Y106_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y106_SLICE_X94Y106_DO5),
.O6(CLBLM_R_X63Y106_SLICE_X94Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333333333333)
  ) CLBLM_R_X63Y106_SLICE_X94Y106_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X64Y106_SLICE_X96Y106_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y106_SLICE_X94Y106_CO5),
.O6(CLBLM_R_X63Y106_SLICE_X94Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333333333333)
  ) CLBLM_R_X63Y106_SLICE_X94Y106_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X62Y105_SLICE_X93Y105_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y106_SLICE_X94Y106_BO5),
.O6(CLBLM_R_X63Y106_SLICE_X94Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffff0000ffff)
  ) CLBLM_R_X63Y106_SLICE_X94Y106_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X63Y104_SLICE_X94Y104_BQ),
.I5(1'b1),
.O5(CLBLM_R_X63Y106_SLICE_X94Y106_AO5),
.O6(CLBLM_R_X63Y106_SLICE_X94Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X63Y106_SLICE_X95Y106_CARRY4 (
.CI(CLBLM_R_X63Y105_SLICE_X95Y105_COUT),
.CO({CLBLM_R_X63Y106_SLICE_X95Y106_D_CY, CLBLM_R_X63Y106_SLICE_X95Y106_C_CY, CLBLM_R_X63Y106_SLICE_X95Y106_B_CY, CLBLM_R_X63Y106_SLICE_X95Y106_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X63Y106_SLICE_X95Y106_D_XOR, CLBLM_R_X63Y106_SLICE_X95Y106_C_XOR, CLBLM_R_X63Y106_SLICE_X95Y106_B_XOR, CLBLM_R_X63Y106_SLICE_X95Y106_A_XOR}),
.S({CLBLM_R_X63Y106_SLICE_X95Y106_DO6, CLBLM_R_X63Y106_SLICE_X95Y106_CO6, CLBLM_R_X63Y106_SLICE_X95Y106_BO6, CLBLM_R_X63Y106_SLICE_X95Y106_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X63Y106_SLICE_X95Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X64Y107_SLICE_X97Y107_BQ),
.O5(CLBLM_R_X63Y106_SLICE_X95Y106_DO5),
.O6(CLBLM_R_X63Y106_SLICE_X95Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X63Y106_SLICE_X95Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X64Y106_SLICE_X96Y106_BQ),
.O5(CLBLM_R_X63Y106_SLICE_X95Y106_CO5),
.O6(CLBLM_R_X63Y106_SLICE_X95Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X63Y106_SLICE_X95Y106_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X64Y106_SLICE_X96Y106_AQ),
.O5(CLBLM_R_X63Y106_SLICE_X95Y106_BO5),
.O6(CLBLM_R_X63Y106_SLICE_X95Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X63Y106_SLICE_X95Y106_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X62Y105_SLICE_X93Y105_BQ),
.O5(CLBLM_R_X63Y106_SLICE_X95Y106_AO5),
.O6(CLBLM_R_X63Y106_SLICE_X95Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X63Y107_SLICE_X94Y107_CARRY4 (
.CI(CLBLM_R_X63Y106_SLICE_X94Y106_COUT),
.CO({CLBLM_R_X63Y107_SLICE_X94Y107_D_CY, CLBLM_R_X63Y107_SLICE_X94Y107_C_CY, CLBLM_R_X63Y107_SLICE_X94Y107_B_CY, CLBLM_R_X63Y107_SLICE_X94Y107_A_CY}),
.CYINIT(1'b0),
.DI({CLBLM_L_X64Y107_SLICE_X97Y107_AQ, CLBLM_L_X64Y107_SLICE_X96Y107_BQ, CLBLM_L_X64Y107_SLICE_X96Y107_AQ, CLBLM_L_X64Y107_SLICE_X97Y107_BQ}),
.O({CLBLM_R_X63Y107_SLICE_X94Y107_D_XOR, CLBLM_R_X63Y107_SLICE_X94Y107_C_XOR, CLBLM_R_X63Y107_SLICE_X94Y107_B_XOR, CLBLM_R_X63Y107_SLICE_X94Y107_A_XOR}),
.S({CLBLM_R_X63Y107_SLICE_X94Y107_DO6, CLBLM_R_X63Y107_SLICE_X94Y107_CO6, CLBLM_R_X63Y107_SLICE_X94Y107_BO6, CLBLM_R_X63Y107_SLICE_X94Y107_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333333333333)
  ) CLBLM_R_X63Y107_SLICE_X94Y107_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X64Y107_SLICE_X97Y107_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y107_SLICE_X94Y107_DO5),
.O6(CLBLM_R_X63Y107_SLICE_X94Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00ff00ff)
  ) CLBLM_R_X63Y107_SLICE_X94Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X64Y107_SLICE_X96Y107_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y107_SLICE_X94Y107_CO5),
.O6(CLBLM_R_X63Y107_SLICE_X94Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555555)
  ) CLBLM_R_X63Y107_SLICE_X94Y107_BLUT (
.I0(CLBLM_L_X64Y107_SLICE_X96Y107_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y107_SLICE_X94Y107_BO5),
.O6(CLBLM_R_X63Y107_SLICE_X94Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0f0f0f)
  ) CLBLM_R_X63Y107_SLICE_X94Y107_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X64Y107_SLICE_X97Y107_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y107_SLICE_X94Y107_AO5),
.O6(CLBLM_R_X63Y107_SLICE_X94Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X63Y107_SLICE_X95Y107_CARRY4 (
.CI(CLBLM_R_X63Y106_SLICE_X95Y106_COUT),
.CO({CLBLM_R_X63Y107_SLICE_X95Y107_D_CY, CLBLM_R_X63Y107_SLICE_X95Y107_C_CY, CLBLM_R_X63Y107_SLICE_X95Y107_B_CY, CLBLM_R_X63Y107_SLICE_X95Y107_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X63Y107_SLICE_X95Y107_D_XOR, CLBLM_R_X63Y107_SLICE_X95Y107_C_XOR, CLBLM_R_X63Y107_SLICE_X95Y107_B_XOR, CLBLM_R_X63Y107_SLICE_X95Y107_A_XOR}),
.S({CLBLM_R_X63Y107_SLICE_X95Y107_DO6, CLBLM_R_X63Y107_SLICE_X95Y107_CO6, CLBLM_R_X63Y107_SLICE_X95Y107_BO6, CLBLM_R_X63Y107_SLICE_X95Y107_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X63Y107_SLICE_X95Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X64Y108_SLICE_X96Y108_AQ),
.O5(CLBLM_R_X63Y107_SLICE_X95Y107_DO5),
.O6(CLBLM_R_X63Y107_SLICE_X95Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X63Y107_SLICE_X95Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X64Y107_SLICE_X97Y107_AQ),
.O5(CLBLM_R_X63Y107_SLICE_X95Y107_CO5),
.O6(CLBLM_R_X63Y107_SLICE_X95Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X63Y107_SLICE_X95Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X64Y107_SLICE_X96Y107_BQ),
.O5(CLBLM_R_X63Y107_SLICE_X95Y107_BO5),
.O6(CLBLM_R_X63Y107_SLICE_X95Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X63Y107_SLICE_X95Y107_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X64Y107_SLICE_X96Y107_AQ),
.O5(CLBLM_R_X63Y107_SLICE_X95Y107_AO5),
.O6(CLBLM_R_X63Y107_SLICE_X95Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X63Y108_SLICE_X94Y108_CARRY4 (
.CI(CLBLM_R_X63Y107_SLICE_X94Y107_COUT),
.CO({CLBLM_R_X63Y108_SLICE_X94Y108_D_CY, CLBLM_R_X63Y108_SLICE_X94Y108_C_CY, CLBLM_R_X63Y108_SLICE_X94Y108_B_CY, CLBLM_R_X63Y108_SLICE_X94Y108_A_CY}),
.CYINIT(1'b0),
.DI({CLBLM_L_X64Y108_SLICE_X96Y108_BQ, CLBLM_R_X63Y110_SLICE_X94Y110_AQ, CLBLM_L_X64Y108_SLICE_X97Y108_AQ, CLBLM_L_X64Y108_SLICE_X96Y108_AQ}),
.O({CLBLM_R_X63Y108_SLICE_X94Y108_D_XOR, CLBLM_R_X63Y108_SLICE_X94Y108_C_XOR, CLBLM_R_X63Y108_SLICE_X94Y108_B_XOR, CLBLM_R_X63Y108_SLICE_X94Y108_A_XOR}),
.S({CLBLM_R_X63Y108_SLICE_X94Y108_DO6, CLBLM_R_X63Y108_SLICE_X94Y108_CO6, CLBLM_R_X63Y108_SLICE_X94Y108_BO6, CLBLM_R_X63Y108_SLICE_X94Y108_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555555)
  ) CLBLM_R_X63Y108_SLICE_X94Y108_DLUT (
.I0(CLBLM_L_X64Y108_SLICE_X96Y108_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y108_SLICE_X94Y108_DO5),
.O6(CLBLM_R_X63Y108_SLICE_X94Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555555)
  ) CLBLM_R_X63Y108_SLICE_X94Y108_CLUT (
.I0(CLBLM_R_X63Y110_SLICE_X94Y110_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y108_SLICE_X94Y108_CO5),
.O6(CLBLM_R_X63Y108_SLICE_X94Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffffffff)
  ) CLBLM_R_X63Y108_SLICE_X94Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X64Y108_SLICE_X97Y108_AQ),
.O5(CLBLM_R_X63Y108_SLICE_X94Y108_BO5),
.O6(CLBLM_R_X63Y108_SLICE_X94Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00ff00ff)
  ) CLBLM_R_X63Y108_SLICE_X94Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X64Y108_SLICE_X96Y108_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y108_SLICE_X94Y108_AO5),
.O6(CLBLM_R_X63Y108_SLICE_X94Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X63Y108_SLICE_X95Y108_CARRY4 (
.CI(CLBLM_R_X63Y107_SLICE_X95Y107_COUT),
.CO({CLBLM_R_X63Y108_SLICE_X95Y108_D_CY, CLBLM_R_X63Y108_SLICE_X95Y108_C_CY, CLBLM_R_X63Y108_SLICE_X95Y108_B_CY, CLBLM_R_X63Y108_SLICE_X95Y108_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X63Y108_SLICE_X95Y108_D_XOR, CLBLM_R_X63Y108_SLICE_X95Y108_C_XOR, CLBLM_R_X63Y108_SLICE_X95Y108_B_XOR, CLBLM_R_X63Y108_SLICE_X95Y108_A_XOR}),
.S({CLBLM_R_X63Y108_SLICE_X95Y108_DO6, CLBLM_R_X63Y108_SLICE_X95Y108_CO6, CLBLM_R_X63Y108_SLICE_X95Y108_BO6, CLBLM_R_X63Y108_SLICE_X95Y108_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X63Y108_SLICE_X95Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X64Y109_SLICE_X96Y109_AQ),
.O5(CLBLM_R_X63Y108_SLICE_X95Y108_DO5),
.O6(CLBLM_R_X63Y108_SLICE_X95Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X63Y108_SLICE_X95Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X64Y108_SLICE_X96Y108_BQ),
.O5(CLBLM_R_X63Y108_SLICE_X95Y108_CO5),
.O6(CLBLM_R_X63Y108_SLICE_X95Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X63Y108_SLICE_X95Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X63Y110_SLICE_X94Y110_AQ),
.O5(CLBLM_R_X63Y108_SLICE_X95Y108_BO5),
.O6(CLBLM_R_X63Y108_SLICE_X95Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X63Y108_SLICE_X95Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X64Y108_SLICE_X97Y108_AQ),
.O5(CLBLM_R_X63Y108_SLICE_X95Y108_AO5),
.O6(CLBLM_R_X63Y108_SLICE_X95Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X63Y109_SLICE_X94Y109_CARRY4 (
.CI(CLBLM_R_X63Y108_SLICE_X94Y108_COUT),
.CO({CLBLM_R_X63Y109_SLICE_X94Y109_D_CY, CLBLM_R_X63Y109_SLICE_X94Y109_C_CY, CLBLM_R_X63Y109_SLICE_X94Y109_B_CY, CLBLM_R_X63Y109_SLICE_X94Y109_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, CLBLM_R_X63Y105_SLICE_X94Y105_AQ, CLBLM_L_X62Y103_SLICE_X93Y103_AQ, CLBLM_L_X64Y109_SLICE_X96Y109_AQ}),
.O({CLBLM_R_X63Y109_SLICE_X94Y109_D_XOR, CLBLM_R_X63Y109_SLICE_X94Y109_C_XOR, CLBLM_R_X63Y109_SLICE_X94Y109_B_XOR, CLBLM_R_X63Y109_SLICE_X94Y109_A_XOR}),
.S({CLBLM_R_X63Y109_SLICE_X94Y109_DO6, CLBLM_R_X63Y109_SLICE_X94Y109_CO6, CLBLM_R_X63Y109_SLICE_X94Y109_BO6, CLBLM_R_X63Y109_SLICE_X94Y109_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffffffff)
  ) CLBLM_R_X63Y109_SLICE_X94Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X64Y109_SLICE_X96Y109_A5Q),
.O5(CLBLM_R_X63Y109_SLICE_X94Y109_DO5),
.O6(CLBLM_R_X63Y109_SLICE_X94Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555555)
  ) CLBLM_R_X63Y109_SLICE_X94Y109_CLUT (
.I0(CLBLM_R_X63Y105_SLICE_X94Y105_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y109_SLICE_X94Y109_CO5),
.O6(CLBLM_R_X63Y109_SLICE_X94Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333333333333)
  ) CLBLM_R_X63Y109_SLICE_X94Y109_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X62Y103_SLICE_X93Y103_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y109_SLICE_X94Y109_BO5),
.O6(CLBLM_R_X63Y109_SLICE_X94Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffff0000ffff)
  ) CLBLM_R_X63Y109_SLICE_X94Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X64Y109_SLICE_X96Y109_AQ),
.I5(1'b1),
.O5(CLBLM_R_X63Y109_SLICE_X94Y109_AO5),
.O6(CLBLM_R_X63Y109_SLICE_X94Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X63Y109_SLICE_X95Y109_CARRY4 (
.CI(CLBLM_R_X63Y108_SLICE_X95Y108_COUT),
.CO({CLBLM_R_X63Y109_SLICE_X95Y109_D_CY, CLBLM_R_X63Y109_SLICE_X95Y109_C_CY, CLBLM_R_X63Y109_SLICE_X95Y109_B_CY, CLBLM_R_X63Y109_SLICE_X95Y109_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X63Y109_SLICE_X95Y109_D_XOR, CLBLM_R_X63Y109_SLICE_X95Y109_C_XOR, CLBLM_R_X63Y109_SLICE_X95Y109_B_XOR, CLBLM_R_X63Y109_SLICE_X95Y109_A_XOR}),
.S({CLBLM_R_X63Y109_SLICE_X95Y109_DO6, CLBLM_R_X63Y109_SLICE_X95Y109_CO6, CLBLM_R_X63Y109_SLICE_X95Y109_BO6, CLBLM_R_X63Y109_SLICE_X95Y109_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y109_SLICE_X95Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y109_SLICE_X95Y109_DO5),
.O6(CLBLM_R_X63Y109_SLICE_X95Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X63Y109_SLICE_X95Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X64Y109_SLICE_X96Y109_A5Q),
.O5(CLBLM_R_X63Y109_SLICE_X95Y109_CO5),
.O6(CLBLM_R_X63Y109_SLICE_X95Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X63Y109_SLICE_X95Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X63Y105_SLICE_X94Y105_AQ),
.O5(CLBLM_R_X63Y109_SLICE_X95Y109_BO5),
.O6(CLBLM_R_X63Y109_SLICE_X95Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X63Y109_SLICE_X95Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X62Y103_SLICE_X93Y103_AQ),
.O5(CLBLM_R_X63Y109_SLICE_X95Y109_AO5),
.O6(CLBLM_R_X63Y109_SLICE_X95Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X63Y110_SLICE_X94Y110_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_R_X63Y100_SLICE_X94Y100_CO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X63Y110_SLICE_X94Y110_AO6),
.Q(CLBLM_R_X63Y110_SLICE_X94Y110_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y110_SLICE_X94Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y110_SLICE_X94Y110_DO5),
.O6(CLBLM_R_X63Y110_SLICE_X94Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff35cf05fa30ca00)
  ) CLBLM_R_X63Y110_SLICE_X94Y110_CLUT (
.I0(CLBLM_L_X62Y105_SLICE_X92Y105_BO5),
.I1(CLBLM_L_X62Y105_SLICE_X93Y105_AO6),
.I2(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I3(CLBLM_R_X63Y109_SLICE_X95Y109_A_XOR),
.I4(CLBLM_R_X63Y109_SLICE_X94Y109_B_XOR),
.I5(CLBLM_L_X62Y103_SLICE_X93Y103_AQ),
.O5(CLBLM_R_X63Y110_SLICE_X94Y110_CO5),
.O6(CLBLM_R_X63Y110_SLICE_X94Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0cacacfc0)
  ) CLBLM_R_X63Y110_SLICE_X94Y110_BLUT (
.I0(CLBLM_R_X63Y108_SLICE_X95Y108_B_XOR),
.I1(CLBLM_L_X50Y107_SLICE_X76Y107_BQ),
.I2(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I3(CLBLM_R_X63Y110_SLICE_X94Y110_AQ),
.I4(CLBLM_L_X62Y105_SLICE_X92Y105_BO5),
.I5(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.O5(CLBLM_R_X63Y110_SLICE_X94Y110_BO5),
.O6(CLBLM_R_X63Y110_SLICE_X94Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0bff08ff00ff00)
  ) CLBLM_R_X63Y110_SLICE_X94Y110_ALUT (
.I0(CLBLM_R_X63Y108_SLICE_X95Y108_B_XOR),
.I1(CLBLM_L_X62Y105_SLICE_X93Y105_AO6),
.I2(CLBLM_L_X62Y112_SLICE_X92Y112_AQ),
.I3(CLBLM_R_X63Y110_SLICE_X94Y110_BO6),
.I4(CLBLM_R_X63Y108_SLICE_X94Y108_C_XOR),
.I5(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.O5(CLBLM_R_X63Y110_SLICE_X94Y110_AO5),
.O6(CLBLM_R_X63Y110_SLICE_X94Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y110_SLICE_X95Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y110_SLICE_X95Y110_DO5),
.O6(CLBLM_R_X63Y110_SLICE_X95Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y110_SLICE_X95Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y110_SLICE_X95Y110_CO5),
.O6(CLBLM_R_X63Y110_SLICE_X95Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y110_SLICE_X95Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y110_SLICE_X95Y110_BO5),
.O6(CLBLM_R_X63Y110_SLICE_X95Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X63Y110_SLICE_X95Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X63Y110_SLICE_X95Y110_AO5),
.O6(CLBLM_R_X63Y110_SLICE_X95Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y96_SLICE_X98Y96_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y96_SLICE_X98Y96_DO5),
.O6(CLBLM_R_X65Y96_SLICE_X98Y96_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y96_SLICE_X98Y96_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y96_SLICE_X98Y96_CO5),
.O6(CLBLM_R_X65Y96_SLICE_X98Y96_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0c0c0c00000808)
  ) CLBLM_R_X65Y96_SLICE_X98Y96_BLUT (
.I0(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I1(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I2(CLBLM_L_X56Y97_SLICE_X85Y97_AQ),
.I3(1'b1),
.I4(CLBLM_R_X63Y95_SLICE_X95Y95_D5Q),
.I5(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.O5(CLBLM_R_X65Y96_SLICE_X98Y96_BO5),
.O6(CLBLM_R_X65Y96_SLICE_X98Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0c0c0c00080008)
  ) CLBLM_R_X65Y96_SLICE_X98Y96_ALUT (
.I0(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I1(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I2(CLBLM_L_X56Y97_SLICE_X85Y97_AQ),
.I3(CLBLM_R_X63Y95_SLICE_X95Y95_CQ),
.I4(1'b1),
.I5(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.O5(CLBLM_R_X65Y96_SLICE_X98Y96_AO5),
.O6(CLBLM_R_X65Y96_SLICE_X98Y96_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y96_SLICE_X99Y96_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y96_SLICE_X99Y96_DO5),
.O6(CLBLM_R_X65Y96_SLICE_X99Y96_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y96_SLICE_X99Y96_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y96_SLICE_X99Y96_CO5),
.O6(CLBLM_R_X65Y96_SLICE_X99Y96_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y96_SLICE_X99Y96_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y96_SLICE_X99Y96_BO5),
.O6(CLBLM_R_X65Y96_SLICE_X99Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y96_SLICE_X99Y96_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y96_SLICE_X99Y96_AO5),
.O6(CLBLM_R_X65Y96_SLICE_X99Y96_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5000500055005000)
  ) CLBLM_R_X65Y97_SLICE_X98Y97_DLUT (
.I0(CLBLM_L_X56Y97_SLICE_X85Y97_AQ),
.I1(1'b1),
.I2(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I3(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I4(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I5(CLBLM_R_X63Y96_SLICE_X95Y96_BQ),
.O5(CLBLM_R_X65Y97_SLICE_X98Y97_DO5),
.O6(CLBLM_R_X65Y97_SLICE_X98Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5500100055001000)
  ) CLBLM_R_X65Y97_SLICE_X98Y97_CLUT (
.I0(CLBLM_L_X56Y97_SLICE_X85Y97_AQ),
.I1(CLBLM_L_X64Y97_SLICE_X97Y97_BQ),
.I2(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I3(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I4(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I5(1'b1),
.O5(CLBLM_R_X65Y97_SLICE_X98Y97_CO5),
.O6(CLBLM_R_X65Y97_SLICE_X98Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0e0c0e00000000)
  ) CLBLM_R_X65Y97_SLICE_X98Y97_BLUT (
.I0(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I1(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I2(CLBLM_L_X56Y97_SLICE_X85Y97_AQ),
.I3(CLBLM_L_X64Y97_SLICE_X97Y97_AQ),
.I4(1'b1),
.I5(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.O5(CLBLM_R_X65Y97_SLICE_X98Y97_BO5),
.O6(CLBLM_R_X65Y97_SLICE_X98Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000033ffa0aa8888)
  ) CLBLM_R_X65Y97_SLICE_X98Y97_ALUT (
.I0(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I1(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I2(CLBLM_L_X60Y98_SLICE_X90Y98_AQ),
.I3(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I4(CLBLM_L_X56Y97_SLICE_X85Y97_AQ),
.I5(1'b1),
.O5(CLBLM_R_X65Y97_SLICE_X98Y97_AO5),
.O6(CLBLM_R_X65Y97_SLICE_X98Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y97_SLICE_X99Y97_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y97_SLICE_X99Y97_DO5),
.O6(CLBLM_R_X65Y97_SLICE_X99Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5500550000005000)
  ) CLBLM_R_X65Y97_SLICE_X99Y97_CLUT (
.I0(CLBLM_L_X56Y97_SLICE_X85Y97_AQ),
.I1(1'b1),
.I2(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I3(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I4(CLBLM_R_X63Y95_SLICE_X95Y95_C5Q),
.I5(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.O5(CLBLM_R_X65Y97_SLICE_X99Y97_CO5),
.O6(CLBLM_R_X65Y97_SLICE_X99Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f050000000000)
  ) CLBLM_R_X65Y97_SLICE_X99Y97_BLUT (
.I0(CLBLM_L_X62Y96_SLICE_X93Y96_CQ),
.I1(1'b1),
.I2(CLBLM_L_X56Y97_SLICE_X85Y97_AQ),
.I3(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I4(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I5(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.O5(CLBLM_R_X65Y97_SLICE_X99Y97_BO5),
.O6(CLBLM_R_X65Y97_SLICE_X99Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f000f0a00000000)
  ) CLBLM_R_X65Y97_SLICE_X99Y97_ALUT (
.I0(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I1(1'b1),
.I2(CLBLM_L_X56Y97_SLICE_X85Y97_AQ),
.I3(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I4(CLBLM_L_X62Y96_SLICE_X93Y96_DQ),
.I5(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.O5(CLBLM_R_X65Y97_SLICE_X99Y97_AO5),
.O6(CLBLM_R_X65Y97_SLICE_X99Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X65Y98_SLICE_X98Y98_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_BQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X65Y98_SLICE_X98Y98_AO6),
.Q(CLBLM_R_X65Y98_SLICE_X98Y98_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X65Y98_SLICE_X98Y98_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_BQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X65Y98_SLICE_X98Y98_BO6),
.Q(CLBLM_R_X65Y98_SLICE_X98Y98_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h50f0505050505050)
  ) CLBLM_R_X65Y98_SLICE_X98Y98_DLUT (
.I0(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I1(1'b1),
.I2(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I3(CLBLM_R_X65Y102_SLICE_X98Y102_A_XOR),
.I4(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I5(CLBLM_L_X60Y98_SLICE_X90Y98_AQ),
.O5(CLBLM_R_X65Y98_SLICE_X98Y98_DO5),
.O6(CLBLM_R_X65Y98_SLICE_X98Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3310333033133333)
  ) CLBLM_R_X65Y98_SLICE_X98Y98_CLUT (
.I0(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I1(CLBLM_R_X65Y101_SLICE_X99Y101_BO6),
.I2(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I3(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I4(CLBLM_L_X64Y100_SLICE_X97Y100_AQ),
.I5(CLBLM_L_X64Y100_SLICE_X96Y100_D_XOR),
.O5(CLBLM_R_X65Y98_SLICE_X98Y98_CO5),
.O6(CLBLM_R_X65Y98_SLICE_X98Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000cccc0000ffff)
  ) CLBLM_R_X65Y98_SLICE_X98Y98_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X65Y97_SLICE_X98Y97_AO5),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X64Y98_SLICE_X96Y98_BO6),
.I5(CLBLM_R_X65Y100_SLICE_X99Y100_CQ),
.O5(CLBLM_R_X65Y98_SLICE_X98Y98_BO5),
.O6(CLBLM_R_X65Y98_SLICE_X98Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3030300032323200)
  ) CLBLM_R_X65Y98_SLICE_X98Y98_ALUT (
.I0(CLBLM_R_X65Y98_SLICE_X99Y98_CO6),
.I1(CLBLM_R_X65Y97_SLICE_X98Y97_BO6),
.I2(CLBLM_R_X65Y97_SLICE_X98Y97_AO6),
.I3(CLBLM_R_X65Y97_SLICE_X98Y97_AO5),
.I4(CLBLM_L_X64Y102_SLICE_X96Y102_C_XOR),
.I5(CLBLM_R_X65Y102_SLICE_X99Y102_BO6),
.O5(CLBLM_R_X65Y98_SLICE_X98Y98_AO5),
.O6(CLBLM_R_X65Y98_SLICE_X98Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X65Y98_SLICE_X99Y98_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_BQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X65Y98_SLICE_X99Y98_AO6),
.Q(CLBLM_R_X65Y98_SLICE_X99Y98_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0c0f0f0c0c0000)
  ) CLBLM_R_X65Y98_SLICE_X99Y98_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X63Y95_SLICE_X95Y95_B5Q),
.I2(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I3(1'b1),
.I4(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I5(CLBLM_L_X64Y100_SLICE_X96Y100_D_XOR),
.O5(CLBLM_R_X65Y98_SLICE_X99Y98_DO5),
.O6(CLBLM_R_X65Y98_SLICE_X99Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcffffaaaaffff)
  ) CLBLM_R_X65Y98_SLICE_X99Y98_CLUT (
.I0(CLBLM_L_X64Y102_SLICE_X97Y102_D_XOR),
.I1(CLBLM_R_X49Y104_SLICE_X75Y104_CQ),
.I2(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I3(1'b1),
.I4(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I5(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.O5(CLBLM_R_X65Y98_SLICE_X99Y98_CO5),
.O6(CLBLM_R_X65Y98_SLICE_X99Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h77007f000000ff00)
  ) CLBLM_R_X65Y98_SLICE_X99Y98_BLUT (
.I0(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I1(CLBLM_L_X60Y98_SLICE_X90Y98_AQ),
.I2(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I3(CLBLM_L_X64Y100_SLICE_X96Y100_D_XOR),
.I4(CLBLM_L_X56Y97_SLICE_X85Y97_AQ),
.I5(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.O5(CLBLM_R_X65Y98_SLICE_X99Y98_BO5),
.O6(CLBLM_R_X65Y98_SLICE_X99Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fff0faaaaff00)
  ) CLBLM_R_X65Y98_SLICE_X99Y98_ALUT (
.I0(CLBLM_R_X65Y98_SLICE_X99Y98_DO6),
.I1(1'b1),
.I2(CLBLM_R_X65Y98_SLICE_X98Y98_CO6),
.I3(CLBLM_R_X65Y98_SLICE_X99Y98_BO6),
.I4(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I5(CLBLM_L_X56Y97_SLICE_X85Y97_AQ),
.O5(CLBLM_R_X65Y98_SLICE_X99Y98_AO5),
.O6(CLBLM_R_X65Y98_SLICE_X99Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X65Y99_SLICE_X98Y99_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_BQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X65Y99_SLICE_X98Y99_AO6),
.Q(CLBLM_R_X65Y99_SLICE_X98Y99_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeeffffe2e2ffff)
  ) CLBLM_R_X65Y99_SLICE_X98Y99_DLUT (
.I0(CLBLM_L_X64Y100_SLICE_X97Y100_C_XOR),
.I1(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I2(CLBLM_L_X62Y101_SLICE_X93Y101_AQ),
.I3(1'b1),
.I4(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I5(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.O5(CLBLM_R_X65Y99_SLICE_X98Y99_DO5),
.O6(CLBLM_R_X65Y99_SLICE_X98Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55dd555500000000)
  ) CLBLM_R_X65Y99_SLICE_X98Y99_CLUT (
.I0(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I1(CLBLM_L_X60Y98_SLICE_X90Y98_AQ),
.I2(1'b1),
.I3(CLBLM_R_X65Y100_SLICE_X98Y100_C_XOR),
.I4(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I5(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.O5(CLBLM_R_X65Y99_SLICE_X98Y99_CO5),
.O6(CLBLM_R_X65Y99_SLICE_X98Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00c000c000e000e0)
  ) CLBLM_R_X65Y99_SLICE_X98Y99_BLUT (
.I0(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I1(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I2(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I3(CLBLM_L_X56Y97_SLICE_X85Y97_AQ),
.I4(1'b1),
.I5(CLBLM_R_X63Y97_SLICE_X94Y97_DQ),
.O5(CLBLM_R_X65Y99_SLICE_X98Y99_BO5),
.O6(CLBLM_R_X65Y99_SLICE_X98Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0c00000f0c0a08)
  ) CLBLM_R_X65Y99_SLICE_X98Y99_ALUT (
.I0(CLBLM_R_X65Y99_SLICE_X98Y99_DO6),
.I1(CLBLM_R_X65Y97_SLICE_X98Y97_AO5),
.I2(CLBLM_R_X65Y96_SLICE_X98Y96_AO6),
.I3(CLBLM_L_X64Y100_SLICE_X96Y100_B_XOR),
.I4(CLBLM_R_X65Y97_SLICE_X98Y97_AO6),
.I5(CLBLM_R_X65Y99_SLICE_X98Y99_CO6),
.O5(CLBLM_R_X65Y99_SLICE_X98Y99_AO5),
.O6(CLBLM_R_X65Y99_SLICE_X98Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X65Y99_SLICE_X99Y99_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_BQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X65Y99_SLICE_X99Y99_AO6),
.Q(CLBLM_R_X65Y99_SLICE_X99Y99_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0ff00ff00000000)
  ) CLBLM_R_X65Y99_SLICE_X99Y99_DLUT (
.I0(CLBLM_R_X65Y100_SLICE_X98Y100_D_XOR),
.I1(1'b1),
.I2(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I3(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I4(CLBLM_L_X60Y98_SLICE_X90Y98_AQ),
.I5(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.O5(CLBLM_R_X65Y99_SLICE_X99Y99_DO5),
.O6(CLBLM_R_X65Y99_SLICE_X99Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55f5555500000000)
  ) CLBLM_R_X65Y99_SLICE_X99Y99_CLUT (
.I0(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I1(1'b1),
.I2(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I3(CLBLM_R_X65Y100_SLICE_X98Y100_B_XOR),
.I4(CLBLM_L_X60Y98_SLICE_X90Y98_AQ),
.I5(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.O5(CLBLM_R_X65Y99_SLICE_X99Y99_CO5),
.O6(CLBLM_R_X65Y99_SLICE_X99Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ff220000)
  ) CLBLM_R_X65Y99_SLICE_X99Y99_BLUT (
.I0(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I1(CLBLM_R_X63Y95_SLICE_X95Y95_BQ),
.I2(1'b1),
.I3(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I4(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I5(CLBLM_L_X56Y97_SLICE_X85Y97_AQ),
.O5(CLBLM_R_X65Y99_SLICE_X99Y99_BO5),
.O6(CLBLM_R_X65Y99_SLICE_X99Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff003000aa0020)
  ) CLBLM_R_X65Y99_SLICE_X99Y99_ALUT (
.I0(CLBLM_L_X64Y100_SLICE_X96Y100_A_XOR),
.I1(CLBLM_R_X65Y99_SLICE_X99Y99_CO6),
.I2(CLBLM_R_X65Y100_SLICE_X99Y100_DO6),
.I3(CLBLM_R_X65Y99_SLICE_X99Y99_BO6),
.I4(CLBLM_R_X65Y97_SLICE_X98Y97_AO6),
.I5(CLBLM_R_X65Y97_SLICE_X98Y97_AO5),
.O5(CLBLM_R_X65Y99_SLICE_X99Y99_AO5),
.O6(CLBLM_R_X65Y99_SLICE_X99Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X65Y100_SLICE_X98Y100_CARRY4 (
.CI(1'b0),
.CO({CLBLM_R_X65Y100_SLICE_X98Y100_D_CY, CLBLM_R_X65Y100_SLICE_X98Y100_C_CY, CLBLM_R_X65Y100_SLICE_X98Y100_B_CY, CLBLM_R_X65Y100_SLICE_X98Y100_A_CY}),
.CYINIT(1'b0),
.DI({CLBLM_L_X64Y106_SLICE_X97Y106_DQ, CLBLM_R_X65Y106_SLICE_X98Y106_CQ, CLBLM_R_X65Y100_SLICE_X99Y100_AQ, CLBLM_R_X65Y100_SLICE_X99Y100_CQ}),
.O({CLBLM_R_X65Y100_SLICE_X98Y100_D_XOR, CLBLM_R_X65Y100_SLICE_X98Y100_C_XOR, CLBLM_R_X65Y100_SLICE_X98Y100_B_XOR, CLBLM_R_X65Y100_SLICE_X98Y100_A_XOR}),
.S({CLBLM_R_X65Y100_SLICE_X98Y100_DO6, CLBLM_R_X65Y100_SLICE_X98Y100_CO6, CLBLM_R_X65Y100_SLICE_X98Y100_BO6, CLBLM_R_X65Y100_SLICE_X98Y100_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0ff0f0f0f0)
  ) CLBLM_R_X65Y100_SLICE_X98Y100_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X64Y106_SLICE_X97Y106_DQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X62Y100_SLICE_X92Y100_CQ),
.O5(CLBLM_R_X65Y100_SLICE_X98Y100_DO5),
.O6(CLBLM_R_X65Y100_SLICE_X98Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3c3c3c3c3c)
  ) CLBLM_R_X65Y100_SLICE_X98Y100_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X62Y101_SLICE_X93Y101_AQ),
.I2(CLBLM_R_X65Y106_SLICE_X98Y106_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y100_SLICE_X98Y100_CO5),
.O6(CLBLM_R_X65Y100_SLICE_X98Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0ff0f00f0ff0f0)
  ) CLBLM_R_X65Y100_SLICE_X98Y100_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X62Y100_SLICE_X92Y100_BQ),
.I3(1'b1),
.I4(CLBLM_R_X65Y100_SLICE_X99Y100_AQ),
.I5(1'b1),
.O5(CLBLM_R_X65Y100_SLICE_X98Y100_BO5),
.O6(CLBLM_R_X65Y100_SLICE_X98Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ffff00ff00)
  ) CLBLM_R_X65Y100_SLICE_X98Y100_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X62Y100_SLICE_X92Y100_AQ),
.I4(1'b1),
.I5(CLBLM_R_X65Y100_SLICE_X99Y100_CQ),
.O5(CLBLM_R_X65Y100_SLICE_X98Y100_AO5),
.O6(CLBLM_R_X65Y100_SLICE_X98Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X65Y100_SLICE_X99Y100_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y105_SLICE_X93Y105_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X65Y100_SLICE_X99Y100_AO6),
.Q(CLBLM_R_X65Y100_SLICE_X99Y100_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X65Y100_SLICE_X99Y100_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y105_SLICE_X93Y105_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X65Y100_SLICE_X99Y100_BO6),
.Q(CLBLM_R_X65Y100_SLICE_X99Y100_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X65Y100_SLICE_X99Y100_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y105_SLICE_X93Y105_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X65Y100_SLICE_X99Y100_CO6),
.Q(CLBLM_R_X65Y100_SLICE_X99Y100_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfdfd5dfdfdfd5d)
  ) CLBLM_R_X65Y100_SLICE_X99Y100_DLUT (
.I0(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I1(CLBLM_L_X64Y100_SLICE_X97Y100_B_XOR),
.I2(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I3(CLBLM_L_X62Y100_SLICE_X92Y100_BQ),
.I4(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I5(1'b1),
.O5(CLBLM_R_X65Y100_SLICE_X99Y100_DO5),
.O6(CLBLM_R_X65Y100_SLICE_X99Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9999f0f00000f0f0)
  ) CLBLM_R_X65Y100_SLICE_X99Y100_CLUT (
.I0(CLBLL_R_X57Y103_SLICE_X86Y103_AQ),
.I1(CLBLL_R_X57Y103_SLICE_X86Y103_A5Q),
.I2(CLBLM_R_X63Y104_SLICE_X94Y104_AQ),
.I3(1'b1),
.I4(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I5(CLBLM_R_X65Y98_SLICE_X98Y98_BQ),
.O5(CLBLM_R_X65Y100_SLICE_X99Y100_CO5),
.O6(CLBLM_R_X65Y100_SLICE_X99Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a055005500f5a0)
  ) CLBLM_R_X65Y100_SLICE_X99Y100_BLUT (
.I0(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I1(1'b1),
.I2(CLBLM_R_X65Y98_SLICE_X99Y98_AQ),
.I3(CLBLM_L_X62Y105_SLICE_X93Y105_BQ),
.I4(CLBLL_R_X57Y103_SLICE_X86Y103_AQ),
.I5(CLBLL_R_X57Y103_SLICE_X86Y103_A5Q),
.O5(CLBLM_R_X65Y100_SLICE_X99Y100_BO5),
.O6(CLBLM_R_X65Y100_SLICE_X99Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd8855005500dd88)
  ) CLBLM_R_X65Y100_SLICE_X99Y100_ALUT (
.I0(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I1(CLBLM_R_X65Y99_SLICE_X99Y99_AQ),
.I2(1'b1),
.I3(CLBLM_L_X64Y105_SLICE_X96Y105_AQ),
.I4(CLBLL_R_X57Y103_SLICE_X86Y103_AQ),
.I5(CLBLL_R_X57Y103_SLICE_X86Y103_A5Q),
.O5(CLBLM_R_X65Y100_SLICE_X99Y100_AO5),
.O6(CLBLM_R_X65Y100_SLICE_X99Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X65Y101_SLICE_X98Y101_CARRY4 (
.CI(CLBLM_R_X65Y100_SLICE_X98Y100_COUT),
.CO({CLBLM_R_X65Y101_SLICE_X98Y101_D_CY, CLBLM_R_X65Y101_SLICE_X98Y101_C_CY, CLBLM_R_X65Y101_SLICE_X98Y101_B_CY, CLBLM_R_X65Y101_SLICE_X98Y101_A_CY}),
.CYINIT(1'b0),
.DI({CLBLM_L_X62Y101_SLICE_X93Y101_CQ, CLBLM_R_X63Y103_SLICE_X95Y103_BQ, CLBLM_R_X65Y106_SLICE_X98Y106_DQ, CLBLM_R_X65Y100_SLICE_X99Y100_BQ}),
.O({CLBLM_R_X65Y101_SLICE_X98Y101_D_XOR, CLBLM_R_X65Y101_SLICE_X98Y101_C_XOR, CLBLM_R_X65Y101_SLICE_X98Y101_B_XOR, CLBLM_R_X65Y101_SLICE_X98Y101_A_XOR}),
.S({CLBLM_R_X65Y101_SLICE_X98Y101_DO6, CLBLM_R_X65Y101_SLICE_X98Y101_CO6, CLBLM_R_X65Y101_SLICE_X98Y101_BO6, CLBLM_R_X65Y101_SLICE_X98Y101_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5a5a5a5a5a)
  ) CLBLM_R_X65Y101_SLICE_X98Y101_DLUT (
.I0(CLBLM_R_X63Y101_SLICE_X95Y101_AQ),
.I1(1'b1),
.I2(CLBLM_L_X62Y101_SLICE_X93Y101_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y101_SLICE_X98Y101_DO5),
.O6(CLBLM_R_X65Y101_SLICE_X98Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0ff0f0f0f0)
  ) CLBLM_R_X65Y101_SLICE_X98Y101_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X62Y101_SLICE_X93Y101_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X63Y103_SLICE_X95Y103_BQ),
.O5(CLBLM_R_X65Y101_SLICE_X98Y101_CO5),
.O6(CLBLM_R_X65Y101_SLICE_X98Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6666666666666666)
  ) CLBLM_R_X65Y101_SLICE_X98Y101_BLUT (
.I0(CLBLM_R_X65Y106_SLICE_X98Y106_DQ),
.I1(CLBLM_L_X64Y100_SLICE_X97Y100_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y101_SLICE_X98Y101_BO5),
.O6(CLBLM_R_X65Y101_SLICE_X98Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0ff0f00f0ff0f0)
  ) CLBLM_R_X65Y101_SLICE_X98Y101_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X64Y100_SLICE_X97Y100_AQ),
.I3(1'b1),
.I4(CLBLM_R_X65Y100_SLICE_X99Y100_BQ),
.I5(1'b1),
.O5(CLBLM_R_X65Y101_SLICE_X98Y101_AO5),
.O6(CLBLM_R_X65Y101_SLICE_X98Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X65Y101_SLICE_X99Y101_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_BQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X65Y101_SLICE_X99Y101_AO6),
.Q(CLBLM_R_X65Y101_SLICE_X99Y101_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffddffddffdd55dd)
  ) CLBLM_R_X65Y101_SLICE_X99Y101_DLUT (
.I0(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I1(CLBLM_L_X64Y101_SLICE_X97Y101_B_XOR),
.I2(1'b1),
.I3(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I4(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I5(CLBLM_L_X64Y100_SLICE_X97Y100_BQ),
.O5(CLBLM_R_X65Y101_SLICE_X99Y101_DO5),
.O6(CLBLM_R_X65Y101_SLICE_X99Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h08cc00cc08cc00cc)
  ) CLBLM_R_X65Y101_SLICE_X99Y101_CLUT (
.I0(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I1(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I2(CLBLM_R_X65Y101_SLICE_X98Y101_B_XOR),
.I3(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I4(CLBLM_L_X60Y98_SLICE_X90Y98_AQ),
.I5(1'b1),
.O5(CLBLM_R_X65Y101_SLICE_X99Y101_CO5),
.O6(CLBLM_R_X65Y101_SLICE_X99Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h80008000fcfccccc)
  ) CLBLM_R_X65Y101_SLICE_X99Y101_BLUT (
.I0(CLBLM_L_X60Y98_SLICE_X90Y98_AQ),
.I1(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I2(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I3(CLBLM_R_X65Y101_SLICE_X98Y101_A_XOR),
.I4(CLBLM_L_X64Y101_SLICE_X97Y101_A_XOR),
.I5(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.O5(CLBLM_R_X65Y101_SLICE_X99Y101_BO5),
.O6(CLBLM_R_X65Y101_SLICE_X99Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3330000033302220)
  ) CLBLM_R_X65Y101_SLICE_X99Y101_ALUT (
.I0(CLBLM_R_X65Y101_SLICE_X99Y101_DO6),
.I1(CLBLM_R_X65Y97_SLICE_X99Y97_CO6),
.I2(CLBLM_L_X64Y101_SLICE_X96Y101_A_XOR),
.I3(CLBLM_R_X65Y97_SLICE_X98Y97_AO5),
.I4(CLBLM_R_X65Y97_SLICE_X98Y97_AO6),
.I5(CLBLM_R_X65Y101_SLICE_X99Y101_CO6),
.O5(CLBLM_R_X65Y101_SLICE_X99Y101_AO5),
.O6(CLBLM_R_X65Y101_SLICE_X99Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X65Y102_SLICE_X98Y102_CARRY4 (
.CI(CLBLM_R_X65Y101_SLICE_X98Y101_COUT),
.CO({CLBLM_R_X65Y102_SLICE_X98Y102_D_CY, CLBLM_R_X65Y102_SLICE_X98Y102_C_CY, CLBLM_R_X65Y102_SLICE_X98Y102_B_CY, CLBLM_R_X65Y102_SLICE_X98Y102_A_CY}),
.CYINIT(1'b0),
.DI({CLBLM_R_X65Y107_SLICE_X98Y107_AQ, CLBLM_R_X65Y107_SLICE_X98Y107_DQ, CLBLM_R_X63Y103_SLICE_X95Y103_CQ, CLBLM_R_X65Y102_SLICE_X98Y102_AO5}),
.O({CLBLM_R_X65Y102_SLICE_X98Y102_D_XOR, CLBLM_R_X65Y102_SLICE_X98Y102_C_XOR, CLBLM_R_X65Y102_SLICE_X98Y102_B_XOR, CLBLM_R_X65Y102_SLICE_X98Y102_A_XOR}),
.S({CLBLM_R_X65Y102_SLICE_X98Y102_DO6, CLBLM_R_X65Y102_SLICE_X98Y102_CO6, CLBLM_R_X65Y102_SLICE_X98Y102_BO6, CLBLM_R_X65Y102_SLICE_X98Y102_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa55555555)
  ) CLBLM_R_X65Y102_SLICE_X98Y102_DLUT (
.I0(CLBLM_R_X65Y107_SLICE_X98Y107_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X65Y107_SLICE_X98Y107_BQ),
.O5(CLBLM_R_X65Y102_SLICE_X98Y102_DO5),
.O6(CLBLM_R_X65Y102_SLICE_X98Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a5a5a5a5a5a5a5)
  ) CLBLM_R_X65Y102_SLICE_X98Y102_CLUT (
.I0(CLBLM_R_X65Y107_SLICE_X98Y107_AQ),
.I1(1'b1),
.I2(CLBLM_R_X65Y107_SLICE_X98Y107_DQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y102_SLICE_X98Y102_CO5),
.O6(CLBLM_R_X65Y102_SLICE_X98Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9999999999999999)
  ) CLBLM_R_X65Y102_SLICE_X98Y102_BLUT (
.I0(CLBLM_R_X65Y107_SLICE_X98Y107_DQ),
.I1(CLBLM_R_X63Y103_SLICE_X95Y103_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y102_SLICE_X98Y102_BO5),
.O6(CLBLM_R_X65Y102_SLICE_X98Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333cccc0000ffff)
  ) CLBLM_R_X65Y102_SLICE_X98Y102_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X63Y103_SLICE_X95Y103_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X62Y101_SLICE_X93Y101_CQ),
.I5(1'b1),
.O5(CLBLM_R_X65Y102_SLICE_X98Y102_AO5),
.O6(CLBLM_R_X65Y102_SLICE_X98Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X65Y102_SLICE_X99Y102_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_BQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X65Y102_SLICE_X99Y102_AO6),
.Q(CLBLM_R_X65Y102_SLICE_X99Y102_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y102_SLICE_X99Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y102_SLICE_X99Y102_DO5),
.O6(CLBLM_R_X65Y102_SLICE_X99Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h08aa08aa00aa00aa)
  ) CLBLM_R_X65Y102_SLICE_X99Y102_CLUT (
.I0(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I1(CLBLM_L_X60Y98_SLICE_X90Y98_AQ),
.I2(CLBLM_R_X65Y102_SLICE_X98Y102_B_XOR),
.I3(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I4(1'b1),
.I5(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.O5(CLBLM_R_X65Y102_SLICE_X99Y102_CO5),
.O6(CLBLM_R_X65Y102_SLICE_X99Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h22000000ffff0000)
  ) CLBLM_R_X65Y102_SLICE_X99Y102_BLUT (
.I0(CLBLM_L_X60Y98_SLICE_X90Y98_AQ),
.I1(CLBLM_R_X65Y102_SLICE_X98Y102_D_XOR),
.I2(1'b1),
.I3(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I4(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I5(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.O5(CLBLM_R_X65Y102_SLICE_X99Y102_BO5),
.O6(CLBLM_R_X65Y102_SLICE_X99Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5040504055445040)
  ) CLBLM_R_X65Y102_SLICE_X99Y102_ALUT (
.I0(CLBLM_L_X64Y99_SLICE_X97Y99_DO6),
.I1(CLBLM_L_X64Y102_SLICE_X96Y102_A_XOR),
.I2(CLBLM_R_X65Y97_SLICE_X98Y97_AO6),
.I3(CLBLM_R_X65Y97_SLICE_X98Y97_AO5),
.I4(CLBLM_R_X63Y102_SLICE_X95Y102_AO6),
.I5(CLBLM_R_X65Y102_SLICE_X99Y102_CO6),
.O5(CLBLM_R_X65Y102_SLICE_X99Y102_AO5),
.O6(CLBLM_R_X65Y102_SLICE_X99Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X65Y103_SLICE_X98Y103_CARRY4 (
.CI(CLBLM_R_X65Y102_SLICE_X98Y102_COUT),
.CO({CLBLM_R_X65Y103_SLICE_X98Y103_D_CY, CLBLM_R_X65Y103_SLICE_X98Y103_C_CY, CLBLM_R_X65Y103_SLICE_X98Y103_B_CY, CLBLM_R_X65Y103_SLICE_X98Y103_A_CY}),
.CYINIT(1'b0),
.DI({CLBLM_L_X64Y106_SLICE_X97Y106_AQ, CLBLM_R_X65Y106_SLICE_X98Y106_AQ, CLBLM_R_X65Y107_SLICE_X98Y107_CQ, CLBLM_R_X65Y107_SLICE_X98Y107_BQ}),
.O({CLBLM_R_X65Y103_SLICE_X98Y103_D_XOR, CLBLM_R_X65Y103_SLICE_X98Y103_C_XOR, CLBLM_R_X65Y103_SLICE_X98Y103_B_XOR, CLBLM_R_X65Y103_SLICE_X98Y103_A_XOR}),
.S({CLBLM_R_X65Y103_SLICE_X98Y103_DO6, CLBLM_R_X65Y103_SLICE_X98Y103_CO6, CLBLM_R_X65Y103_SLICE_X98Y103_BO6, CLBLM_R_X65Y103_SLICE_X98Y103_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a5a5a5a5a5a5a5)
  ) CLBLM_R_X65Y103_SLICE_X98Y103_DLUT (
.I0(CLBLM_R_X63Y103_SLICE_X95Y103_AQ),
.I1(1'b1),
.I2(CLBLM_L_X64Y106_SLICE_X97Y106_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y103_SLICE_X98Y103_DO5),
.O6(CLBLM_R_X65Y103_SLICE_X98Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00f0ff0f00f0f)
  ) CLBLM_R_X65Y103_SLICE_X98Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X65Y106_SLICE_X98Y106_AQ),
.I3(1'b1),
.I4(CLBLM_L_X64Y106_SLICE_X97Y106_AQ),
.I5(1'b1),
.O5(CLBLM_R_X65Y103_SLICE_X98Y103_CO5),
.O6(CLBLM_R_X65Y103_SLICE_X98Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a5a5a5a5a5a5a5)
  ) CLBLM_R_X65Y103_SLICE_X98Y103_BLUT (
.I0(CLBLM_R_X65Y107_SLICE_X98Y107_CQ),
.I1(1'b1),
.I2(CLBLM_R_X65Y106_SLICE_X98Y106_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y103_SLICE_X98Y103_BO5),
.O6(CLBLM_R_X65Y103_SLICE_X98Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa55aa55aa55aa55)
  ) CLBLM_R_X65Y103_SLICE_X98Y103_ALUT (
.I0(CLBLM_R_X65Y107_SLICE_X98Y107_CQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X65Y107_SLICE_X98Y107_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y103_SLICE_X98Y103_AO5),
.O6(CLBLM_R_X65Y103_SLICE_X98Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X65Y103_SLICE_X99Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_BQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X65Y103_SLICE_X99Y103_AO6),
.Q(CLBLM_R_X65Y103_SLICE_X99Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X65Y103_SLICE_X99Y103_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_BQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X65Y103_SLICE_X99Y103_BO6),
.Q(CLBLM_R_X65Y103_SLICE_X99Y103_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h08cc08cc00cc00cc)
  ) CLBLM_R_X65Y103_SLICE_X99Y103_DLUT (
.I0(CLBLM_L_X60Y98_SLICE_X90Y98_AQ),
.I1(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I2(CLBLM_R_X65Y103_SLICE_X98Y103_D_XOR),
.I3(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I4(1'b1),
.I5(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.O5(CLBLM_R_X65Y103_SLICE_X99Y103_DO5),
.O6(CLBLM_R_X65Y103_SLICE_X99Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2f002f000f000f00)
  ) CLBLM_R_X65Y103_SLICE_X99Y103_CLUT (
.I0(CLBLM_L_X60Y98_SLICE_X90Y98_AQ),
.I1(CLBLM_R_X65Y103_SLICE_X98Y103_C_XOR),
.I2(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I3(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I4(1'b1),
.I5(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.O5(CLBLM_R_X65Y103_SLICE_X99Y103_CO5),
.O6(CLBLM_R_X65Y103_SLICE_X99Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000f5c4f0c0)
  ) CLBLM_R_X65Y103_SLICE_X99Y103_BLUT (
.I0(CLBLM_R_X65Y103_SLICE_X99Y103_DO6),
.I1(CLBLM_L_X64Y103_SLICE_X96Y103_C_XOR),
.I2(CLBLM_R_X65Y97_SLICE_X98Y97_AO6),
.I3(CLBLM_R_X65Y97_SLICE_X98Y97_AO5),
.I4(CLBLM_R_X63Y103_SLICE_X95Y103_DO6),
.I5(CLBLM_R_X65Y97_SLICE_X99Y97_AO6),
.O5(CLBLM_R_X65Y103_SLICE_X99Y103_BO5),
.O6(CLBLM_R_X65Y103_SLICE_X99Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3030323230003200)
  ) CLBLM_R_X65Y103_SLICE_X99Y103_ALUT (
.I0(CLBLM_L_X64Y105_SLICE_X96Y105_CO6),
.I1(CLBLM_R_X63Y98_SLICE_X94Y98_DO6),
.I2(CLBLM_R_X65Y97_SLICE_X98Y97_AO6),
.I3(CLBLM_R_X65Y97_SLICE_X98Y97_AO5),
.I4(CLBLM_R_X65Y103_SLICE_X99Y103_CO6),
.I5(CLBLM_L_X64Y103_SLICE_X96Y103_B_XOR),
.O5(CLBLM_R_X65Y103_SLICE_X99Y103_AO5),
.O6(CLBLM_R_X65Y103_SLICE_X99Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X65Y104_SLICE_X98Y104_CARRY4 (
.CI(CLBLM_R_X65Y103_SLICE_X98Y103_COUT),
.CO({CLBLM_R_X65Y104_SLICE_X98Y104_D_CY, CLBLM_R_X65Y104_SLICE_X98Y104_C_CY, CLBLM_R_X65Y104_SLICE_X98Y104_B_CY, CLBLM_R_X65Y104_SLICE_X98Y104_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, CLBLM_R_X65Y106_SLICE_X98Y106_BQ, CLBLM_R_X63Y103_SLICE_X95Y103_AQ}),
.O({CLBLM_R_X65Y104_SLICE_X98Y104_D_XOR, CLBLM_R_X65Y104_SLICE_X98Y104_C_XOR, CLBLM_R_X65Y104_SLICE_X98Y104_B_XOR, CLBLM_R_X65Y104_SLICE_X98Y104_A_XOR}),
.S({CLBLM_R_X65Y104_SLICE_X98Y104_DO6, CLBLM_R_X65Y104_SLICE_X98Y104_CO6, CLBLM_R_X65Y104_SLICE_X98Y104_BO6, CLBLM_R_X65Y104_SLICE_X98Y104_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y104_SLICE_X98Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y104_SLICE_X98Y104_DO5),
.O6(CLBLM_R_X65Y104_SLICE_X98Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00f0ff0f00f0f)
  ) CLBLM_R_X65Y104_SLICE_X98Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X64Y106_SLICE_X97Y106_BQ),
.I3(1'b1),
.I4(CLBLM_L_X64Y106_SLICE_X97Y106_CQ),
.I5(1'b1),
.O5(CLBLM_R_X65Y104_SLICE_X98Y104_CO5),
.O6(CLBLM_R_X65Y104_SLICE_X98Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0000ff00ff)
  ) CLBLM_R_X65Y104_SLICE_X98Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X65Y106_SLICE_X98Y106_BQ),
.I4(1'b1),
.I5(CLBLM_L_X64Y106_SLICE_X97Y106_BQ),
.O5(CLBLM_R_X65Y104_SLICE_X98Y104_BO5),
.O6(CLBLM_R_X65Y104_SLICE_X98Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf00ff00ff00ff00f)
  ) CLBLM_R_X65Y104_SLICE_X98Y104_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X63Y103_SLICE_X95Y103_AQ),
.I3(CLBLM_R_X65Y106_SLICE_X98Y106_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y104_SLICE_X98Y104_AO5),
.O6(CLBLM_R_X65Y104_SLICE_X98Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X65Y104_SLICE_X99Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_BQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X65Y104_SLICE_X99Y104_AO6),
.Q(CLBLM_R_X65Y104_SLICE_X99Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X65Y104_SLICE_X99Y104_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_BQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X65Y104_SLICE_X99Y104_BO6),
.Q(CLBLM_R_X65Y104_SLICE_X99Y104_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h30ff00ff00000000)
  ) CLBLM_R_X65Y104_SLICE_X99Y104_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X65Y104_SLICE_X98Y104_A_XOR),
.I2(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I3(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I4(CLBLM_L_X60Y98_SLICE_X90Y98_AQ),
.I5(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.O5(CLBLM_R_X65Y104_SLICE_X99Y104_DO5),
.O6(CLBLM_R_X65Y104_SLICE_X99Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00aaa0aa00aa)
  ) CLBLM_R_X65Y104_SLICE_X99Y104_CLUT (
.I0(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I1(1'b1),
.I2(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I3(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I4(CLBLM_L_X60Y98_SLICE_X90Y98_AQ),
.I5(CLBLM_R_X65Y103_SLICE_X98Y103_A_XOR),
.O5(CLBLM_R_X65Y104_SLICE_X99Y104_CO5),
.O6(CLBLM_R_X65Y104_SLICE_X99Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3131303031003000)
  ) CLBLM_R_X65Y104_SLICE_X99Y104_BLUT (
.I0(CLBLM_R_X65Y104_SLICE_X99Y104_DO6),
.I1(CLBLM_R_X65Y97_SLICE_X98Y97_DO6),
.I2(CLBLM_R_X65Y97_SLICE_X98Y97_AO6),
.I3(CLBLM_L_X64Y103_SLICE_X96Y103_D_XOR),
.I4(CLBLM_R_X63Y104_SLICE_X95Y104_AO6),
.I5(CLBLM_R_X65Y97_SLICE_X98Y97_AO5),
.O5(CLBLM_R_X65Y104_SLICE_X99Y104_BO5),
.O6(CLBLM_R_X65Y104_SLICE_X99Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff002200f00020)
  ) CLBLM_R_X65Y104_SLICE_X99Y104_ALUT (
.I0(CLBLM_L_X64Y105_SLICE_X97Y105_CO6),
.I1(CLBLM_R_X65Y104_SLICE_X99Y104_CO6),
.I2(CLBLM_L_X64Y102_SLICE_X96Y102_D_XOR),
.I3(CLBLM_L_X62Y97_SLICE_X93Y97_DO6),
.I4(CLBLM_R_X65Y97_SLICE_X98Y97_AO6),
.I5(CLBLM_R_X65Y97_SLICE_X98Y97_AO5),
.O5(CLBLM_R_X65Y104_SLICE_X99Y104_AO5),
.O6(CLBLM_R_X65Y104_SLICE_X99Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X65Y105_SLICE_X98Y105_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_BQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X65Y105_SLICE_X98Y105_AO6),
.Q(CLBLM_R_X65Y105_SLICE_X98Y105_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X65Y105_SLICE_X98Y105_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_BQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X65Y105_SLICE_X98Y105_BO6),
.Q(CLBLM_R_X65Y105_SLICE_X98Y105_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaafffff0f0ffff)
  ) CLBLM_R_X65Y105_SLICE_X98Y105_DLUT (
.I0(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I1(1'b1),
.I2(CLBLM_L_X64Y104_SLICE_X97Y104_B_XOR),
.I3(CLBLM_R_X49Y107_SLICE_X75Y107_DQ),
.I4(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I5(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.O5(CLBLM_R_X65Y105_SLICE_X98Y105_DO5),
.O6(CLBLM_R_X65Y105_SLICE_X98Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbc8fffffbc8ffff)
  ) CLBLM_R_X65Y105_SLICE_X98Y105_CLUT (
.I0(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I1(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I2(CLBLM_R_X49Y106_SLICE_X75Y106_CQ),
.I3(CLBLM_L_X64Y103_SLICE_X97Y103_B_XOR),
.I4(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I5(1'b1),
.O5(CLBLM_R_X65Y105_SLICE_X98Y105_CO5),
.O6(CLBLM_R_X65Y105_SLICE_X98Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f000a0c0c0008)
  ) CLBLM_R_X65Y105_SLICE_X98Y105_BLUT (
.I0(CLBLM_R_X65Y105_SLICE_X98Y105_DO6),
.I1(CLBLM_R_X65Y97_SLICE_X98Y97_AO5),
.I2(CLBLM_R_X65Y99_SLICE_X98Y99_BO6),
.I3(CLBLM_R_X65Y105_SLICE_X99Y105_CO6),
.I4(CLBLM_R_X65Y97_SLICE_X98Y97_AO6),
.I5(CLBLM_L_X64Y104_SLICE_X96Y104_A_XOR),
.O5(CLBLM_R_X65Y105_SLICE_X98Y105_BO5),
.O6(CLBLM_R_X65Y105_SLICE_X98Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5151510050505000)
  ) CLBLM_R_X65Y105_SLICE_X98Y105_ALUT (
.I0(CLBLM_R_X65Y97_SLICE_X98Y97_CO6),
.I1(CLBLM_R_X65Y105_SLICE_X99Y105_BO6),
.I2(CLBLM_R_X65Y97_SLICE_X98Y97_AO6),
.I3(CLBLM_L_X64Y103_SLICE_X96Y103_A_XOR),
.I4(CLBLM_R_X65Y97_SLICE_X98Y97_AO5),
.I5(CLBLM_R_X65Y105_SLICE_X98Y105_CO6),
.O5(CLBLM_R_X65Y105_SLICE_X98Y105_AO5),
.O6(CLBLM_R_X65Y105_SLICE_X98Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X65Y105_SLICE_X99Y105_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X60Y98_SLICE_X91Y98_BQ),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X65Y105_SLICE_X99Y105_AO6),
.Q(CLBLM_R_X65Y105_SLICE_X99Y105_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cc00cc80cc80cc)
  ) CLBLM_R_X65Y105_SLICE_X99Y105_DLUT (
.I0(CLBLM_L_X60Y98_SLICE_X90Y98_AQ),
.I1(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I2(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I3(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I4(1'b1),
.I5(CLBLM_R_X65Y104_SLICE_X98Y104_C_XOR),
.O5(CLBLM_R_X65Y105_SLICE_X99Y105_DO5),
.O6(CLBLM_R_X65Y105_SLICE_X99Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h20ff20ff00000000)
  ) CLBLM_R_X65Y105_SLICE_X99Y105_CLUT (
.I0(CLBLM_L_X60Y98_SLICE_X90Y98_AQ),
.I1(CLBLM_R_X65Y104_SLICE_X98Y104_B_XOR),
.I2(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I3(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I4(1'b1),
.I5(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.O5(CLBLM_R_X65Y105_SLICE_X99Y105_CO5),
.O6(CLBLM_R_X65Y105_SLICE_X99Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7030303070303030)
  ) CLBLM_R_X65Y105_SLICE_X99Y105_BLUT (
.I0(CLBLM_R_X65Y103_SLICE_X98Y103_B_XOR),
.I1(CLBLM_L_X56Y97_SLICE_X84Y97_BQ),
.I2(CLBLM_L_X60Y97_SLICE_X90Y97_CQ),
.I3(CLBLM_L_X60Y97_SLICE_X90Y97_AQ),
.I4(CLBLM_L_X60Y98_SLICE_X90Y98_AQ),
.I5(1'b1),
.O5(CLBLM_R_X65Y105_SLICE_X99Y105_BO5),
.O6(CLBLM_R_X65Y105_SLICE_X99Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f500c400f000c0)
  ) CLBLM_R_X65Y105_SLICE_X99Y105_ALUT (
.I0(CLBLM_R_X65Y105_SLICE_X99Y105_DO6),
.I1(CLBLM_R_X65Y97_SLICE_X98Y97_AO5),
.I2(CLBLM_R_X65Y97_SLICE_X98Y97_AO6),
.I3(CLBLM_R_X65Y97_SLICE_X99Y97_BO6),
.I4(CLBLM_L_X64Y104_SLICE_X96Y104_B_XOR),
.I5(CLBLM_L_X64Y105_SLICE_X97Y105_DO6),
.O5(CLBLM_R_X65Y105_SLICE_X99Y105_AO5),
.O6(CLBLM_R_X65Y105_SLICE_X99Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X65Y106_SLICE_X98Y106_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y105_SLICE_X93Y105_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X65Y106_SLICE_X98Y106_AO6),
.Q(CLBLM_R_X65Y106_SLICE_X98Y106_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X65Y106_SLICE_X98Y106_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y105_SLICE_X93Y105_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X65Y106_SLICE_X98Y106_BO6),
.Q(CLBLM_R_X65Y106_SLICE_X98Y106_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X65Y106_SLICE_X98Y106_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y105_SLICE_X93Y105_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X65Y106_SLICE_X98Y106_CO6),
.Q(CLBLM_R_X65Y106_SLICE_X98Y106_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X65Y106_SLICE_X98Y106_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y105_SLICE_X93Y105_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X65Y106_SLICE_X98Y106_DO6),
.Q(CLBLM_R_X65Y106_SLICE_X98Y106_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h88228822f0f0f0f0)
  ) CLBLM_R_X65Y106_SLICE_X98Y106_DLUT (
.I0(CLBLM_R_X65Y101_SLICE_X99Y101_AQ),
.I1(CLBLL_R_X57Y103_SLICE_X86Y103_A5Q),
.I2(CLBLM_L_X64Y106_SLICE_X96Y106_AQ),
.I3(CLBLL_R_X57Y103_SLICE_X86Y103_AQ),
.I4(1'b1),
.I5(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.O5(CLBLM_R_X65Y106_SLICE_X98Y106_DO5),
.O6(CLBLM_R_X65Y106_SLICE_X98Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3c3caaaaaaaa)
  ) CLBLM_R_X65Y106_SLICE_X98Y106_CLUT (
.I0(CLBLM_L_X64Y105_SLICE_X97Y105_AQ),
.I1(CLBLL_R_X57Y103_SLICE_X86Y103_A5Q),
.I2(CLBLL_R_X57Y103_SLICE_X86Y103_AQ),
.I3(1'b1),
.I4(CLBLM_R_X65Y99_SLICE_X98Y99_AQ),
.I5(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.O5(CLBLM_R_X65Y106_SLICE_X98Y106_CO5),
.O6(CLBLM_R_X65Y106_SLICE_X98Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc3c30000aaaaaaaa)
  ) CLBLM_R_X65Y106_SLICE_X98Y106_BLUT (
.I0(CLBLM_L_X62Y103_SLICE_X93Y103_AQ),
.I1(CLBLL_R_X57Y103_SLICE_X86Y103_A5Q),
.I2(CLBLL_R_X57Y103_SLICE_X86Y103_AQ),
.I3(1'b1),
.I4(CLBLM_R_X65Y104_SLICE_X99Y104_BQ),
.I5(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.O5(CLBLM_R_X65Y106_SLICE_X98Y106_BO5),
.O6(CLBLM_R_X65Y106_SLICE_X98Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc330000f0f0f0f0)
  ) CLBLM_R_X65Y106_SLICE_X98Y106_ALUT (
.I0(1'b1),
.I1(CLBLL_R_X57Y103_SLICE_X86Y103_AQ),
.I2(CLBLM_R_X63Y110_SLICE_X94Y110_AQ),
.I3(CLBLL_R_X57Y103_SLICE_X86Y103_A5Q),
.I4(CLBLM_R_X65Y105_SLICE_X98Y105_AQ),
.I5(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.O5(CLBLM_R_X65Y106_SLICE_X98Y106_AO5),
.O6(CLBLM_R_X65Y106_SLICE_X98Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y106_SLICE_X99Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y106_SLICE_X99Y106_DO5),
.O6(CLBLM_R_X65Y106_SLICE_X99Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y106_SLICE_X99Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y106_SLICE_X99Y106_CO5),
.O6(CLBLM_R_X65Y106_SLICE_X99Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y106_SLICE_X99Y106_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y106_SLICE_X99Y106_BO5),
.O6(CLBLM_R_X65Y106_SLICE_X99Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y106_SLICE_X99Y106_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y106_SLICE_X99Y106_AO5),
.O6(CLBLM_R_X65Y106_SLICE_X99Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X65Y107_SLICE_X98Y107_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y105_SLICE_X93Y105_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X65Y107_SLICE_X98Y107_AO6),
.Q(CLBLM_R_X65Y107_SLICE_X98Y107_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X65Y107_SLICE_X98Y107_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y105_SLICE_X93Y105_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X65Y107_SLICE_X98Y107_BO6),
.Q(CLBLM_R_X65Y107_SLICE_X98Y107_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X65Y107_SLICE_X98Y107_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y105_SLICE_X93Y105_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X65Y107_SLICE_X98Y107_CO6),
.Q(CLBLM_R_X65Y107_SLICE_X98Y107_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(1)
  ) CLBLM_R_X65Y107_SLICE_X98Y107_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(CLBLM_L_X62Y105_SLICE_X93Y105_DO6),
.CLR(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.D(CLBLM_R_X65Y107_SLICE_X98Y107_DO6),
.Q(CLBLM_R_X65Y107_SLICE_X98Y107_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd580d58075207520)
  ) CLBLM_R_X65Y107_SLICE_X98Y107_DLUT (
.I0(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I1(CLBLL_R_X57Y103_SLICE_X86Y103_AQ),
.I2(CLBLM_R_X65Y102_SLICE_X99Y102_AQ),
.I3(CLBLM_L_X64Y107_SLICE_X96Y107_BQ),
.I4(1'b1),
.I5(CLBLL_R_X57Y103_SLICE_X86Y103_A5Q),
.O5(CLBLM_R_X65Y107_SLICE_X98Y107_DO5),
.O6(CLBLM_R_X65Y107_SLICE_X98Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8505072725050)
  ) CLBLM_R_X65Y107_SLICE_X98Y107_CLUT (
.I0(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I1(CLBLL_R_X57Y103_SLICE_X86Y103_AQ),
.I2(CLBLM_L_X64Y108_SLICE_X97Y108_AQ),
.I3(1'b1),
.I4(CLBLM_R_X65Y104_SLICE_X99Y104_AQ),
.I5(CLBLL_R_X57Y103_SLICE_X86Y103_A5Q),
.O5(CLBLM_R_X65Y107_SLICE_X98Y107_CO5),
.O6(CLBLM_R_X65Y107_SLICE_X98Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa55f0f00000f0f0)
  ) CLBLM_R_X65Y107_SLICE_X98Y107_BLUT (
.I0(CLBLL_R_X57Y103_SLICE_X86Y103_AQ),
.I1(1'b1),
.I2(CLBLM_L_X64Y108_SLICE_X96Y108_AQ),
.I3(CLBLL_R_X57Y103_SLICE_X86Y103_A5Q),
.I4(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I5(CLBLM_R_X65Y98_SLICE_X98Y98_AQ),
.O5(CLBLM_R_X65Y107_SLICE_X98Y107_BO5),
.O6(CLBLM_R_X65Y107_SLICE_X98Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h9090ffff90900000)
  ) CLBLM_R_X65Y107_SLICE_X98Y107_ALUT (
.I0(CLBLL_R_X57Y103_SLICE_X86Y103_AQ),
.I1(CLBLL_R_X57Y103_SLICE_X86Y103_A5Q),
.I2(CLBLM_L_X64Y99_SLICE_X96Y99_AQ),
.I3(1'b1),
.I4(CLBLM_L_X60Y98_SLICE_X91Y98_A5Q),
.I5(CLBLM_L_X64Y107_SLICE_X97Y107_AQ),
.O5(CLBLM_R_X65Y107_SLICE_X98Y107_AO5),
.O6(CLBLM_R_X65Y107_SLICE_X98Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y107_SLICE_X99Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y107_SLICE_X99Y107_DO5),
.O6(CLBLM_R_X65Y107_SLICE_X99Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y107_SLICE_X99Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y107_SLICE_X99Y107_CO5),
.O6(CLBLM_R_X65Y107_SLICE_X99Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y107_SLICE_X99Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y107_SLICE_X99Y107_BO5),
.O6(CLBLM_R_X65Y107_SLICE_X99Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X65Y107_SLICE_X99Y107_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X65Y107_SLICE_X99Y107_AO5),
.O6(CLBLM_R_X65Y107_SLICE_X99Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(RIOB33_X105Y127_IOB_X1Y128_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X139Y78_BUFHCE_X0Y20_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X139Y78_BUFHCE_X0Y20_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y101_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y101_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y102_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y102_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y103_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y103_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y104_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y104_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y105_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y105_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y106_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y106_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y107_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y107_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y108_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y108_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y109_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y109_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y110_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y110_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y111_IOB_X0Y111_IBUF (
.I(LIOB33_X0Y111_IOB_X0Y111_IPAD),
.O(LIOB33_X0Y111_IOB_X0Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y111_IOB_X0Y112_IBUF (
.I(LIOB33_X0Y111_IOB_X0Y112_IPAD),
.O(LIOB33_X0Y111_IOB_X0Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y113_IOB_X0Y113_IBUF (
.I(LIOB33_X0Y113_IOB_X0Y113_IPAD),
.O(LIOB33_X0Y113_IOB_X0Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y113_IOB_X0Y114_IBUF (
.I(LIOB33_X0Y113_IOB_X0Y114_IPAD),
.O(LIOB33_X0Y113_IOB_X0Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y115_IOB_X0Y115_IBUF (
.I(LIOB33_X0Y115_IOB_X0Y115_IPAD),
.O(LIOB33_X0Y115_IOB_X0Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y115_IOB_X0Y116_IBUF (
.I(LIOB33_X0Y115_IOB_X0Y116_IPAD),
.O(LIOB33_X0Y115_IOB_X0Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y117_IOB_X0Y117_IBUF (
.I(LIOB33_X0Y117_IOB_X0Y117_IPAD),
.O(LIOB33_X0Y117_IOB_X0Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y117_IOB_X0Y118_IBUF (
.I(LIOB33_X0Y117_IOB_X0Y118_IPAD),
.O(LIOB33_X0Y117_IOB_X0Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y119_IOB_X0Y119_IBUF (
.I(LIOB33_X0Y119_IOB_X0Y119_IPAD),
.O(LIOB33_X0Y119_IOB_X0Y119_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y119_IOB_X0Y120_IBUF (
.I(LIOB33_X0Y119_IOB_X0Y120_IPAD),
.O(LIOB33_X0Y119_IOB_X0Y120_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y121_IOB_X0Y121_IBUF (
.I(LIOB33_X0Y121_IOB_X0Y121_IPAD),
.O(LIOB33_X0Y121_IOB_X0Y121_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y121_IOB_X0Y122_IBUF (
.I(LIOB33_X0Y121_IOB_X0Y122_IPAD),
.O(LIOB33_X0Y121_IOB_X0Y122_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y123_IOB_X0Y123_IBUF (
.I(LIOB33_X0Y123_IOB_X0Y123_IPAD),
.O(LIOB33_X0Y123_IOB_X0Y123_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y124_OBUF (
.I(CLBLM_R_X49Y109_SLICE_X74Y109_DQ),
.O(LIOB33_X0Y123_IOB_X0Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y125_OBUF (
.I(CLBLM_R_X49Y107_SLICE_X74Y107_AQ),
.O(LIOB33_X0Y125_IOB_X0Y125_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y126_OBUF (
.I(CLBLM_R_X49Y111_SLICE_X74Y111_AQ),
.O(LIOB33_X0Y125_IOB_X0Y126_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y127_OBUF (
.I(CLBLM_R_X49Y111_SLICE_X74Y111_BQ),
.O(LIOB33_X0Y127_IOB_X0Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y128_OBUF (
.I(CLBLM_R_X49Y109_SLICE_X74Y109_AQ),
.O(LIOB33_X0Y127_IOB_X0Y128_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y129_OBUF (
.I(CLBLM_R_X49Y109_SLICE_X74Y109_BQ),
.O(LIOB33_X0Y129_IOB_X0Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y130_OBUF (
.I(CLBLM_R_X49Y111_SLICE_X74Y111_CQ),
.O(LIOB33_X0Y129_IOB_X0Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y131_OBUF (
.I(CLBLM_R_X49Y109_SLICE_X74Y109_CQ),
.O(LIOB33_X0Y131_IOB_X0Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y132_OBUF (
.I(CLBLM_R_X49Y109_SLICE_X74Y109_DQ),
.O(LIOB33_X0Y131_IOB_X0Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y133_OBUF (
.I(CLBLM_R_X49Y107_SLICE_X74Y107_AQ),
.O(LIOB33_X0Y133_IOB_X0Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y134_OBUF (
.I(CLBLM_R_X49Y111_SLICE_X74Y111_AQ),
.O(LIOB33_X0Y133_IOB_X0Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y135_OBUF (
.I(CLBLM_R_X49Y111_SLICE_X74Y111_BQ),
.O(LIOB33_X0Y135_IOB_X0Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y136_OBUF (
.I(CLBLM_R_X49Y109_SLICE_X74Y109_AQ),
.O(LIOB33_X0Y135_IOB_X0Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y137_OBUF (
.I(CLBLM_R_X49Y109_SLICE_X74Y109_BQ),
.O(LIOB33_X0Y137_IOB_X0Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y138_OBUF (
.I(CLBLM_R_X49Y111_SLICE_X74Y111_CQ),
.O(LIOB33_X0Y137_IOB_X0Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y139_OBUF (
.I(CLBLM_R_X49Y109_SLICE_X74Y109_CQ),
.O(LIOB33_X0Y139_IOB_X0Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y140_OBUF (
.I(CLBLM_L_X50Y104_SLICE_X76Y104_AQ),
.O(LIOB33_X0Y139_IOB_X0Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y141_OBUF (
.I(CLBLM_L_X50Y105_SLICE_X77Y105_AQ),
.O(LIOB33_X0Y141_IOB_X0Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y142_OBUF (
.I(CLBLM_R_X49Y105_SLICE_X75Y105_CQ),
.O(LIOB33_X0Y141_IOB_X0Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y143_IOB_X0Y143_OBUF (
.I(CLBLM_R_X49Y106_SLICE_X74Y106_AQ),
.O(LIOB33_X0Y143_IOB_X0Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y145_OBUF (
.I(CLBLM_L_X50Y106_SLICE_X76Y106_CQ),
.O(LIOB33_X0Y145_IOB_X0Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y146_OBUF (
.I(CLBLM_L_X50Y107_SLICE_X76Y107_BQ),
.O(LIOB33_X0Y145_IOB_X0Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y147_OBUF (
.I(CLBLM_L_X50Y107_SLICE_X77Y107_AQ),
.O(LIOB33_X0Y147_IOB_X0Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y148_OBUF (
.I(CLBLM_R_X49Y111_SLICE_X75Y111_AQ),
.O(LIOB33_X0Y147_IOB_X0Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y100_IOB_X0Y100_IBUF (
.I(LIOB33_SING_X0Y100_IOB_X0Y100_IPAD),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y149_IOB_X0Y149_OBUF (
.I(CLBLM_R_X49Y111_SLICE_X75Y111_A5Q),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y101_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y102_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y103_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y104_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y105_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y105_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y106_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y107_IOB_X1Y107_OBUF (
.I(1'b0),
.O(RIOB33_X105Y107_IOB_X1Y107_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y107_IOB_X1Y108_OBUF (
.I(CLBLM_R_X65Y100_SLICE_X99Y100_CQ),
.O(RIOB33_X105Y107_IOB_X1Y108_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y109_IOB_X1Y109_OBUF (
.I(CLBLM_R_X65Y100_SLICE_X99Y100_AQ),
.O(RIOB33_X105Y109_IOB_X1Y109_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y109_IOB_X1Y110_OBUF (
.I(CLBLM_R_X65Y106_SLICE_X98Y106_CQ),
.O(RIOB33_X105Y109_IOB_X1Y110_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y111_IOB_X1Y111_OBUF (
.I(CLBLM_L_X64Y106_SLICE_X97Y106_DQ),
.O(RIOB33_X105Y111_IOB_X1Y111_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y111_IOB_X1Y112_OBUF (
.I(CLBLM_R_X65Y100_SLICE_X99Y100_BQ),
.O(RIOB33_X105Y111_IOB_X1Y112_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y113_IOB_X1Y113_OBUF (
.I(CLBLM_R_X65Y106_SLICE_X98Y106_DQ),
.O(RIOB33_X105Y113_IOB_X1Y113_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y113_IOB_X1Y114_OBUF (
.I(CLBLM_R_X63Y103_SLICE_X95Y103_BQ),
.O(RIOB33_X105Y113_IOB_X1Y114_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y115_IOB_X1Y115_OBUF (
.I(CLBLM_R_X63Y101_SLICE_X95Y101_AQ),
.O(RIOB33_X105Y115_IOB_X1Y115_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y115_IOB_X1Y116_OBUF (
.I(CLBLM_R_X63Y103_SLICE_X95Y103_CQ),
.O(RIOB33_X105Y115_IOB_X1Y116_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y117_IOB_X1Y117_OBUF (
.I(CLBLM_R_X65Y107_SLICE_X98Y107_DQ),
.O(RIOB33_X105Y117_IOB_X1Y117_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y117_IOB_X1Y118_OBUF (
.I(CLBLM_R_X65Y107_SLICE_X98Y107_AQ),
.O(RIOB33_X105Y117_IOB_X1Y118_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y119_IOB_X1Y119_OBUF (
.I(CLBLM_R_X65Y107_SLICE_X98Y107_BQ),
.O(RIOB33_X105Y119_IOB_X1Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y119_IOB_X1Y120_OBUF (
.I(CLBLM_R_X65Y107_SLICE_X98Y107_CQ),
.O(RIOB33_X105Y119_IOB_X1Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y121_IOB_X1Y121_OBUF (
.I(CLBLM_R_X65Y106_SLICE_X98Y106_AQ),
.O(RIOB33_X105Y121_IOB_X1Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y121_IOB_X1Y122_OBUF (
.I(CLBLM_L_X64Y106_SLICE_X97Y106_AQ),
.O(RIOB33_X105Y121_IOB_X1Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y123_IOB_X1Y123_OBUF (
.I(CLBLM_R_X63Y103_SLICE_X95Y103_AQ),
.O(RIOB33_X105Y123_IOB_X1Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y123_IOB_X1Y124_OBUF (
.I(CLBLM_R_X65Y106_SLICE_X98Y106_BQ),
.O(RIOB33_X105Y123_IOB_X1Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y125_IOB_X1Y125_OBUF (
.I(CLBLM_L_X64Y106_SLICE_X97Y106_BQ),
.O(RIOB33_X105Y125_IOB_X1Y125_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y125_IOB_X1Y126_OBUF (
.I(CLBLM_L_X64Y106_SLICE_X97Y106_CQ),
.O(RIOB33_X105Y125_IOB_X1Y126_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y127_IOB_X1Y127_OBUF (
.I(CLBLM_R_X59Y102_SLICE_X88Y102_AQ),
.O(RIOB33_X105Y127_IOB_X1Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y128_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y129_IOB_X1Y129_OBUF (
.I(CLBLM_L_X62Y104_SLICE_X93Y104_AQ),
.O(RIOB33_X105Y129_IOB_X1Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y129_IOB_X1Y130_OBUF (
.I(CLBLM_L_X62Y103_SLICE_X92Y103_AQ),
.O(RIOB33_X105Y129_IOB_X1Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y131_IOB_X1Y131_OBUF (
.I(CLBLM_R_X59Y102_SLICE_X89Y102_AQ),
.O(RIOB33_X105Y131_IOB_X1Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y131_IOB_X1Y132_OBUF (
.I(CLBLM_L_X60Y110_SLICE_X91Y110_AQ),
.O(RIOB33_X105Y131_IOB_X1Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y133_IOB_X1Y133_OBUF (
.I(CLBLM_L_X62Y106_SLICE_X93Y106_AQ),
.O(RIOB33_X105Y133_IOB_X1Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y133_IOB_X1Y134_OBUF (
.I(CLBLM_L_X62Y110_SLICE_X92Y110_AQ),
.O(RIOB33_X105Y133_IOB_X1Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y135_IOB_X1Y135_OBUF (
.I(CLBLM_L_X62Y108_SLICE_X93Y108_AQ),
.O(RIOB33_X105Y135_IOB_X1Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y135_IOB_X1Y136_OBUF (
.I(CLBLM_L_X60Y111_SLICE_X91Y111_BQ),
.O(RIOB33_X105Y135_IOB_X1Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y137_IOB_X1Y137_OBUF (
.I(CLBLM_L_X60Y111_SLICE_X90Y111_AQ),
.O(RIOB33_X105Y137_IOB_X1Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y137_IOB_X1Y138_OBUF (
.I(CLBLM_L_X62Y110_SLICE_X92Y110_BQ),
.O(RIOB33_X105Y137_IOB_X1Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y139_IOB_X1Y139_OBUF (
.I(CLBLM_L_X60Y111_SLICE_X91Y111_AQ),
.O(RIOB33_X105Y139_IOB_X1Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y139_IOB_X1Y140_OBUF (
.I(CLBLL_R_X57Y99_SLICE_X87Y99_AQ),
.O(RIOB33_X105Y139_IOB_X1Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y141_IOB_X1Y141_OBUF (
.I(CLBLM_L_X60Y98_SLICE_X90Y98_BQ),
.O(RIOB33_X105Y141_IOB_X1Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y141_IOB_X1Y142_OBUF (
.I(CLBLM_L_X62Y110_SLICE_X93Y110_AQ),
.O(RIOB33_X105Y141_IOB_X1Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y143_IOB_X1Y143_OBUF (
.I(CLBLM_L_X56Y111_SLICE_X84Y111_AQ),
.O(RIOB33_X105Y143_IOB_X1Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y143_IOB_X1Y144_OBUF (
.I(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.O(RIOB33_X105Y143_IOB_X1Y144_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y145_IOB_X1Y145_OBUF (
.I(CLBLL_L_X54Y109_SLICE_X82Y109_AO6),
.O(RIOB33_X105Y145_IOB_X1Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y100_IOB_X1Y100_IBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_IPAD),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_I)
  );
  assign CLBLL_L_X52Y99_SLICE_X78Y99_A = CLBLL_L_X52Y99_SLICE_X78Y99_AO6;
  assign CLBLL_L_X52Y99_SLICE_X78Y99_B = CLBLL_L_X52Y99_SLICE_X78Y99_BO6;
  assign CLBLL_L_X52Y99_SLICE_X78Y99_C = CLBLL_L_X52Y99_SLICE_X78Y99_CO6;
  assign CLBLL_L_X52Y99_SLICE_X78Y99_D = CLBLL_L_X52Y99_SLICE_X78Y99_DO6;
  assign CLBLL_L_X52Y99_SLICE_X79Y99_A = CLBLL_L_X52Y99_SLICE_X79Y99_AO6;
  assign CLBLL_L_X52Y99_SLICE_X79Y99_B = CLBLL_L_X52Y99_SLICE_X79Y99_BO6;
  assign CLBLL_L_X52Y99_SLICE_X79Y99_C = CLBLL_L_X52Y99_SLICE_X79Y99_CO6;
  assign CLBLL_L_X52Y99_SLICE_X79Y99_D = CLBLL_L_X52Y99_SLICE_X79Y99_DO6;
  assign CLBLL_L_X52Y99_SLICE_X79Y99_AMUX = CLBLL_L_X52Y99_SLICE_X79Y99_AO6;
  assign CLBLL_L_X52Y101_SLICE_X78Y101_A = CLBLL_L_X52Y101_SLICE_X78Y101_AO6;
  assign CLBLL_L_X52Y101_SLICE_X78Y101_B = CLBLL_L_X52Y101_SLICE_X78Y101_BO6;
  assign CLBLL_L_X52Y101_SLICE_X78Y101_C = CLBLL_L_X52Y101_SLICE_X78Y101_CO6;
  assign CLBLL_L_X52Y101_SLICE_X78Y101_D = CLBLL_L_X52Y101_SLICE_X78Y101_DO6;
  assign CLBLL_L_X52Y101_SLICE_X79Y101_A = CLBLL_L_X52Y101_SLICE_X79Y101_AO6;
  assign CLBLL_L_X52Y101_SLICE_X79Y101_B = CLBLL_L_X52Y101_SLICE_X79Y101_BO6;
  assign CLBLL_L_X52Y101_SLICE_X79Y101_C = CLBLL_L_X52Y101_SLICE_X79Y101_CO6;
  assign CLBLL_L_X52Y101_SLICE_X79Y101_D = CLBLL_L_X52Y101_SLICE_X79Y101_DO6;
  assign CLBLL_L_X52Y105_SLICE_X78Y105_A = CLBLL_L_X52Y105_SLICE_X78Y105_AO6;
  assign CLBLL_L_X52Y105_SLICE_X78Y105_B = CLBLL_L_X52Y105_SLICE_X78Y105_BO6;
  assign CLBLL_L_X52Y105_SLICE_X78Y105_C = CLBLL_L_X52Y105_SLICE_X78Y105_CO6;
  assign CLBLL_L_X52Y105_SLICE_X78Y105_D = CLBLL_L_X52Y105_SLICE_X78Y105_DO6;
  assign CLBLL_L_X52Y105_SLICE_X78Y105_AMUX = CLBLL_L_X52Y105_SLICE_X78Y105_AO5;
  assign CLBLL_L_X52Y105_SLICE_X78Y105_BMUX = CLBLL_L_X52Y105_SLICE_X78Y105_BO5;
  assign CLBLL_L_X52Y105_SLICE_X79Y105_A = CLBLL_L_X52Y105_SLICE_X79Y105_AO6;
  assign CLBLL_L_X52Y105_SLICE_X79Y105_B = CLBLL_L_X52Y105_SLICE_X79Y105_BO6;
  assign CLBLL_L_X52Y105_SLICE_X79Y105_C = CLBLL_L_X52Y105_SLICE_X79Y105_CO6;
  assign CLBLL_L_X52Y105_SLICE_X79Y105_D = CLBLL_L_X52Y105_SLICE_X79Y105_DO6;
  assign CLBLL_L_X52Y106_SLICE_X78Y106_A = CLBLL_L_X52Y106_SLICE_X78Y106_AO6;
  assign CLBLL_L_X52Y106_SLICE_X78Y106_B = CLBLL_L_X52Y106_SLICE_X78Y106_BO6;
  assign CLBLL_L_X52Y106_SLICE_X78Y106_C = CLBLL_L_X52Y106_SLICE_X78Y106_CO6;
  assign CLBLL_L_X52Y106_SLICE_X78Y106_D = CLBLL_L_X52Y106_SLICE_X78Y106_DO6;
  assign CLBLL_L_X52Y106_SLICE_X78Y106_AMUX = CLBLL_L_X52Y106_SLICE_X78Y106_AO5;
  assign CLBLL_L_X52Y106_SLICE_X79Y106_A = CLBLL_L_X52Y106_SLICE_X79Y106_AO6;
  assign CLBLL_L_X52Y106_SLICE_X79Y106_B = CLBLL_L_X52Y106_SLICE_X79Y106_BO6;
  assign CLBLL_L_X52Y106_SLICE_X79Y106_C = CLBLL_L_X52Y106_SLICE_X79Y106_CO6;
  assign CLBLL_L_X52Y106_SLICE_X79Y106_D = CLBLL_L_X52Y106_SLICE_X79Y106_DO6;
  assign CLBLL_L_X52Y106_SLICE_X79Y106_AMUX = CLBLL_L_X52Y106_SLICE_X79Y106_AO5;
  assign CLBLL_L_X52Y107_SLICE_X78Y107_A = CLBLL_L_X52Y107_SLICE_X78Y107_AO6;
  assign CLBLL_L_X52Y107_SLICE_X78Y107_B = CLBLL_L_X52Y107_SLICE_X78Y107_BO6;
  assign CLBLL_L_X52Y107_SLICE_X78Y107_C = CLBLL_L_X52Y107_SLICE_X78Y107_CO6;
  assign CLBLL_L_X52Y107_SLICE_X78Y107_D = CLBLL_L_X52Y107_SLICE_X78Y107_DO6;
  assign CLBLL_L_X52Y107_SLICE_X78Y107_AMUX = CLBLL_L_X52Y107_SLICE_X78Y107_AO5;
  assign CLBLL_L_X52Y107_SLICE_X78Y107_BMUX = CLBLL_L_X52Y107_SLICE_X78Y107_BO5;
  assign CLBLL_L_X52Y107_SLICE_X79Y107_A = CLBLL_L_X52Y107_SLICE_X79Y107_AO6;
  assign CLBLL_L_X52Y107_SLICE_X79Y107_B = CLBLL_L_X52Y107_SLICE_X79Y107_BO6;
  assign CLBLL_L_X52Y107_SLICE_X79Y107_C = CLBLL_L_X52Y107_SLICE_X79Y107_CO6;
  assign CLBLL_L_X52Y107_SLICE_X79Y107_D = CLBLL_L_X52Y107_SLICE_X79Y107_DO6;
  assign CLBLL_L_X54Y97_SLICE_X82Y97_A = CLBLL_L_X54Y97_SLICE_X82Y97_AO6;
  assign CLBLL_L_X54Y97_SLICE_X82Y97_B = CLBLL_L_X54Y97_SLICE_X82Y97_BO6;
  assign CLBLL_L_X54Y97_SLICE_X82Y97_C = CLBLL_L_X54Y97_SLICE_X82Y97_CO6;
  assign CLBLL_L_X54Y97_SLICE_X82Y97_D = CLBLL_L_X54Y97_SLICE_X82Y97_DO6;
  assign CLBLL_L_X54Y97_SLICE_X83Y97_A = CLBLL_L_X54Y97_SLICE_X83Y97_AO6;
  assign CLBLL_L_X54Y97_SLICE_X83Y97_B = CLBLL_L_X54Y97_SLICE_X83Y97_BO6;
  assign CLBLL_L_X54Y97_SLICE_X83Y97_C = CLBLL_L_X54Y97_SLICE_X83Y97_CO6;
  assign CLBLL_L_X54Y97_SLICE_X83Y97_D = CLBLL_L_X54Y97_SLICE_X83Y97_DO6;
  assign CLBLL_L_X54Y98_SLICE_X82Y98_A = CLBLL_L_X54Y98_SLICE_X82Y98_AO6;
  assign CLBLL_L_X54Y98_SLICE_X82Y98_B = CLBLL_L_X54Y98_SLICE_X82Y98_BO6;
  assign CLBLL_L_X54Y98_SLICE_X82Y98_C = CLBLL_L_X54Y98_SLICE_X82Y98_CO6;
  assign CLBLL_L_X54Y98_SLICE_X82Y98_D = CLBLL_L_X54Y98_SLICE_X82Y98_DO6;
  assign CLBLL_L_X54Y98_SLICE_X82Y98_BMUX = CLBLL_L_X54Y98_SLICE_X82Y98_BO6;
  assign CLBLL_L_X54Y98_SLICE_X83Y98_A = CLBLL_L_X54Y98_SLICE_X83Y98_AO6;
  assign CLBLL_L_X54Y98_SLICE_X83Y98_B = CLBLL_L_X54Y98_SLICE_X83Y98_BO6;
  assign CLBLL_L_X54Y98_SLICE_X83Y98_C = CLBLL_L_X54Y98_SLICE_X83Y98_CO6;
  assign CLBLL_L_X54Y98_SLICE_X83Y98_D = CLBLL_L_X54Y98_SLICE_X83Y98_DO6;
  assign CLBLL_L_X54Y98_SLICE_X83Y98_CMUX = CLBLL_L_X54Y98_SLICE_X83Y98_CO5;
  assign CLBLL_L_X54Y99_SLICE_X82Y99_A = CLBLL_L_X54Y99_SLICE_X82Y99_AO6;
  assign CLBLL_L_X54Y99_SLICE_X82Y99_B = CLBLL_L_X54Y99_SLICE_X82Y99_BO6;
  assign CLBLL_L_X54Y99_SLICE_X82Y99_C = CLBLL_L_X54Y99_SLICE_X82Y99_CO6;
  assign CLBLL_L_X54Y99_SLICE_X82Y99_D = CLBLL_L_X54Y99_SLICE_X82Y99_DO6;
  assign CLBLL_L_X54Y99_SLICE_X82Y99_AMUX = CLBLL_L_X54Y99_SLICE_X82Y99_AO5;
  assign CLBLL_L_X54Y99_SLICE_X82Y99_BMUX = CLBLL_L_X54Y99_SLICE_X82Y99_BO5;
  assign CLBLL_L_X54Y99_SLICE_X83Y99_A = CLBLL_L_X54Y99_SLICE_X83Y99_AO6;
  assign CLBLL_L_X54Y99_SLICE_X83Y99_B = CLBLL_L_X54Y99_SLICE_X83Y99_BO6;
  assign CLBLL_L_X54Y99_SLICE_X83Y99_C = CLBLL_L_X54Y99_SLICE_X83Y99_CO6;
  assign CLBLL_L_X54Y99_SLICE_X83Y99_D = CLBLL_L_X54Y99_SLICE_X83Y99_DO6;
  assign CLBLL_L_X54Y99_SLICE_X83Y99_AMUX = CLBLL_L_X54Y99_SLICE_X83Y99_A5Q;
  assign CLBLL_L_X54Y99_SLICE_X83Y99_BMUX = CLBLL_L_X54Y99_SLICE_X83Y99_BO5;
  assign CLBLL_L_X54Y100_SLICE_X82Y100_A = CLBLL_L_X54Y100_SLICE_X82Y100_AO6;
  assign CLBLL_L_X54Y100_SLICE_X82Y100_B = CLBLL_L_X54Y100_SLICE_X82Y100_BO6;
  assign CLBLL_L_X54Y100_SLICE_X82Y100_C = CLBLL_L_X54Y100_SLICE_X82Y100_CO6;
  assign CLBLL_L_X54Y100_SLICE_X82Y100_D = CLBLL_L_X54Y100_SLICE_X82Y100_DO6;
  assign CLBLL_L_X54Y100_SLICE_X82Y100_AMUX = CLBLL_L_X54Y100_SLICE_X82Y100_AO5;
  assign CLBLL_L_X54Y100_SLICE_X83Y100_A = CLBLL_L_X54Y100_SLICE_X83Y100_AO6;
  assign CLBLL_L_X54Y100_SLICE_X83Y100_B = CLBLL_L_X54Y100_SLICE_X83Y100_BO6;
  assign CLBLL_L_X54Y100_SLICE_X83Y100_C = CLBLL_L_X54Y100_SLICE_X83Y100_CO6;
  assign CLBLL_L_X54Y100_SLICE_X83Y100_D = CLBLL_L_X54Y100_SLICE_X83Y100_DO6;
  assign CLBLL_L_X54Y100_SLICE_X83Y100_AMUX = CLBLL_L_X54Y100_SLICE_X83Y100_AO5;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_A = CLBLL_L_X54Y101_SLICE_X82Y101_AO6;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_B = CLBLL_L_X54Y101_SLICE_X82Y101_BO6;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_C = CLBLL_L_X54Y101_SLICE_X82Y101_CO6;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_D = CLBLL_L_X54Y101_SLICE_X82Y101_DO6;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_AMUX = CLBLL_L_X54Y101_SLICE_X82Y101_AO5;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_A = CLBLL_L_X54Y101_SLICE_X83Y101_AO6;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_B = CLBLL_L_X54Y101_SLICE_X83Y101_BO6;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_C = CLBLL_L_X54Y101_SLICE_X83Y101_CO6;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_D = CLBLL_L_X54Y101_SLICE_X83Y101_DO6;
  assign CLBLL_L_X54Y102_SLICE_X82Y102_A = CLBLL_L_X54Y102_SLICE_X82Y102_AO6;
  assign CLBLL_L_X54Y102_SLICE_X82Y102_B = CLBLL_L_X54Y102_SLICE_X82Y102_BO6;
  assign CLBLL_L_X54Y102_SLICE_X82Y102_C = CLBLL_L_X54Y102_SLICE_X82Y102_CO6;
  assign CLBLL_L_X54Y102_SLICE_X82Y102_D = CLBLL_L_X54Y102_SLICE_X82Y102_DO6;
  assign CLBLL_L_X54Y102_SLICE_X82Y102_AMUX = CLBLL_L_X54Y102_SLICE_X82Y102_AO5;
  assign CLBLL_L_X54Y102_SLICE_X83Y102_A = CLBLL_L_X54Y102_SLICE_X83Y102_AO6;
  assign CLBLL_L_X54Y102_SLICE_X83Y102_B = CLBLL_L_X54Y102_SLICE_X83Y102_BO6;
  assign CLBLL_L_X54Y102_SLICE_X83Y102_C = CLBLL_L_X54Y102_SLICE_X83Y102_CO6;
  assign CLBLL_L_X54Y102_SLICE_X83Y102_D = CLBLL_L_X54Y102_SLICE_X83Y102_DO6;
  assign CLBLL_L_X54Y103_SLICE_X82Y103_A = CLBLL_L_X54Y103_SLICE_X82Y103_AO6;
  assign CLBLL_L_X54Y103_SLICE_X82Y103_B = CLBLL_L_X54Y103_SLICE_X82Y103_BO6;
  assign CLBLL_L_X54Y103_SLICE_X82Y103_C = CLBLL_L_X54Y103_SLICE_X82Y103_CO6;
  assign CLBLL_L_X54Y103_SLICE_X82Y103_D = CLBLL_L_X54Y103_SLICE_X82Y103_DO6;
  assign CLBLL_L_X54Y103_SLICE_X83Y103_A = CLBLL_L_X54Y103_SLICE_X83Y103_AO6;
  assign CLBLL_L_X54Y103_SLICE_X83Y103_B = CLBLL_L_X54Y103_SLICE_X83Y103_BO6;
  assign CLBLL_L_X54Y103_SLICE_X83Y103_C = CLBLL_L_X54Y103_SLICE_X83Y103_CO6;
  assign CLBLL_L_X54Y103_SLICE_X83Y103_D = CLBLL_L_X54Y103_SLICE_X83Y103_DO6;
  assign CLBLL_L_X54Y104_SLICE_X82Y104_A = CLBLL_L_X54Y104_SLICE_X82Y104_AO6;
  assign CLBLL_L_X54Y104_SLICE_X82Y104_B = CLBLL_L_X54Y104_SLICE_X82Y104_BO6;
  assign CLBLL_L_X54Y104_SLICE_X82Y104_C = CLBLL_L_X54Y104_SLICE_X82Y104_CO6;
  assign CLBLL_L_X54Y104_SLICE_X82Y104_D = CLBLL_L_X54Y104_SLICE_X82Y104_DO6;
  assign CLBLL_L_X54Y104_SLICE_X83Y104_A = CLBLL_L_X54Y104_SLICE_X83Y104_AO6;
  assign CLBLL_L_X54Y104_SLICE_X83Y104_B = CLBLL_L_X54Y104_SLICE_X83Y104_BO6;
  assign CLBLL_L_X54Y104_SLICE_X83Y104_C = CLBLL_L_X54Y104_SLICE_X83Y104_CO6;
  assign CLBLL_L_X54Y104_SLICE_X83Y104_D = CLBLL_L_X54Y104_SLICE_X83Y104_DO6;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_A = CLBLL_L_X54Y105_SLICE_X82Y105_AO6;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_B = CLBLL_L_X54Y105_SLICE_X82Y105_BO6;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_C = CLBLL_L_X54Y105_SLICE_X82Y105_CO6;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_D = CLBLL_L_X54Y105_SLICE_X82Y105_DO6;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_BMUX = CLBLL_L_X54Y105_SLICE_X82Y105_B_XOR;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_CMUX = CLBLL_L_X54Y105_SLICE_X82Y105_C_XOR;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_DMUX = CLBLL_L_X54Y105_SLICE_X82Y105_D_XOR;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_A = CLBLL_L_X54Y105_SLICE_X83Y105_AO6;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_B = CLBLL_L_X54Y105_SLICE_X83Y105_BO6;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_C = CLBLL_L_X54Y105_SLICE_X83Y105_CO6;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_D = CLBLL_L_X54Y105_SLICE_X83Y105_DO6;
  assign CLBLL_L_X54Y106_SLICE_X82Y106_A = CLBLL_L_X54Y106_SLICE_X82Y106_AO6;
  assign CLBLL_L_X54Y106_SLICE_X82Y106_B = CLBLL_L_X54Y106_SLICE_X82Y106_BO6;
  assign CLBLL_L_X54Y106_SLICE_X82Y106_C = CLBLL_L_X54Y106_SLICE_X82Y106_CO6;
  assign CLBLL_L_X54Y106_SLICE_X82Y106_D = CLBLL_L_X54Y106_SLICE_X82Y106_DO6;
  assign CLBLL_L_X54Y106_SLICE_X82Y106_AMUX = CLBLL_L_X54Y106_SLICE_X82Y106_A_XOR;
  assign CLBLL_L_X54Y106_SLICE_X82Y106_BMUX = CLBLL_L_X54Y106_SLICE_X82Y106_B_XOR;
  assign CLBLL_L_X54Y106_SLICE_X82Y106_CMUX = CLBLL_L_X54Y106_SLICE_X82Y106_C_XOR;
  assign CLBLL_L_X54Y106_SLICE_X82Y106_DMUX = CLBLL_L_X54Y106_SLICE_X82Y106_D_XOR;
  assign CLBLL_L_X54Y106_SLICE_X83Y106_A = CLBLL_L_X54Y106_SLICE_X83Y106_AO6;
  assign CLBLL_L_X54Y106_SLICE_X83Y106_B = CLBLL_L_X54Y106_SLICE_X83Y106_BO6;
  assign CLBLL_L_X54Y106_SLICE_X83Y106_C = CLBLL_L_X54Y106_SLICE_X83Y106_CO6;
  assign CLBLL_L_X54Y106_SLICE_X83Y106_D = CLBLL_L_X54Y106_SLICE_X83Y106_DO6;
  assign CLBLL_L_X54Y106_SLICE_X83Y106_AMUX = CLBLL_L_X54Y106_SLICE_X83Y106_AO5;
  assign CLBLL_L_X54Y106_SLICE_X83Y106_BMUX = CLBLL_L_X54Y106_SLICE_X83Y106_BO6;
  assign CLBLL_L_X54Y106_SLICE_X83Y106_CMUX = CLBLL_L_X54Y106_SLICE_X83Y106_CO6;
  assign CLBLL_L_X54Y107_SLICE_X82Y107_A = CLBLL_L_X54Y107_SLICE_X82Y107_AO6;
  assign CLBLL_L_X54Y107_SLICE_X82Y107_B = CLBLL_L_X54Y107_SLICE_X82Y107_BO6;
  assign CLBLL_L_X54Y107_SLICE_X82Y107_C = CLBLL_L_X54Y107_SLICE_X82Y107_CO6;
  assign CLBLL_L_X54Y107_SLICE_X82Y107_D = CLBLL_L_X54Y107_SLICE_X82Y107_DO6;
  assign CLBLL_L_X54Y107_SLICE_X82Y107_AMUX = CLBLL_L_X54Y107_SLICE_X82Y107_A_XOR;
  assign CLBLL_L_X54Y107_SLICE_X82Y107_BMUX = CLBLL_L_X54Y107_SLICE_X82Y107_B_XOR;
  assign CLBLL_L_X54Y107_SLICE_X82Y107_CMUX = CLBLL_L_X54Y107_SLICE_X82Y107_C_XOR;
  assign CLBLL_L_X54Y107_SLICE_X82Y107_DMUX = CLBLL_L_X54Y107_SLICE_X82Y107_D_XOR;
  assign CLBLL_L_X54Y107_SLICE_X83Y107_A = CLBLL_L_X54Y107_SLICE_X83Y107_AO6;
  assign CLBLL_L_X54Y107_SLICE_X83Y107_B = CLBLL_L_X54Y107_SLICE_X83Y107_BO6;
  assign CLBLL_L_X54Y107_SLICE_X83Y107_C = CLBLL_L_X54Y107_SLICE_X83Y107_CO6;
  assign CLBLL_L_X54Y107_SLICE_X83Y107_D = CLBLL_L_X54Y107_SLICE_X83Y107_DO6;
  assign CLBLL_L_X54Y107_SLICE_X83Y107_AMUX = CLBLL_L_X54Y107_SLICE_X83Y107_AO5;
  assign CLBLL_L_X54Y107_SLICE_X83Y107_BMUX = CLBLL_L_X54Y107_SLICE_X83Y107_BO6;
  assign CLBLL_L_X54Y107_SLICE_X83Y107_DMUX = CLBLL_L_X54Y107_SLICE_X83Y107_DO6;
  assign CLBLL_L_X54Y108_SLICE_X82Y108_A = CLBLL_L_X54Y108_SLICE_X82Y108_AO6;
  assign CLBLL_L_X54Y108_SLICE_X82Y108_B = CLBLL_L_X54Y108_SLICE_X82Y108_BO6;
  assign CLBLL_L_X54Y108_SLICE_X82Y108_C = CLBLL_L_X54Y108_SLICE_X82Y108_CO6;
  assign CLBLL_L_X54Y108_SLICE_X82Y108_D = CLBLL_L_X54Y108_SLICE_X82Y108_DO6;
  assign CLBLL_L_X54Y108_SLICE_X82Y108_AMUX = CLBLL_L_X54Y108_SLICE_X82Y108_A_XOR;
  assign CLBLL_L_X54Y108_SLICE_X83Y108_A = CLBLL_L_X54Y108_SLICE_X83Y108_AO6;
  assign CLBLL_L_X54Y108_SLICE_X83Y108_B = CLBLL_L_X54Y108_SLICE_X83Y108_BO6;
  assign CLBLL_L_X54Y108_SLICE_X83Y108_C = CLBLL_L_X54Y108_SLICE_X83Y108_CO6;
  assign CLBLL_L_X54Y108_SLICE_X83Y108_D = CLBLL_L_X54Y108_SLICE_X83Y108_DO6;
  assign CLBLL_L_X54Y108_SLICE_X83Y108_AMUX = CLBLL_L_X54Y108_SLICE_X83Y108_AO5;
  assign CLBLL_L_X54Y109_SLICE_X82Y109_A = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLL_L_X54Y109_SLICE_X82Y109_B = CLBLL_L_X54Y109_SLICE_X82Y109_BO6;
  assign CLBLL_L_X54Y109_SLICE_X82Y109_C = CLBLL_L_X54Y109_SLICE_X82Y109_CO6;
  assign CLBLL_L_X54Y109_SLICE_X82Y109_D = CLBLL_L_X54Y109_SLICE_X82Y109_DO6;
  assign CLBLL_L_X54Y109_SLICE_X83Y109_A = CLBLL_L_X54Y109_SLICE_X83Y109_AO6;
  assign CLBLL_L_X54Y109_SLICE_X83Y109_B = CLBLL_L_X54Y109_SLICE_X83Y109_BO6;
  assign CLBLL_L_X54Y109_SLICE_X83Y109_C = CLBLL_L_X54Y109_SLICE_X83Y109_CO6;
  assign CLBLL_L_X54Y109_SLICE_X83Y109_D = CLBLL_L_X54Y109_SLICE_X83Y109_DO6;
  assign CLBLL_R_X57Y97_SLICE_X86Y97_A = CLBLL_R_X57Y97_SLICE_X86Y97_AO6;
  assign CLBLL_R_X57Y97_SLICE_X86Y97_B = CLBLL_R_X57Y97_SLICE_X86Y97_BO6;
  assign CLBLL_R_X57Y97_SLICE_X86Y97_C = CLBLL_R_X57Y97_SLICE_X86Y97_CO6;
  assign CLBLL_R_X57Y97_SLICE_X86Y97_D = CLBLL_R_X57Y97_SLICE_X86Y97_DO6;
  assign CLBLL_R_X57Y97_SLICE_X86Y97_BMUX = CLBLL_R_X57Y97_SLICE_X86Y97_BO6;
  assign CLBLL_R_X57Y97_SLICE_X87Y97_A = CLBLL_R_X57Y97_SLICE_X87Y97_AO6;
  assign CLBLL_R_X57Y97_SLICE_X87Y97_B = CLBLL_R_X57Y97_SLICE_X87Y97_BO6;
  assign CLBLL_R_X57Y97_SLICE_X87Y97_C = CLBLL_R_X57Y97_SLICE_X87Y97_CO6;
  assign CLBLL_R_X57Y97_SLICE_X87Y97_D = CLBLL_R_X57Y97_SLICE_X87Y97_DO6;
  assign CLBLL_R_X57Y98_SLICE_X86Y98_A = CLBLL_R_X57Y98_SLICE_X86Y98_AO6;
  assign CLBLL_R_X57Y98_SLICE_X86Y98_B = CLBLL_R_X57Y98_SLICE_X86Y98_BO6;
  assign CLBLL_R_X57Y98_SLICE_X86Y98_C = CLBLL_R_X57Y98_SLICE_X86Y98_CO6;
  assign CLBLL_R_X57Y98_SLICE_X86Y98_D = CLBLL_R_X57Y98_SLICE_X86Y98_DO6;
  assign CLBLL_R_X57Y98_SLICE_X87Y98_A = CLBLL_R_X57Y98_SLICE_X87Y98_AO6;
  assign CLBLL_R_X57Y98_SLICE_X87Y98_B = CLBLL_R_X57Y98_SLICE_X87Y98_BO6;
  assign CLBLL_R_X57Y98_SLICE_X87Y98_C = CLBLL_R_X57Y98_SLICE_X87Y98_CO6;
  assign CLBLL_R_X57Y98_SLICE_X87Y98_D = CLBLL_R_X57Y98_SLICE_X87Y98_DO6;
  assign CLBLL_R_X57Y99_SLICE_X86Y99_A = CLBLL_R_X57Y99_SLICE_X86Y99_AO6;
  assign CLBLL_R_X57Y99_SLICE_X86Y99_B = CLBLL_R_X57Y99_SLICE_X86Y99_BO6;
  assign CLBLL_R_X57Y99_SLICE_X86Y99_C = CLBLL_R_X57Y99_SLICE_X86Y99_CO6;
  assign CLBLL_R_X57Y99_SLICE_X86Y99_D = CLBLL_R_X57Y99_SLICE_X86Y99_DO6;
  assign CLBLL_R_X57Y99_SLICE_X87Y99_A = CLBLL_R_X57Y99_SLICE_X87Y99_AO6;
  assign CLBLL_R_X57Y99_SLICE_X87Y99_B = CLBLL_R_X57Y99_SLICE_X87Y99_BO6;
  assign CLBLL_R_X57Y99_SLICE_X87Y99_C = CLBLL_R_X57Y99_SLICE_X87Y99_CO6;
  assign CLBLL_R_X57Y99_SLICE_X87Y99_D = CLBLL_R_X57Y99_SLICE_X87Y99_DO6;
  assign CLBLL_R_X57Y100_SLICE_X86Y100_A = CLBLL_R_X57Y100_SLICE_X86Y100_AO6;
  assign CLBLL_R_X57Y100_SLICE_X86Y100_B = CLBLL_R_X57Y100_SLICE_X86Y100_BO6;
  assign CLBLL_R_X57Y100_SLICE_X86Y100_C = CLBLL_R_X57Y100_SLICE_X86Y100_CO6;
  assign CLBLL_R_X57Y100_SLICE_X86Y100_D = CLBLL_R_X57Y100_SLICE_X86Y100_DO6;
  assign CLBLL_R_X57Y100_SLICE_X86Y100_AMUX = CLBLL_R_X57Y100_SLICE_X86Y100_AO6;
  assign CLBLL_R_X57Y100_SLICE_X87Y100_A = CLBLL_R_X57Y100_SLICE_X87Y100_AO6;
  assign CLBLL_R_X57Y100_SLICE_X87Y100_B = CLBLL_R_X57Y100_SLICE_X87Y100_BO6;
  assign CLBLL_R_X57Y100_SLICE_X87Y100_C = CLBLL_R_X57Y100_SLICE_X87Y100_CO6;
  assign CLBLL_R_X57Y100_SLICE_X87Y100_D = CLBLL_R_X57Y100_SLICE_X87Y100_DO6;
  assign CLBLL_R_X57Y101_SLICE_X86Y101_A = CLBLL_R_X57Y101_SLICE_X86Y101_AO6;
  assign CLBLL_R_X57Y101_SLICE_X86Y101_B = CLBLL_R_X57Y101_SLICE_X86Y101_BO6;
  assign CLBLL_R_X57Y101_SLICE_X86Y101_C = CLBLL_R_X57Y101_SLICE_X86Y101_CO6;
  assign CLBLL_R_X57Y101_SLICE_X86Y101_D = CLBLL_R_X57Y101_SLICE_X86Y101_DO6;
  assign CLBLL_R_X57Y101_SLICE_X86Y101_AMUX = CLBLL_R_X57Y101_SLICE_X86Y101_AO5;
  assign CLBLL_R_X57Y101_SLICE_X87Y101_A = CLBLL_R_X57Y101_SLICE_X87Y101_AO6;
  assign CLBLL_R_X57Y101_SLICE_X87Y101_B = CLBLL_R_X57Y101_SLICE_X87Y101_BO6;
  assign CLBLL_R_X57Y101_SLICE_X87Y101_C = CLBLL_R_X57Y101_SLICE_X87Y101_CO6;
  assign CLBLL_R_X57Y101_SLICE_X87Y101_D = CLBLL_R_X57Y101_SLICE_X87Y101_DO6;
  assign CLBLL_R_X57Y101_SLICE_X87Y101_BMUX = CLBLL_R_X57Y101_SLICE_X87Y101_BO5;
  assign CLBLL_R_X57Y102_SLICE_X86Y102_A = CLBLL_R_X57Y102_SLICE_X86Y102_AO6;
  assign CLBLL_R_X57Y102_SLICE_X86Y102_B = CLBLL_R_X57Y102_SLICE_X86Y102_BO6;
  assign CLBLL_R_X57Y102_SLICE_X86Y102_C = CLBLL_R_X57Y102_SLICE_X86Y102_CO6;
  assign CLBLL_R_X57Y102_SLICE_X86Y102_D = CLBLL_R_X57Y102_SLICE_X86Y102_DO6;
  assign CLBLL_R_X57Y102_SLICE_X86Y102_AMUX = CLBLL_R_X57Y102_SLICE_X86Y102_AO5;
  assign CLBLL_R_X57Y102_SLICE_X86Y102_CMUX = CLBLL_R_X57Y102_SLICE_X86Y102_CO6;
  assign CLBLL_R_X57Y102_SLICE_X87Y102_A = CLBLL_R_X57Y102_SLICE_X87Y102_AO6;
  assign CLBLL_R_X57Y102_SLICE_X87Y102_B = CLBLL_R_X57Y102_SLICE_X87Y102_BO6;
  assign CLBLL_R_X57Y102_SLICE_X87Y102_C = CLBLL_R_X57Y102_SLICE_X87Y102_CO6;
  assign CLBLL_R_X57Y102_SLICE_X87Y102_D = CLBLL_R_X57Y102_SLICE_X87Y102_DO6;
  assign CLBLL_R_X57Y103_SLICE_X86Y103_A = CLBLL_R_X57Y103_SLICE_X86Y103_AO6;
  assign CLBLL_R_X57Y103_SLICE_X86Y103_B = CLBLL_R_X57Y103_SLICE_X86Y103_BO6;
  assign CLBLL_R_X57Y103_SLICE_X86Y103_C = CLBLL_R_X57Y103_SLICE_X86Y103_CO6;
  assign CLBLL_R_X57Y103_SLICE_X86Y103_D = CLBLL_R_X57Y103_SLICE_X86Y103_DO6;
  assign CLBLL_R_X57Y103_SLICE_X86Y103_AMUX = CLBLL_R_X57Y103_SLICE_X86Y103_A5Q;
  assign CLBLL_R_X57Y103_SLICE_X87Y103_A = CLBLL_R_X57Y103_SLICE_X87Y103_AO6;
  assign CLBLL_R_X57Y103_SLICE_X87Y103_B = CLBLL_R_X57Y103_SLICE_X87Y103_BO6;
  assign CLBLL_R_X57Y103_SLICE_X87Y103_C = CLBLL_R_X57Y103_SLICE_X87Y103_CO6;
  assign CLBLL_R_X57Y103_SLICE_X87Y103_D = CLBLL_R_X57Y103_SLICE_X87Y103_DO6;
  assign CLBLL_R_X57Y104_SLICE_X86Y104_A = CLBLL_R_X57Y104_SLICE_X86Y104_AO6;
  assign CLBLL_R_X57Y104_SLICE_X86Y104_B = CLBLL_R_X57Y104_SLICE_X86Y104_BO6;
  assign CLBLL_R_X57Y104_SLICE_X86Y104_C = CLBLL_R_X57Y104_SLICE_X86Y104_CO6;
  assign CLBLL_R_X57Y104_SLICE_X86Y104_D = CLBLL_R_X57Y104_SLICE_X86Y104_DO6;
  assign CLBLL_R_X57Y104_SLICE_X87Y104_A = CLBLL_R_X57Y104_SLICE_X87Y104_AO6;
  assign CLBLL_R_X57Y104_SLICE_X87Y104_B = CLBLL_R_X57Y104_SLICE_X87Y104_BO6;
  assign CLBLL_R_X57Y104_SLICE_X87Y104_C = CLBLL_R_X57Y104_SLICE_X87Y104_CO6;
  assign CLBLL_R_X57Y104_SLICE_X87Y104_D = CLBLL_R_X57Y104_SLICE_X87Y104_DO6;
  assign CLBLL_R_X57Y105_SLICE_X86Y105_A = CLBLL_R_X57Y105_SLICE_X86Y105_AO6;
  assign CLBLL_R_X57Y105_SLICE_X86Y105_B = CLBLL_R_X57Y105_SLICE_X86Y105_BO6;
  assign CLBLL_R_X57Y105_SLICE_X86Y105_C = CLBLL_R_X57Y105_SLICE_X86Y105_CO6;
  assign CLBLL_R_X57Y105_SLICE_X86Y105_D = CLBLL_R_X57Y105_SLICE_X86Y105_DO6;
  assign CLBLL_R_X57Y105_SLICE_X87Y105_A = CLBLL_R_X57Y105_SLICE_X87Y105_AO6;
  assign CLBLL_R_X57Y105_SLICE_X87Y105_B = CLBLL_R_X57Y105_SLICE_X87Y105_BO6;
  assign CLBLL_R_X57Y105_SLICE_X87Y105_C = CLBLL_R_X57Y105_SLICE_X87Y105_CO6;
  assign CLBLL_R_X57Y105_SLICE_X87Y105_D = CLBLL_R_X57Y105_SLICE_X87Y105_DO6;
  assign CLBLL_R_X57Y105_SLICE_X87Y105_AMUX = CLBLL_R_X57Y105_SLICE_X87Y105_A_XOR;
  assign CLBLL_R_X57Y105_SLICE_X87Y105_BMUX = CLBLL_R_X57Y105_SLICE_X87Y105_B_XOR;
  assign CLBLL_R_X57Y105_SLICE_X87Y105_CMUX = CLBLL_R_X57Y105_SLICE_X87Y105_C_XOR;
  assign CLBLL_R_X57Y105_SLICE_X87Y105_DMUX = CLBLL_R_X57Y105_SLICE_X87Y105_D_XOR;
  assign CLBLL_R_X57Y106_SLICE_X86Y106_A = CLBLL_R_X57Y106_SLICE_X86Y106_AO6;
  assign CLBLL_R_X57Y106_SLICE_X86Y106_B = CLBLL_R_X57Y106_SLICE_X86Y106_BO6;
  assign CLBLL_R_X57Y106_SLICE_X86Y106_C = CLBLL_R_X57Y106_SLICE_X86Y106_CO6;
  assign CLBLL_R_X57Y106_SLICE_X86Y106_D = CLBLL_R_X57Y106_SLICE_X86Y106_DO6;
  assign CLBLL_R_X57Y106_SLICE_X86Y106_AMUX = CLBLL_R_X57Y106_SLICE_X86Y106_A_XOR;
  assign CLBLL_R_X57Y106_SLICE_X86Y106_BMUX = CLBLL_R_X57Y106_SLICE_X86Y106_B_XOR;
  assign CLBLL_R_X57Y106_SLICE_X86Y106_CMUX = CLBLL_R_X57Y106_SLICE_X86Y106_C_XOR;
  assign CLBLL_R_X57Y106_SLICE_X86Y106_DMUX = CLBLL_R_X57Y106_SLICE_X86Y106_D_XOR;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_A = CLBLL_R_X57Y106_SLICE_X87Y106_AO6;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_B = CLBLL_R_X57Y106_SLICE_X87Y106_BO6;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_C = CLBLL_R_X57Y106_SLICE_X87Y106_CO6;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_D = CLBLL_R_X57Y106_SLICE_X87Y106_DO6;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_AMUX = CLBLL_R_X57Y106_SLICE_X87Y106_A_XOR;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_BMUX = CLBLL_R_X57Y106_SLICE_X87Y106_B_XOR;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_CMUX = CLBLL_R_X57Y106_SLICE_X87Y106_C_XOR;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_DMUX = CLBLL_R_X57Y106_SLICE_X87Y106_D_XOR;
  assign CLBLL_R_X57Y107_SLICE_X86Y107_A = CLBLL_R_X57Y107_SLICE_X86Y107_AO6;
  assign CLBLL_R_X57Y107_SLICE_X86Y107_B = CLBLL_R_X57Y107_SLICE_X86Y107_BO6;
  assign CLBLL_R_X57Y107_SLICE_X86Y107_C = CLBLL_R_X57Y107_SLICE_X86Y107_CO6;
  assign CLBLL_R_X57Y107_SLICE_X86Y107_D = CLBLL_R_X57Y107_SLICE_X86Y107_DO6;
  assign CLBLL_R_X57Y107_SLICE_X86Y107_AMUX = CLBLL_R_X57Y107_SLICE_X86Y107_A_XOR;
  assign CLBLL_R_X57Y107_SLICE_X86Y107_BMUX = CLBLL_R_X57Y107_SLICE_X86Y107_B_XOR;
  assign CLBLL_R_X57Y107_SLICE_X86Y107_CMUX = CLBLL_R_X57Y107_SLICE_X86Y107_C_XOR;
  assign CLBLL_R_X57Y107_SLICE_X86Y107_DMUX = CLBLL_R_X57Y107_SLICE_X86Y107_D_XOR;
  assign CLBLL_R_X57Y107_SLICE_X87Y107_A = CLBLL_R_X57Y107_SLICE_X87Y107_AO6;
  assign CLBLL_R_X57Y107_SLICE_X87Y107_B = CLBLL_R_X57Y107_SLICE_X87Y107_BO6;
  assign CLBLL_R_X57Y107_SLICE_X87Y107_C = CLBLL_R_X57Y107_SLICE_X87Y107_CO6;
  assign CLBLL_R_X57Y107_SLICE_X87Y107_D = CLBLL_R_X57Y107_SLICE_X87Y107_DO6;
  assign CLBLL_R_X57Y107_SLICE_X87Y107_AMUX = CLBLL_R_X57Y107_SLICE_X87Y107_A_XOR;
  assign CLBLL_R_X57Y107_SLICE_X87Y107_BMUX = CLBLL_R_X57Y107_SLICE_X87Y107_B_XOR;
  assign CLBLL_R_X57Y107_SLICE_X87Y107_CMUX = CLBLL_R_X57Y107_SLICE_X87Y107_C_XOR;
  assign CLBLL_R_X57Y108_SLICE_X86Y108_A = CLBLL_R_X57Y108_SLICE_X86Y108_AO6;
  assign CLBLL_R_X57Y108_SLICE_X86Y108_B = CLBLL_R_X57Y108_SLICE_X86Y108_BO6;
  assign CLBLL_R_X57Y108_SLICE_X86Y108_C = CLBLL_R_X57Y108_SLICE_X86Y108_CO6;
  assign CLBLL_R_X57Y108_SLICE_X86Y108_D = CLBLL_R_X57Y108_SLICE_X86Y108_DO6;
  assign CLBLL_R_X57Y108_SLICE_X86Y108_AMUX = CLBLL_R_X57Y108_SLICE_X86Y108_A_XOR;
  assign CLBLL_R_X57Y108_SLICE_X86Y108_BMUX = CLBLL_R_X57Y108_SLICE_X86Y108_B_XOR;
  assign CLBLL_R_X57Y108_SLICE_X86Y108_CMUX = CLBLL_R_X57Y108_SLICE_X86Y108_C_XOR;
  assign CLBLL_R_X57Y108_SLICE_X87Y108_A = CLBLL_R_X57Y108_SLICE_X87Y108_AO6;
  assign CLBLL_R_X57Y108_SLICE_X87Y108_B = CLBLL_R_X57Y108_SLICE_X87Y108_BO6;
  assign CLBLL_R_X57Y108_SLICE_X87Y108_C = CLBLL_R_X57Y108_SLICE_X87Y108_CO6;
  assign CLBLL_R_X57Y108_SLICE_X87Y108_D = CLBLL_R_X57Y108_SLICE_X87Y108_DO6;
  assign CLBLL_R_X57Y109_SLICE_X86Y109_A = CLBLL_R_X57Y109_SLICE_X86Y109_AO6;
  assign CLBLL_R_X57Y109_SLICE_X86Y109_B = CLBLL_R_X57Y109_SLICE_X86Y109_BO6;
  assign CLBLL_R_X57Y109_SLICE_X86Y109_C = CLBLL_R_X57Y109_SLICE_X86Y109_CO6;
  assign CLBLL_R_X57Y109_SLICE_X86Y109_D = CLBLL_R_X57Y109_SLICE_X86Y109_DO6;
  assign CLBLL_R_X57Y109_SLICE_X87Y109_A = CLBLL_R_X57Y109_SLICE_X87Y109_AO6;
  assign CLBLL_R_X57Y109_SLICE_X87Y109_B = CLBLL_R_X57Y109_SLICE_X87Y109_BO6;
  assign CLBLL_R_X57Y109_SLICE_X87Y109_C = CLBLL_R_X57Y109_SLICE_X87Y109_CO6;
  assign CLBLL_R_X57Y109_SLICE_X87Y109_D = CLBLL_R_X57Y109_SLICE_X87Y109_DO6;
  assign CLBLL_R_X57Y109_SLICE_X87Y109_AMUX = CLBLL_R_X57Y109_SLICE_X87Y109_A_XOR;
  assign CLBLL_R_X57Y109_SLICE_X87Y109_BMUX = CLBLL_R_X57Y109_SLICE_X87Y109_B_XOR;
  assign CLBLL_R_X57Y109_SLICE_X87Y109_CMUX = CLBLL_R_X57Y109_SLICE_X87Y109_C_XOR;
  assign CLBLL_R_X57Y109_SLICE_X87Y109_DMUX = CLBLL_R_X57Y109_SLICE_X87Y109_D_XOR;
  assign CLBLL_R_X57Y110_SLICE_X86Y110_A = CLBLL_R_X57Y110_SLICE_X86Y110_AO6;
  assign CLBLL_R_X57Y110_SLICE_X86Y110_B = CLBLL_R_X57Y110_SLICE_X86Y110_BO6;
  assign CLBLL_R_X57Y110_SLICE_X86Y110_C = CLBLL_R_X57Y110_SLICE_X86Y110_CO6;
  assign CLBLL_R_X57Y110_SLICE_X86Y110_D = CLBLL_R_X57Y110_SLICE_X86Y110_DO6;
  assign CLBLL_R_X57Y110_SLICE_X87Y110_A = CLBLL_R_X57Y110_SLICE_X87Y110_AO6;
  assign CLBLL_R_X57Y110_SLICE_X87Y110_B = CLBLL_R_X57Y110_SLICE_X87Y110_BO6;
  assign CLBLL_R_X57Y110_SLICE_X87Y110_C = CLBLL_R_X57Y110_SLICE_X87Y110_CO6;
  assign CLBLL_R_X57Y110_SLICE_X87Y110_D = CLBLL_R_X57Y110_SLICE_X87Y110_DO6;
  assign CLBLL_R_X57Y110_SLICE_X87Y110_AMUX = CLBLL_R_X57Y110_SLICE_X87Y110_A_XOR;
  assign CLBLL_R_X57Y110_SLICE_X87Y110_BMUX = CLBLL_R_X57Y110_SLICE_X87Y110_B_XOR;
  assign CLBLL_R_X57Y110_SLICE_X87Y110_CMUX = CLBLL_R_X57Y110_SLICE_X87Y110_C_XOR;
  assign CLBLL_R_X57Y110_SLICE_X87Y110_DMUX = CLBLL_R_X57Y110_SLICE_X87Y110_D_XOR;
  assign CLBLL_R_X57Y111_SLICE_X86Y111_A = CLBLL_R_X57Y111_SLICE_X86Y111_AO6;
  assign CLBLL_R_X57Y111_SLICE_X86Y111_B = CLBLL_R_X57Y111_SLICE_X86Y111_BO6;
  assign CLBLL_R_X57Y111_SLICE_X86Y111_C = CLBLL_R_X57Y111_SLICE_X86Y111_CO6;
  assign CLBLL_R_X57Y111_SLICE_X86Y111_D = CLBLL_R_X57Y111_SLICE_X86Y111_DO6;
  assign CLBLL_R_X57Y111_SLICE_X87Y111_A = CLBLL_R_X57Y111_SLICE_X87Y111_AO6;
  assign CLBLL_R_X57Y111_SLICE_X87Y111_B = CLBLL_R_X57Y111_SLICE_X87Y111_BO6;
  assign CLBLL_R_X57Y111_SLICE_X87Y111_C = CLBLL_R_X57Y111_SLICE_X87Y111_CO6;
  assign CLBLL_R_X57Y111_SLICE_X87Y111_D = CLBLL_R_X57Y111_SLICE_X87Y111_DO6;
  assign CLBLL_R_X57Y111_SLICE_X87Y111_AMUX = CLBLL_R_X57Y111_SLICE_X87Y111_A_XOR;
  assign CLBLL_R_X57Y111_SLICE_X87Y111_BMUX = CLBLL_R_X57Y111_SLICE_X87Y111_B_XOR;
  assign CLBLL_R_X57Y111_SLICE_X87Y111_CMUX = CLBLL_R_X57Y111_SLICE_X87Y111_C_XOR;
  assign CLBLL_R_X57Y111_SLICE_X87Y111_DMUX = CLBLL_R_X57Y111_SLICE_X87Y111_D_XOR;
  assign CLBLM_L_X32Y119_SLICE_X46Y119_A = CLBLM_L_X32Y119_SLICE_X46Y119_AO6;
  assign CLBLM_L_X32Y119_SLICE_X46Y119_B = CLBLM_L_X32Y119_SLICE_X46Y119_BO6;
  assign CLBLM_L_X32Y119_SLICE_X46Y119_C = CLBLM_L_X32Y119_SLICE_X46Y119_CO6;
  assign CLBLM_L_X32Y119_SLICE_X46Y119_D = CLBLM_L_X32Y119_SLICE_X46Y119_DO6;
  assign CLBLM_L_X32Y119_SLICE_X47Y119_A = CLBLM_L_X32Y119_SLICE_X47Y119_AO6;
  assign CLBLM_L_X32Y119_SLICE_X47Y119_B = CLBLM_L_X32Y119_SLICE_X47Y119_BO6;
  assign CLBLM_L_X32Y119_SLICE_X47Y119_C = CLBLM_L_X32Y119_SLICE_X47Y119_CO6;
  assign CLBLM_L_X32Y119_SLICE_X47Y119_D = CLBLM_L_X32Y119_SLICE_X47Y119_DO6;
  assign CLBLM_L_X50Y104_SLICE_X76Y104_A = CLBLM_L_X50Y104_SLICE_X76Y104_AO6;
  assign CLBLM_L_X50Y104_SLICE_X76Y104_B = CLBLM_L_X50Y104_SLICE_X76Y104_BO6;
  assign CLBLM_L_X50Y104_SLICE_X76Y104_C = CLBLM_L_X50Y104_SLICE_X76Y104_CO6;
  assign CLBLM_L_X50Y104_SLICE_X76Y104_D = CLBLM_L_X50Y104_SLICE_X76Y104_DO6;
  assign CLBLM_L_X50Y104_SLICE_X77Y104_A = CLBLM_L_X50Y104_SLICE_X77Y104_AO6;
  assign CLBLM_L_X50Y104_SLICE_X77Y104_B = CLBLM_L_X50Y104_SLICE_X77Y104_BO6;
  assign CLBLM_L_X50Y104_SLICE_X77Y104_C = CLBLM_L_X50Y104_SLICE_X77Y104_CO6;
  assign CLBLM_L_X50Y104_SLICE_X77Y104_D = CLBLM_L_X50Y104_SLICE_X77Y104_DO6;
  assign CLBLM_L_X50Y105_SLICE_X76Y105_A = CLBLM_L_X50Y105_SLICE_X76Y105_AO6;
  assign CLBLM_L_X50Y105_SLICE_X76Y105_B = CLBLM_L_X50Y105_SLICE_X76Y105_BO6;
  assign CLBLM_L_X50Y105_SLICE_X76Y105_C = CLBLM_L_X50Y105_SLICE_X76Y105_CO6;
  assign CLBLM_L_X50Y105_SLICE_X76Y105_D = CLBLM_L_X50Y105_SLICE_X76Y105_DO6;
  assign CLBLM_L_X50Y105_SLICE_X76Y105_BMUX = CLBLM_L_X50Y105_SLICE_X76Y105_BO5;
  assign CLBLM_L_X50Y105_SLICE_X76Y105_CMUX = CLBLM_L_X50Y105_SLICE_X76Y105_CO5;
  assign CLBLM_L_X50Y105_SLICE_X77Y105_A = CLBLM_L_X50Y105_SLICE_X77Y105_AO6;
  assign CLBLM_L_X50Y105_SLICE_X77Y105_B = CLBLM_L_X50Y105_SLICE_X77Y105_BO6;
  assign CLBLM_L_X50Y105_SLICE_X77Y105_C = CLBLM_L_X50Y105_SLICE_X77Y105_CO6;
  assign CLBLM_L_X50Y105_SLICE_X77Y105_D = CLBLM_L_X50Y105_SLICE_X77Y105_DO6;
  assign CLBLM_L_X50Y106_SLICE_X76Y106_A = CLBLM_L_X50Y106_SLICE_X76Y106_AO6;
  assign CLBLM_L_X50Y106_SLICE_X76Y106_B = CLBLM_L_X50Y106_SLICE_X76Y106_BO6;
  assign CLBLM_L_X50Y106_SLICE_X76Y106_C = CLBLM_L_X50Y106_SLICE_X76Y106_CO6;
  assign CLBLM_L_X50Y106_SLICE_X76Y106_D = CLBLM_L_X50Y106_SLICE_X76Y106_DO6;
  assign CLBLM_L_X50Y106_SLICE_X76Y106_BMUX = CLBLM_L_X50Y106_SLICE_X76Y106_BO5;
  assign CLBLM_L_X50Y106_SLICE_X77Y106_A = CLBLM_L_X50Y106_SLICE_X77Y106_AO6;
  assign CLBLM_L_X50Y106_SLICE_X77Y106_B = CLBLM_L_X50Y106_SLICE_X77Y106_BO6;
  assign CLBLM_L_X50Y106_SLICE_X77Y106_C = CLBLM_L_X50Y106_SLICE_X77Y106_CO6;
  assign CLBLM_L_X50Y106_SLICE_X77Y106_D = CLBLM_L_X50Y106_SLICE_X77Y106_DO6;
  assign CLBLM_L_X50Y106_SLICE_X77Y106_AMUX = CLBLM_L_X50Y106_SLICE_X77Y106_AO5;
  assign CLBLM_L_X50Y106_SLICE_X77Y106_BMUX = CLBLM_L_X50Y106_SLICE_X77Y106_BO5;
  assign CLBLM_L_X50Y107_SLICE_X76Y107_A = CLBLM_L_X50Y107_SLICE_X76Y107_AO6;
  assign CLBLM_L_X50Y107_SLICE_X76Y107_B = CLBLM_L_X50Y107_SLICE_X76Y107_BO6;
  assign CLBLM_L_X50Y107_SLICE_X76Y107_C = CLBLM_L_X50Y107_SLICE_X76Y107_CO6;
  assign CLBLM_L_X50Y107_SLICE_X76Y107_D = CLBLM_L_X50Y107_SLICE_X76Y107_DO6;
  assign CLBLM_L_X50Y107_SLICE_X76Y107_AMUX = CLBLM_L_X50Y107_SLICE_X76Y107_AO5;
  assign CLBLM_L_X50Y107_SLICE_X77Y107_A = CLBLM_L_X50Y107_SLICE_X77Y107_AO6;
  assign CLBLM_L_X50Y107_SLICE_X77Y107_B = CLBLM_L_X50Y107_SLICE_X77Y107_BO6;
  assign CLBLM_L_X50Y107_SLICE_X77Y107_C = CLBLM_L_X50Y107_SLICE_X77Y107_CO6;
  assign CLBLM_L_X50Y107_SLICE_X77Y107_D = CLBLM_L_X50Y107_SLICE_X77Y107_DO6;
  assign CLBLM_L_X50Y108_SLICE_X76Y108_A = CLBLM_L_X50Y108_SLICE_X76Y108_AO6;
  assign CLBLM_L_X50Y108_SLICE_X76Y108_B = CLBLM_L_X50Y108_SLICE_X76Y108_BO6;
  assign CLBLM_L_X50Y108_SLICE_X76Y108_C = CLBLM_L_X50Y108_SLICE_X76Y108_CO6;
  assign CLBLM_L_X50Y108_SLICE_X76Y108_D = CLBLM_L_X50Y108_SLICE_X76Y108_DO6;
  assign CLBLM_L_X50Y108_SLICE_X76Y108_AMUX = CLBLM_L_X50Y108_SLICE_X76Y108_A_XOR;
  assign CLBLM_L_X50Y108_SLICE_X76Y108_BMUX = CLBLM_L_X50Y108_SLICE_X76Y108_B_XOR;
  assign CLBLM_L_X50Y108_SLICE_X76Y108_CMUX = CLBLM_L_X50Y108_SLICE_X76Y108_C_XOR;
  assign CLBLM_L_X50Y108_SLICE_X76Y108_DMUX = CLBLM_L_X50Y108_SLICE_X76Y108_D_XOR;
  assign CLBLM_L_X50Y108_SLICE_X77Y108_A = CLBLM_L_X50Y108_SLICE_X77Y108_AO6;
  assign CLBLM_L_X50Y108_SLICE_X77Y108_B = CLBLM_L_X50Y108_SLICE_X77Y108_BO6;
  assign CLBLM_L_X50Y108_SLICE_X77Y108_C = CLBLM_L_X50Y108_SLICE_X77Y108_CO6;
  assign CLBLM_L_X50Y108_SLICE_X77Y108_D = CLBLM_L_X50Y108_SLICE_X77Y108_DO6;
  assign CLBLM_L_X50Y108_SLICE_X77Y108_AMUX = CLBLM_L_X50Y108_SLICE_X77Y108_A_XOR;
  assign CLBLM_L_X50Y108_SLICE_X77Y108_BMUX = CLBLM_L_X50Y108_SLICE_X77Y108_B_XOR;
  assign CLBLM_L_X50Y108_SLICE_X77Y108_CMUX = CLBLM_L_X50Y108_SLICE_X77Y108_C_XOR;
  assign CLBLM_L_X50Y108_SLICE_X77Y108_DMUX = CLBLM_L_X50Y108_SLICE_X77Y108_D_XOR;
  assign CLBLM_L_X50Y109_SLICE_X76Y109_A = CLBLM_L_X50Y109_SLICE_X76Y109_AO6;
  assign CLBLM_L_X50Y109_SLICE_X76Y109_B = CLBLM_L_X50Y109_SLICE_X76Y109_BO6;
  assign CLBLM_L_X50Y109_SLICE_X76Y109_C = CLBLM_L_X50Y109_SLICE_X76Y109_CO6;
  assign CLBLM_L_X50Y109_SLICE_X76Y109_D = CLBLM_L_X50Y109_SLICE_X76Y109_DO6;
  assign CLBLM_L_X50Y109_SLICE_X76Y109_AMUX = CLBLM_L_X50Y109_SLICE_X76Y109_A_XOR;
  assign CLBLM_L_X50Y109_SLICE_X76Y109_BMUX = CLBLM_L_X50Y109_SLICE_X76Y109_B_XOR;
  assign CLBLM_L_X50Y109_SLICE_X76Y109_CMUX = CLBLM_L_X50Y109_SLICE_X76Y109_C_XOR;
  assign CLBLM_L_X50Y109_SLICE_X76Y109_DMUX = CLBLM_L_X50Y109_SLICE_X76Y109_D_XOR;
  assign CLBLM_L_X50Y109_SLICE_X77Y109_A = CLBLM_L_X50Y109_SLICE_X77Y109_AO6;
  assign CLBLM_L_X50Y109_SLICE_X77Y109_B = CLBLM_L_X50Y109_SLICE_X77Y109_BO6;
  assign CLBLM_L_X50Y109_SLICE_X77Y109_C = CLBLM_L_X50Y109_SLICE_X77Y109_CO6;
  assign CLBLM_L_X50Y109_SLICE_X77Y109_D = CLBLM_L_X50Y109_SLICE_X77Y109_DO6;
  assign CLBLM_L_X50Y109_SLICE_X77Y109_AMUX = CLBLM_L_X50Y109_SLICE_X77Y109_A_XOR;
  assign CLBLM_L_X50Y109_SLICE_X77Y109_BMUX = CLBLM_L_X50Y109_SLICE_X77Y109_B_XOR;
  assign CLBLM_L_X50Y109_SLICE_X77Y109_CMUX = CLBLM_L_X50Y109_SLICE_X77Y109_C_XOR;
  assign CLBLM_L_X50Y109_SLICE_X77Y109_DMUX = CLBLM_L_X50Y109_SLICE_X77Y109_D_XOR;
  assign CLBLM_L_X50Y110_SLICE_X76Y110_A = CLBLM_L_X50Y110_SLICE_X76Y110_AO6;
  assign CLBLM_L_X50Y110_SLICE_X76Y110_B = CLBLM_L_X50Y110_SLICE_X76Y110_BO6;
  assign CLBLM_L_X50Y110_SLICE_X76Y110_C = CLBLM_L_X50Y110_SLICE_X76Y110_CO6;
  assign CLBLM_L_X50Y110_SLICE_X76Y110_D = CLBLM_L_X50Y110_SLICE_X76Y110_DO6;
  assign CLBLM_L_X50Y110_SLICE_X76Y110_AMUX = CLBLM_L_X50Y110_SLICE_X76Y110_A_CY;
  assign CLBLM_L_X50Y110_SLICE_X77Y110_A = CLBLM_L_X50Y110_SLICE_X77Y110_AO6;
  assign CLBLM_L_X50Y110_SLICE_X77Y110_B = CLBLM_L_X50Y110_SLICE_X77Y110_BO6;
  assign CLBLM_L_X50Y110_SLICE_X77Y110_C = CLBLM_L_X50Y110_SLICE_X77Y110_CO6;
  assign CLBLM_L_X50Y110_SLICE_X77Y110_D = CLBLM_L_X50Y110_SLICE_X77Y110_DO6;
  assign CLBLM_L_X50Y110_SLICE_X77Y110_AMUX = CLBLM_L_X50Y110_SLICE_X77Y110_A_XOR;
  assign CLBLM_L_X50Y111_SLICE_X76Y111_A = CLBLM_L_X50Y111_SLICE_X76Y111_AO6;
  assign CLBLM_L_X50Y111_SLICE_X76Y111_B = CLBLM_L_X50Y111_SLICE_X76Y111_BO6;
  assign CLBLM_L_X50Y111_SLICE_X76Y111_C = CLBLM_L_X50Y111_SLICE_X76Y111_CO6;
  assign CLBLM_L_X50Y111_SLICE_X76Y111_D = CLBLM_L_X50Y111_SLICE_X76Y111_DO6;
  assign CLBLM_L_X50Y111_SLICE_X76Y111_CMUX = CLBLM_L_X50Y111_SLICE_X76Y111_CO6;
  assign CLBLM_L_X50Y111_SLICE_X77Y111_A = CLBLM_L_X50Y111_SLICE_X77Y111_AO6;
  assign CLBLM_L_X50Y111_SLICE_X77Y111_B = CLBLM_L_X50Y111_SLICE_X77Y111_BO6;
  assign CLBLM_L_X50Y111_SLICE_X77Y111_C = CLBLM_L_X50Y111_SLICE_X77Y111_CO6;
  assign CLBLM_L_X50Y111_SLICE_X77Y111_D = CLBLM_L_X50Y111_SLICE_X77Y111_DO6;
  assign CLBLM_L_X56Y97_SLICE_X84Y97_A = CLBLM_L_X56Y97_SLICE_X84Y97_AO6;
  assign CLBLM_L_X56Y97_SLICE_X84Y97_B = CLBLM_L_X56Y97_SLICE_X84Y97_BO6;
  assign CLBLM_L_X56Y97_SLICE_X84Y97_C = CLBLM_L_X56Y97_SLICE_X84Y97_CO6;
  assign CLBLM_L_X56Y97_SLICE_X84Y97_D = CLBLM_L_X56Y97_SLICE_X84Y97_DO6;
  assign CLBLM_L_X56Y97_SLICE_X84Y97_AMUX = CLBLM_L_X56Y97_SLICE_X84Y97_AO5;
  assign CLBLM_L_X56Y97_SLICE_X84Y97_CMUX = CLBLM_L_X56Y97_SLICE_X84Y97_CO5;
  assign CLBLM_L_X56Y97_SLICE_X85Y97_A = CLBLM_L_X56Y97_SLICE_X85Y97_AO6;
  assign CLBLM_L_X56Y97_SLICE_X85Y97_B = CLBLM_L_X56Y97_SLICE_X85Y97_BO6;
  assign CLBLM_L_X56Y97_SLICE_X85Y97_C = CLBLM_L_X56Y97_SLICE_X85Y97_CO6;
  assign CLBLM_L_X56Y97_SLICE_X85Y97_D = CLBLM_L_X56Y97_SLICE_X85Y97_DO6;
  assign CLBLM_L_X56Y97_SLICE_X85Y97_BMUX = CLBLM_L_X56Y97_SLICE_X85Y97_BO5;
  assign CLBLM_L_X56Y98_SLICE_X84Y98_A = CLBLM_L_X56Y98_SLICE_X84Y98_AO6;
  assign CLBLM_L_X56Y98_SLICE_X84Y98_B = CLBLM_L_X56Y98_SLICE_X84Y98_BO6;
  assign CLBLM_L_X56Y98_SLICE_X84Y98_C = CLBLM_L_X56Y98_SLICE_X84Y98_CO6;
  assign CLBLM_L_X56Y98_SLICE_X84Y98_D = CLBLM_L_X56Y98_SLICE_X84Y98_DO6;
  assign CLBLM_L_X56Y98_SLICE_X84Y98_AMUX = CLBLM_L_X56Y98_SLICE_X84Y98_AO5;
  assign CLBLM_L_X56Y98_SLICE_X84Y98_BMUX = CLBLM_L_X56Y98_SLICE_X84Y98_BO6;
  assign CLBLM_L_X56Y98_SLICE_X84Y98_CMUX = CLBLM_L_X56Y98_SLICE_X84Y98_CO6;
  assign CLBLM_L_X56Y98_SLICE_X84Y98_DMUX = CLBLM_L_X56Y98_SLICE_X84Y98_DO5;
  assign CLBLM_L_X56Y98_SLICE_X85Y98_A = CLBLM_L_X56Y98_SLICE_X85Y98_AO6;
  assign CLBLM_L_X56Y98_SLICE_X85Y98_B = CLBLM_L_X56Y98_SLICE_X85Y98_BO6;
  assign CLBLM_L_X56Y98_SLICE_X85Y98_C = CLBLM_L_X56Y98_SLICE_X85Y98_CO6;
  assign CLBLM_L_X56Y98_SLICE_X85Y98_D = CLBLM_L_X56Y98_SLICE_X85Y98_DO6;
  assign CLBLM_L_X56Y98_SLICE_X85Y98_AMUX = CLBLM_L_X56Y98_SLICE_X85Y98_A5Q;
  assign CLBLM_L_X56Y98_SLICE_X85Y98_BMUX = CLBLM_L_X56Y98_SLICE_X85Y98_BO5;
  assign CLBLM_L_X56Y99_SLICE_X84Y99_A = CLBLM_L_X56Y99_SLICE_X84Y99_AO6;
  assign CLBLM_L_X56Y99_SLICE_X84Y99_B = CLBLM_L_X56Y99_SLICE_X84Y99_BO6;
  assign CLBLM_L_X56Y99_SLICE_X84Y99_C = CLBLM_L_X56Y99_SLICE_X84Y99_CO6;
  assign CLBLM_L_X56Y99_SLICE_X84Y99_D = CLBLM_L_X56Y99_SLICE_X84Y99_DO6;
  assign CLBLM_L_X56Y99_SLICE_X85Y99_A = CLBLM_L_X56Y99_SLICE_X85Y99_AO6;
  assign CLBLM_L_X56Y99_SLICE_X85Y99_B = CLBLM_L_X56Y99_SLICE_X85Y99_BO6;
  assign CLBLM_L_X56Y99_SLICE_X85Y99_C = CLBLM_L_X56Y99_SLICE_X85Y99_CO6;
  assign CLBLM_L_X56Y99_SLICE_X85Y99_D = CLBLM_L_X56Y99_SLICE_X85Y99_DO6;
  assign CLBLM_L_X56Y99_SLICE_X85Y99_AMUX = CLBLM_L_X56Y99_SLICE_X85Y99_A5Q;
  assign CLBLM_L_X56Y100_SLICE_X84Y100_A = CLBLM_L_X56Y100_SLICE_X84Y100_AO6;
  assign CLBLM_L_X56Y100_SLICE_X84Y100_B = CLBLM_L_X56Y100_SLICE_X84Y100_BO6;
  assign CLBLM_L_X56Y100_SLICE_X84Y100_C = CLBLM_L_X56Y100_SLICE_X84Y100_CO6;
  assign CLBLM_L_X56Y100_SLICE_X84Y100_D = CLBLM_L_X56Y100_SLICE_X84Y100_DO6;
  assign CLBLM_L_X56Y100_SLICE_X85Y100_A = CLBLM_L_X56Y100_SLICE_X85Y100_AO6;
  assign CLBLM_L_X56Y100_SLICE_X85Y100_B = CLBLM_L_X56Y100_SLICE_X85Y100_BO6;
  assign CLBLM_L_X56Y100_SLICE_X85Y100_C = CLBLM_L_X56Y100_SLICE_X85Y100_CO6;
  assign CLBLM_L_X56Y100_SLICE_X85Y100_D = CLBLM_L_X56Y100_SLICE_X85Y100_DO6;
  assign CLBLM_L_X56Y100_SLICE_X85Y100_AMUX = CLBLM_L_X56Y100_SLICE_X85Y100_AO5;
  assign CLBLM_L_X56Y100_SLICE_X85Y100_BMUX = CLBLM_L_X56Y100_SLICE_X85Y100_BO5;
  assign CLBLM_L_X56Y101_SLICE_X84Y101_A = CLBLM_L_X56Y101_SLICE_X84Y101_AO6;
  assign CLBLM_L_X56Y101_SLICE_X84Y101_B = CLBLM_L_X56Y101_SLICE_X84Y101_BO6;
  assign CLBLM_L_X56Y101_SLICE_X84Y101_C = CLBLM_L_X56Y101_SLICE_X84Y101_CO6;
  assign CLBLM_L_X56Y101_SLICE_X84Y101_D = CLBLM_L_X56Y101_SLICE_X84Y101_DO6;
  assign CLBLM_L_X56Y101_SLICE_X85Y101_A = CLBLM_L_X56Y101_SLICE_X85Y101_AO6;
  assign CLBLM_L_X56Y101_SLICE_X85Y101_B = CLBLM_L_X56Y101_SLICE_X85Y101_BO6;
  assign CLBLM_L_X56Y101_SLICE_X85Y101_C = CLBLM_L_X56Y101_SLICE_X85Y101_CO6;
  assign CLBLM_L_X56Y101_SLICE_X85Y101_D = CLBLM_L_X56Y101_SLICE_X85Y101_DO6;
  assign CLBLM_L_X56Y102_SLICE_X84Y102_A = CLBLM_L_X56Y102_SLICE_X84Y102_AO6;
  assign CLBLM_L_X56Y102_SLICE_X84Y102_B = CLBLM_L_X56Y102_SLICE_X84Y102_BO6;
  assign CLBLM_L_X56Y102_SLICE_X84Y102_C = CLBLM_L_X56Y102_SLICE_X84Y102_CO6;
  assign CLBLM_L_X56Y102_SLICE_X84Y102_D = CLBLM_L_X56Y102_SLICE_X84Y102_DO6;
  assign CLBLM_L_X56Y102_SLICE_X85Y102_A = CLBLM_L_X56Y102_SLICE_X85Y102_AO6;
  assign CLBLM_L_X56Y102_SLICE_X85Y102_B = CLBLM_L_X56Y102_SLICE_X85Y102_BO6;
  assign CLBLM_L_X56Y102_SLICE_X85Y102_C = CLBLM_L_X56Y102_SLICE_X85Y102_CO6;
  assign CLBLM_L_X56Y102_SLICE_X85Y102_D = CLBLM_L_X56Y102_SLICE_X85Y102_DO6;
  assign CLBLM_L_X56Y102_SLICE_X85Y102_AMUX = CLBLM_L_X56Y102_SLICE_X85Y102_A5Q;
  assign CLBLM_L_X56Y103_SLICE_X84Y103_A = CLBLM_L_X56Y103_SLICE_X84Y103_AO6;
  assign CLBLM_L_X56Y103_SLICE_X84Y103_B = CLBLM_L_X56Y103_SLICE_X84Y103_BO6;
  assign CLBLM_L_X56Y103_SLICE_X84Y103_C = CLBLM_L_X56Y103_SLICE_X84Y103_CO6;
  assign CLBLM_L_X56Y103_SLICE_X84Y103_D = CLBLM_L_X56Y103_SLICE_X84Y103_DO6;
  assign CLBLM_L_X56Y103_SLICE_X85Y103_A = CLBLM_L_X56Y103_SLICE_X85Y103_AO6;
  assign CLBLM_L_X56Y103_SLICE_X85Y103_B = CLBLM_L_X56Y103_SLICE_X85Y103_BO6;
  assign CLBLM_L_X56Y103_SLICE_X85Y103_C = CLBLM_L_X56Y103_SLICE_X85Y103_CO6;
  assign CLBLM_L_X56Y103_SLICE_X85Y103_D = CLBLM_L_X56Y103_SLICE_X85Y103_DO6;
  assign CLBLM_L_X56Y104_SLICE_X84Y104_A = CLBLM_L_X56Y104_SLICE_X84Y104_AO6;
  assign CLBLM_L_X56Y104_SLICE_X84Y104_B = CLBLM_L_X56Y104_SLICE_X84Y104_BO6;
  assign CLBLM_L_X56Y104_SLICE_X84Y104_C = CLBLM_L_X56Y104_SLICE_X84Y104_CO6;
  assign CLBLM_L_X56Y104_SLICE_X84Y104_D = CLBLM_L_X56Y104_SLICE_X84Y104_DO6;
  assign CLBLM_L_X56Y104_SLICE_X85Y104_A = CLBLM_L_X56Y104_SLICE_X85Y104_AO6;
  assign CLBLM_L_X56Y104_SLICE_X85Y104_B = CLBLM_L_X56Y104_SLICE_X85Y104_BO6;
  assign CLBLM_L_X56Y104_SLICE_X85Y104_C = CLBLM_L_X56Y104_SLICE_X85Y104_CO6;
  assign CLBLM_L_X56Y104_SLICE_X85Y104_D = CLBLM_L_X56Y104_SLICE_X85Y104_DO6;
  assign CLBLM_L_X56Y105_SLICE_X84Y105_A = CLBLM_L_X56Y105_SLICE_X84Y105_AO6;
  assign CLBLM_L_X56Y105_SLICE_X84Y105_B = CLBLM_L_X56Y105_SLICE_X84Y105_BO6;
  assign CLBLM_L_X56Y105_SLICE_X84Y105_C = CLBLM_L_X56Y105_SLICE_X84Y105_CO6;
  assign CLBLM_L_X56Y105_SLICE_X84Y105_D = CLBLM_L_X56Y105_SLICE_X84Y105_DO6;
  assign CLBLM_L_X56Y105_SLICE_X85Y105_A = CLBLM_L_X56Y105_SLICE_X85Y105_AO6;
  assign CLBLM_L_X56Y105_SLICE_X85Y105_B = CLBLM_L_X56Y105_SLICE_X85Y105_BO6;
  assign CLBLM_L_X56Y105_SLICE_X85Y105_C = CLBLM_L_X56Y105_SLICE_X85Y105_CO6;
  assign CLBLM_L_X56Y105_SLICE_X85Y105_D = CLBLM_L_X56Y105_SLICE_X85Y105_DO6;
  assign CLBLM_L_X56Y111_SLICE_X84Y111_A = CLBLM_L_X56Y111_SLICE_X84Y111_AO6;
  assign CLBLM_L_X56Y111_SLICE_X84Y111_B = CLBLM_L_X56Y111_SLICE_X84Y111_BO6;
  assign CLBLM_L_X56Y111_SLICE_X84Y111_C = CLBLM_L_X56Y111_SLICE_X84Y111_CO6;
  assign CLBLM_L_X56Y111_SLICE_X84Y111_D = CLBLM_L_X56Y111_SLICE_X84Y111_DO6;
  assign CLBLM_L_X56Y111_SLICE_X85Y111_A = CLBLM_L_X56Y111_SLICE_X85Y111_AO6;
  assign CLBLM_L_X56Y111_SLICE_X85Y111_B = CLBLM_L_X56Y111_SLICE_X85Y111_BO6;
  assign CLBLM_L_X56Y111_SLICE_X85Y111_C = CLBLM_L_X56Y111_SLICE_X85Y111_CO6;
  assign CLBLM_L_X56Y111_SLICE_X85Y111_D = CLBLM_L_X56Y111_SLICE_X85Y111_DO6;
  assign CLBLM_L_X60Y96_SLICE_X90Y96_A = CLBLM_L_X60Y96_SLICE_X90Y96_AO6;
  assign CLBLM_L_X60Y96_SLICE_X90Y96_B = CLBLM_L_X60Y96_SLICE_X90Y96_BO6;
  assign CLBLM_L_X60Y96_SLICE_X90Y96_C = CLBLM_L_X60Y96_SLICE_X90Y96_CO6;
  assign CLBLM_L_X60Y96_SLICE_X90Y96_D = CLBLM_L_X60Y96_SLICE_X90Y96_DO6;
  assign CLBLM_L_X60Y96_SLICE_X91Y96_A = CLBLM_L_X60Y96_SLICE_X91Y96_AO6;
  assign CLBLM_L_X60Y96_SLICE_X91Y96_B = CLBLM_L_X60Y96_SLICE_X91Y96_BO6;
  assign CLBLM_L_X60Y96_SLICE_X91Y96_C = CLBLM_L_X60Y96_SLICE_X91Y96_CO6;
  assign CLBLM_L_X60Y96_SLICE_X91Y96_D = CLBLM_L_X60Y96_SLICE_X91Y96_DO6;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_A = CLBLM_L_X60Y97_SLICE_X90Y97_AO6;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_B = CLBLM_L_X60Y97_SLICE_X90Y97_BO6;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_C = CLBLM_L_X60Y97_SLICE_X90Y97_CO6;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_D = CLBLM_L_X60Y97_SLICE_X90Y97_DO6;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_AMUX = CLBLM_L_X60Y97_SLICE_X90Y97_A5Q;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_A = CLBLM_L_X60Y97_SLICE_X91Y97_AO6;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_B = CLBLM_L_X60Y97_SLICE_X91Y97_BO6;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_C = CLBLM_L_X60Y97_SLICE_X91Y97_CO6;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_D = CLBLM_L_X60Y97_SLICE_X91Y97_DO6;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_AMUX = CLBLM_L_X60Y97_SLICE_X91Y97_AO5;
  assign CLBLM_L_X60Y98_SLICE_X90Y98_A = CLBLM_L_X60Y98_SLICE_X90Y98_AO6;
  assign CLBLM_L_X60Y98_SLICE_X90Y98_B = CLBLM_L_X60Y98_SLICE_X90Y98_BO6;
  assign CLBLM_L_X60Y98_SLICE_X90Y98_C = CLBLM_L_X60Y98_SLICE_X90Y98_CO6;
  assign CLBLM_L_X60Y98_SLICE_X90Y98_D = CLBLM_L_X60Y98_SLICE_X90Y98_DO6;
  assign CLBLM_L_X60Y98_SLICE_X90Y98_CMUX = CLBLM_L_X60Y98_SLICE_X90Y98_CO5;
  assign CLBLM_L_X60Y98_SLICE_X91Y98_A = CLBLM_L_X60Y98_SLICE_X91Y98_AO6;
  assign CLBLM_L_X60Y98_SLICE_X91Y98_B = CLBLM_L_X60Y98_SLICE_X91Y98_BO6;
  assign CLBLM_L_X60Y98_SLICE_X91Y98_C = CLBLM_L_X60Y98_SLICE_X91Y98_CO6;
  assign CLBLM_L_X60Y98_SLICE_X91Y98_D = CLBLM_L_X60Y98_SLICE_X91Y98_DO6;
  assign CLBLM_L_X60Y98_SLICE_X91Y98_AMUX = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_A = CLBLM_L_X60Y99_SLICE_X90Y99_AO6;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_B = CLBLM_L_X60Y99_SLICE_X90Y99_BO6;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_C = CLBLM_L_X60Y99_SLICE_X90Y99_CO6;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_D = CLBLM_L_X60Y99_SLICE_X90Y99_DO6;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_AMUX = CLBLM_L_X60Y99_SLICE_X90Y99_AO5;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_BMUX = CLBLM_L_X60Y99_SLICE_X90Y99_BO5;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_A = CLBLM_L_X60Y99_SLICE_X91Y99_AO6;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_B = CLBLM_L_X60Y99_SLICE_X91Y99_BO6;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_C = CLBLM_L_X60Y99_SLICE_X91Y99_CO6;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_D = CLBLM_L_X60Y99_SLICE_X91Y99_DO6;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_AMUX = CLBLM_L_X60Y99_SLICE_X91Y99_AO5;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_BMUX = CLBLM_L_X60Y99_SLICE_X91Y99_BO5;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_CMUX = CLBLM_L_X60Y99_SLICE_X91Y99_CO6;
  assign CLBLM_L_X60Y100_SLICE_X90Y100_A = CLBLM_L_X60Y100_SLICE_X90Y100_AO6;
  assign CLBLM_L_X60Y100_SLICE_X90Y100_B = CLBLM_L_X60Y100_SLICE_X90Y100_BO6;
  assign CLBLM_L_X60Y100_SLICE_X90Y100_C = CLBLM_L_X60Y100_SLICE_X90Y100_CO6;
  assign CLBLM_L_X60Y100_SLICE_X90Y100_D = CLBLM_L_X60Y100_SLICE_X90Y100_DO6;
  assign CLBLM_L_X60Y100_SLICE_X90Y100_AMUX = CLBLM_L_X60Y100_SLICE_X90Y100_AO5;
  assign CLBLM_L_X60Y100_SLICE_X91Y100_A = CLBLM_L_X60Y100_SLICE_X91Y100_AO6;
  assign CLBLM_L_X60Y100_SLICE_X91Y100_B = CLBLM_L_X60Y100_SLICE_X91Y100_BO6;
  assign CLBLM_L_X60Y100_SLICE_X91Y100_C = CLBLM_L_X60Y100_SLICE_X91Y100_CO6;
  assign CLBLM_L_X60Y100_SLICE_X91Y100_D = CLBLM_L_X60Y100_SLICE_X91Y100_DO6;
  assign CLBLM_L_X60Y100_SLICE_X91Y100_AMUX = CLBLM_L_X60Y100_SLICE_X91Y100_AO5;
  assign CLBLM_L_X60Y100_SLICE_X91Y100_CMUX = CLBLM_L_X60Y100_SLICE_X91Y100_CO5;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_A = CLBLM_L_X60Y101_SLICE_X90Y101_AO6;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_B = CLBLM_L_X60Y101_SLICE_X90Y101_BO6;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_C = CLBLM_L_X60Y101_SLICE_X90Y101_CO6;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_D = CLBLM_L_X60Y101_SLICE_X90Y101_DO6;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_A = CLBLM_L_X60Y101_SLICE_X91Y101_AO6;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_B = CLBLM_L_X60Y101_SLICE_X91Y101_BO6;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_C = CLBLM_L_X60Y101_SLICE_X91Y101_CO6;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_D = CLBLM_L_X60Y101_SLICE_X91Y101_DO6;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_CMUX = CLBLM_L_X60Y101_SLICE_X91Y101_CO5;
  assign CLBLM_L_X60Y102_SLICE_X90Y102_A = CLBLM_L_X60Y102_SLICE_X90Y102_AO6;
  assign CLBLM_L_X60Y102_SLICE_X90Y102_B = CLBLM_L_X60Y102_SLICE_X90Y102_BO6;
  assign CLBLM_L_X60Y102_SLICE_X90Y102_C = CLBLM_L_X60Y102_SLICE_X90Y102_CO6;
  assign CLBLM_L_X60Y102_SLICE_X90Y102_D = CLBLM_L_X60Y102_SLICE_X90Y102_DO6;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_A = CLBLM_L_X60Y102_SLICE_X91Y102_AO6;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_B = CLBLM_L_X60Y102_SLICE_X91Y102_BO6;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_C = CLBLM_L_X60Y102_SLICE_X91Y102_CO6;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_D = CLBLM_L_X60Y102_SLICE_X91Y102_DO6;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_AMUX = CLBLM_L_X60Y102_SLICE_X91Y102_A_XOR;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_BMUX = CLBLM_L_X60Y102_SLICE_X91Y102_B_XOR;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_CMUX = CLBLM_L_X60Y102_SLICE_X91Y102_C_XOR;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_DMUX = CLBLM_L_X60Y102_SLICE_X91Y102_D_XOR;
  assign CLBLM_L_X60Y103_SLICE_X90Y103_A = CLBLM_L_X60Y103_SLICE_X90Y103_AO6;
  assign CLBLM_L_X60Y103_SLICE_X90Y103_B = CLBLM_L_X60Y103_SLICE_X90Y103_BO6;
  assign CLBLM_L_X60Y103_SLICE_X90Y103_C = CLBLM_L_X60Y103_SLICE_X90Y103_CO6;
  assign CLBLM_L_X60Y103_SLICE_X90Y103_D = CLBLM_L_X60Y103_SLICE_X90Y103_DO6;
  assign CLBLM_L_X60Y103_SLICE_X90Y103_BMUX = CLBLM_L_X60Y103_SLICE_X90Y103_F8MUX_O;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_A = CLBLM_L_X60Y103_SLICE_X91Y103_AO6;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_B = CLBLM_L_X60Y103_SLICE_X91Y103_BO6;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_C = CLBLM_L_X60Y103_SLICE_X91Y103_CO6;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_D = CLBLM_L_X60Y103_SLICE_X91Y103_DO6;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_AMUX = CLBLM_L_X60Y103_SLICE_X91Y103_A_XOR;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_BMUX = CLBLM_L_X60Y103_SLICE_X91Y103_B_XOR;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_CMUX = CLBLM_L_X60Y103_SLICE_X91Y103_C_XOR;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_DMUX = CLBLM_L_X60Y103_SLICE_X91Y103_D_XOR;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_A = CLBLM_L_X60Y104_SLICE_X90Y104_AO6;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_B = CLBLM_L_X60Y104_SLICE_X90Y104_BO6;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_C = CLBLM_L_X60Y104_SLICE_X90Y104_CO6;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_D = CLBLM_L_X60Y104_SLICE_X90Y104_DO6;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_A = CLBLM_L_X60Y104_SLICE_X91Y104_AO6;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_B = CLBLM_L_X60Y104_SLICE_X91Y104_BO6;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_C = CLBLM_L_X60Y104_SLICE_X91Y104_CO6;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_D = CLBLM_L_X60Y104_SLICE_X91Y104_DO6;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_AMUX = CLBLM_L_X60Y104_SLICE_X91Y104_A_XOR;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_BMUX = CLBLM_L_X60Y104_SLICE_X91Y104_B_XOR;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_CMUX = CLBLM_L_X60Y104_SLICE_X91Y104_C_XOR;
  assign CLBLM_L_X60Y105_SLICE_X90Y105_A = CLBLM_L_X60Y105_SLICE_X90Y105_AO6;
  assign CLBLM_L_X60Y105_SLICE_X90Y105_B = CLBLM_L_X60Y105_SLICE_X90Y105_BO6;
  assign CLBLM_L_X60Y105_SLICE_X90Y105_C = CLBLM_L_X60Y105_SLICE_X90Y105_CO6;
  assign CLBLM_L_X60Y105_SLICE_X90Y105_D = CLBLM_L_X60Y105_SLICE_X90Y105_DO6;
  assign CLBLM_L_X60Y105_SLICE_X90Y105_AMUX = CLBLM_L_X60Y105_SLICE_X90Y105_A_XOR;
  assign CLBLM_L_X60Y105_SLICE_X90Y105_BMUX = CLBLM_L_X60Y105_SLICE_X90Y105_B_XOR;
  assign CLBLM_L_X60Y105_SLICE_X90Y105_CMUX = CLBLM_L_X60Y105_SLICE_X90Y105_C_XOR;
  assign CLBLM_L_X60Y105_SLICE_X90Y105_DMUX = CLBLM_L_X60Y105_SLICE_X90Y105_D_XOR;
  assign CLBLM_L_X60Y105_SLICE_X91Y105_A = CLBLM_L_X60Y105_SLICE_X91Y105_AO6;
  assign CLBLM_L_X60Y105_SLICE_X91Y105_B = CLBLM_L_X60Y105_SLICE_X91Y105_BO6;
  assign CLBLM_L_X60Y105_SLICE_X91Y105_C = CLBLM_L_X60Y105_SLICE_X91Y105_CO6;
  assign CLBLM_L_X60Y105_SLICE_X91Y105_D = CLBLM_L_X60Y105_SLICE_X91Y105_DO6;
  assign CLBLM_L_X60Y105_SLICE_X91Y105_AMUX = CLBLM_L_X60Y105_SLICE_X91Y105_A_XOR;
  assign CLBLM_L_X60Y105_SLICE_X91Y105_BMUX = CLBLM_L_X60Y105_SLICE_X91Y105_B_XOR;
  assign CLBLM_L_X60Y105_SLICE_X91Y105_CMUX = CLBLM_L_X60Y105_SLICE_X91Y105_C_XOR;
  assign CLBLM_L_X60Y105_SLICE_X91Y105_DMUX = CLBLM_L_X60Y105_SLICE_X91Y105_D_XOR;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_A = CLBLM_L_X60Y106_SLICE_X90Y106_AO6;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_B = CLBLM_L_X60Y106_SLICE_X90Y106_BO6;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_C = CLBLM_L_X60Y106_SLICE_X90Y106_CO6;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_D = CLBLM_L_X60Y106_SLICE_X90Y106_DO6;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_AMUX = CLBLM_L_X60Y106_SLICE_X90Y106_A_XOR;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_BMUX = CLBLM_L_X60Y106_SLICE_X90Y106_B_XOR;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_CMUX = CLBLM_L_X60Y106_SLICE_X90Y106_C_XOR;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_DMUX = CLBLM_L_X60Y106_SLICE_X90Y106_D_XOR;
  assign CLBLM_L_X60Y106_SLICE_X91Y106_A = CLBLM_L_X60Y106_SLICE_X91Y106_AO6;
  assign CLBLM_L_X60Y106_SLICE_X91Y106_B = CLBLM_L_X60Y106_SLICE_X91Y106_BO6;
  assign CLBLM_L_X60Y106_SLICE_X91Y106_C = CLBLM_L_X60Y106_SLICE_X91Y106_CO6;
  assign CLBLM_L_X60Y106_SLICE_X91Y106_D = CLBLM_L_X60Y106_SLICE_X91Y106_DO6;
  assign CLBLM_L_X60Y106_SLICE_X91Y106_AMUX = CLBLM_L_X60Y106_SLICE_X91Y106_A_XOR;
  assign CLBLM_L_X60Y106_SLICE_X91Y106_BMUX = CLBLM_L_X60Y106_SLICE_X91Y106_B_XOR;
  assign CLBLM_L_X60Y106_SLICE_X91Y106_CMUX = CLBLM_L_X60Y106_SLICE_X91Y106_C_XOR;
  assign CLBLM_L_X60Y106_SLICE_X91Y106_DMUX = CLBLM_L_X60Y106_SLICE_X91Y106_D_XOR;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_A = CLBLM_L_X60Y107_SLICE_X90Y107_AO6;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_B = CLBLM_L_X60Y107_SLICE_X90Y107_BO6;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_C = CLBLM_L_X60Y107_SLICE_X90Y107_CO6;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_D = CLBLM_L_X60Y107_SLICE_X90Y107_DO6;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_AMUX = CLBLM_L_X60Y107_SLICE_X90Y107_A_XOR;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_BMUX = CLBLM_L_X60Y107_SLICE_X90Y107_B_XOR;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_CMUX = CLBLM_L_X60Y107_SLICE_X90Y107_C_XOR;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_DMUX = CLBLM_L_X60Y107_SLICE_X90Y107_D_XOR;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_A = CLBLM_L_X60Y107_SLICE_X91Y107_AO6;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_B = CLBLM_L_X60Y107_SLICE_X91Y107_BO6;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_C = CLBLM_L_X60Y107_SLICE_X91Y107_CO6;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_D = CLBLM_L_X60Y107_SLICE_X91Y107_DO6;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_AMUX = CLBLM_L_X60Y107_SLICE_X91Y107_A_XOR;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_BMUX = CLBLM_L_X60Y107_SLICE_X91Y107_B_XOR;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_CMUX = CLBLM_L_X60Y107_SLICE_X91Y107_C_XOR;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_A = CLBLM_L_X60Y108_SLICE_X90Y108_AO6;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_B = CLBLM_L_X60Y108_SLICE_X90Y108_BO6;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_C = CLBLM_L_X60Y108_SLICE_X90Y108_CO6;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_D = CLBLM_L_X60Y108_SLICE_X90Y108_DO6;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_AMUX = CLBLM_L_X60Y108_SLICE_X90Y108_A_XOR;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_BMUX = CLBLM_L_X60Y108_SLICE_X90Y108_B_XOR;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_CMUX = CLBLM_L_X60Y108_SLICE_X90Y108_C_XOR;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_DMUX = CLBLM_L_X60Y108_SLICE_X90Y108_D_XOR;
  assign CLBLM_L_X60Y108_SLICE_X91Y108_A = CLBLM_L_X60Y108_SLICE_X91Y108_AO6;
  assign CLBLM_L_X60Y108_SLICE_X91Y108_B = CLBLM_L_X60Y108_SLICE_X91Y108_BO6;
  assign CLBLM_L_X60Y108_SLICE_X91Y108_C = CLBLM_L_X60Y108_SLICE_X91Y108_CO6;
  assign CLBLM_L_X60Y108_SLICE_X91Y108_D = CLBLM_L_X60Y108_SLICE_X91Y108_DO6;
  assign CLBLM_L_X60Y109_SLICE_X90Y109_A = CLBLM_L_X60Y109_SLICE_X90Y109_AO6;
  assign CLBLM_L_X60Y109_SLICE_X90Y109_B = CLBLM_L_X60Y109_SLICE_X90Y109_BO6;
  assign CLBLM_L_X60Y109_SLICE_X90Y109_C = CLBLM_L_X60Y109_SLICE_X90Y109_CO6;
  assign CLBLM_L_X60Y109_SLICE_X90Y109_D = CLBLM_L_X60Y109_SLICE_X90Y109_DO6;
  assign CLBLM_L_X60Y109_SLICE_X90Y109_AMUX = CLBLM_L_X60Y109_SLICE_X90Y109_A_XOR;
  assign CLBLM_L_X60Y109_SLICE_X90Y109_BMUX = CLBLM_L_X60Y109_SLICE_X90Y109_B_XOR;
  assign CLBLM_L_X60Y109_SLICE_X90Y109_CMUX = CLBLM_L_X60Y109_SLICE_X90Y109_C_XOR;
  assign CLBLM_L_X60Y109_SLICE_X90Y109_DMUX = CLBLM_L_X60Y109_SLICE_X90Y109_D_XOR;
  assign CLBLM_L_X60Y109_SLICE_X91Y109_A = CLBLM_L_X60Y109_SLICE_X91Y109_AO6;
  assign CLBLM_L_X60Y109_SLICE_X91Y109_B = CLBLM_L_X60Y109_SLICE_X91Y109_BO6;
  assign CLBLM_L_X60Y109_SLICE_X91Y109_C = CLBLM_L_X60Y109_SLICE_X91Y109_CO6;
  assign CLBLM_L_X60Y109_SLICE_X91Y109_D = CLBLM_L_X60Y109_SLICE_X91Y109_DO6;
  assign CLBLM_L_X60Y110_SLICE_X90Y110_A = CLBLM_L_X60Y110_SLICE_X90Y110_AO6;
  assign CLBLM_L_X60Y110_SLICE_X90Y110_B = CLBLM_L_X60Y110_SLICE_X90Y110_BO6;
  assign CLBLM_L_X60Y110_SLICE_X90Y110_C = CLBLM_L_X60Y110_SLICE_X90Y110_CO6;
  assign CLBLM_L_X60Y110_SLICE_X90Y110_D = CLBLM_L_X60Y110_SLICE_X90Y110_DO6;
  assign CLBLM_L_X60Y110_SLICE_X90Y110_AMUX = CLBLM_L_X60Y110_SLICE_X90Y110_A_XOR;
  assign CLBLM_L_X60Y110_SLICE_X90Y110_BMUX = CLBLM_L_X60Y110_SLICE_X90Y110_B_XOR;
  assign CLBLM_L_X60Y110_SLICE_X90Y110_CMUX = CLBLM_L_X60Y110_SLICE_X90Y110_C_XOR;
  assign CLBLM_L_X60Y110_SLICE_X91Y110_A = CLBLM_L_X60Y110_SLICE_X91Y110_AO6;
  assign CLBLM_L_X60Y110_SLICE_X91Y110_B = CLBLM_L_X60Y110_SLICE_X91Y110_BO6;
  assign CLBLM_L_X60Y110_SLICE_X91Y110_C = CLBLM_L_X60Y110_SLICE_X91Y110_CO6;
  assign CLBLM_L_X60Y110_SLICE_X91Y110_D = CLBLM_L_X60Y110_SLICE_X91Y110_DO6;
  assign CLBLM_L_X60Y111_SLICE_X90Y111_A = CLBLM_L_X60Y111_SLICE_X90Y111_AO6;
  assign CLBLM_L_X60Y111_SLICE_X90Y111_B = CLBLM_L_X60Y111_SLICE_X90Y111_BO6;
  assign CLBLM_L_X60Y111_SLICE_X90Y111_C = CLBLM_L_X60Y111_SLICE_X90Y111_CO6;
  assign CLBLM_L_X60Y111_SLICE_X90Y111_D = CLBLM_L_X60Y111_SLICE_X90Y111_DO6;
  assign CLBLM_L_X60Y111_SLICE_X91Y111_A = CLBLM_L_X60Y111_SLICE_X91Y111_AO6;
  assign CLBLM_L_X60Y111_SLICE_X91Y111_B = CLBLM_L_X60Y111_SLICE_X91Y111_BO6;
  assign CLBLM_L_X60Y111_SLICE_X91Y111_C = CLBLM_L_X60Y111_SLICE_X91Y111_CO6;
  assign CLBLM_L_X60Y111_SLICE_X91Y111_D = CLBLM_L_X60Y111_SLICE_X91Y111_DO6;
  assign CLBLM_L_X60Y112_SLICE_X90Y112_A = CLBLM_L_X60Y112_SLICE_X90Y112_AO6;
  assign CLBLM_L_X60Y112_SLICE_X90Y112_B = CLBLM_L_X60Y112_SLICE_X90Y112_BO6;
  assign CLBLM_L_X60Y112_SLICE_X90Y112_C = CLBLM_L_X60Y112_SLICE_X90Y112_CO6;
  assign CLBLM_L_X60Y112_SLICE_X90Y112_D = CLBLM_L_X60Y112_SLICE_X90Y112_DO6;
  assign CLBLM_L_X60Y112_SLICE_X91Y112_A = CLBLM_L_X60Y112_SLICE_X91Y112_AO6;
  assign CLBLM_L_X60Y112_SLICE_X91Y112_B = CLBLM_L_X60Y112_SLICE_X91Y112_BO6;
  assign CLBLM_L_X60Y112_SLICE_X91Y112_C = CLBLM_L_X60Y112_SLICE_X91Y112_CO6;
  assign CLBLM_L_X60Y112_SLICE_X91Y112_D = CLBLM_L_X60Y112_SLICE_X91Y112_DO6;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_A = CLBLM_L_X62Y95_SLICE_X92Y95_AO6;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_B = CLBLM_L_X62Y95_SLICE_X92Y95_BO6;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_C = CLBLM_L_X62Y95_SLICE_X92Y95_CO6;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_D = CLBLM_L_X62Y95_SLICE_X92Y95_DO6;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_AMUX = CLBLM_L_X62Y95_SLICE_X92Y95_A5Q;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_A = CLBLM_L_X62Y95_SLICE_X93Y95_AO6;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_B = CLBLM_L_X62Y95_SLICE_X93Y95_BO6;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_C = CLBLM_L_X62Y95_SLICE_X93Y95_CO6;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_D = CLBLM_L_X62Y95_SLICE_X93Y95_DO6;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_AMUX = CLBLM_L_X62Y95_SLICE_X93Y95_AO5;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_BMUX = CLBLM_L_X62Y95_SLICE_X93Y95_BO5;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_DMUX = CLBLM_L_X62Y95_SLICE_X93Y95_D5Q;
  assign CLBLM_L_X62Y96_SLICE_X92Y96_A = CLBLM_L_X62Y96_SLICE_X92Y96_AO6;
  assign CLBLM_L_X62Y96_SLICE_X92Y96_B = CLBLM_L_X62Y96_SLICE_X92Y96_BO6;
  assign CLBLM_L_X62Y96_SLICE_X92Y96_C = CLBLM_L_X62Y96_SLICE_X92Y96_CO6;
  assign CLBLM_L_X62Y96_SLICE_X92Y96_D = CLBLM_L_X62Y96_SLICE_X92Y96_DO6;
  assign CLBLM_L_X62Y96_SLICE_X92Y96_AMUX = CLBLM_L_X62Y96_SLICE_X92Y96_F7AMUX_O;
  assign CLBLM_L_X62Y96_SLICE_X93Y96_A = CLBLM_L_X62Y96_SLICE_X93Y96_AO6;
  assign CLBLM_L_X62Y96_SLICE_X93Y96_B = CLBLM_L_X62Y96_SLICE_X93Y96_BO6;
  assign CLBLM_L_X62Y96_SLICE_X93Y96_C = CLBLM_L_X62Y96_SLICE_X93Y96_CO6;
  assign CLBLM_L_X62Y96_SLICE_X93Y96_D = CLBLM_L_X62Y96_SLICE_X93Y96_DO6;
  assign CLBLM_L_X62Y96_SLICE_X93Y96_AMUX = CLBLM_L_X62Y96_SLICE_X93Y96_F7AMUX_O;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_A = CLBLM_L_X62Y97_SLICE_X92Y97_AO6;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_B = CLBLM_L_X62Y97_SLICE_X92Y97_BO6;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_C = CLBLM_L_X62Y97_SLICE_X92Y97_CO6;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_D = CLBLM_L_X62Y97_SLICE_X92Y97_DO6;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_CMUX = CLBLM_L_X62Y97_SLICE_X92Y97_C5Q;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_DMUX = CLBLM_L_X62Y97_SLICE_X92Y97_D5Q;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_A = CLBLM_L_X62Y97_SLICE_X93Y97_AO6;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_B = CLBLM_L_X62Y97_SLICE_X93Y97_BO6;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_C = CLBLM_L_X62Y97_SLICE_X93Y97_CO6;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_D = CLBLM_L_X62Y97_SLICE_X93Y97_DO6;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_AMUX = CLBLM_L_X62Y97_SLICE_X93Y97_F7AMUX_O;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_CMUX = CLBLM_L_X62Y97_SLICE_X93Y97_CO5;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_A = CLBLM_L_X62Y98_SLICE_X92Y98_AO6;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_B = CLBLM_L_X62Y98_SLICE_X92Y98_BO6;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_C = CLBLM_L_X62Y98_SLICE_X92Y98_CO6;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_D = CLBLM_L_X62Y98_SLICE_X92Y98_DO6;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_A = CLBLM_L_X62Y98_SLICE_X93Y98_AO6;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_B = CLBLM_L_X62Y98_SLICE_X93Y98_BO6;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_C = CLBLM_L_X62Y98_SLICE_X93Y98_CO6;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_D = CLBLM_L_X62Y98_SLICE_X93Y98_DO6;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_A = CLBLM_L_X62Y99_SLICE_X92Y99_AO6;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_B = CLBLM_L_X62Y99_SLICE_X92Y99_BO6;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_C = CLBLM_L_X62Y99_SLICE_X92Y99_CO6;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_D = CLBLM_L_X62Y99_SLICE_X92Y99_DO6;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_AMUX = CLBLM_L_X62Y99_SLICE_X92Y99_AO5;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_A = CLBLM_L_X62Y99_SLICE_X93Y99_AO6;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_B = CLBLM_L_X62Y99_SLICE_X93Y99_BO6;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_C = CLBLM_L_X62Y99_SLICE_X93Y99_CO6;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_D = CLBLM_L_X62Y99_SLICE_X93Y99_DO6;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_BMUX = CLBLM_L_X62Y99_SLICE_X93Y99_BO6;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_A = CLBLM_L_X62Y100_SLICE_X92Y100_AO6;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_B = CLBLM_L_X62Y100_SLICE_X92Y100_BO6;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_C = CLBLM_L_X62Y100_SLICE_X92Y100_CO6;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_D = CLBLM_L_X62Y100_SLICE_X92Y100_DO6;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_AMUX = CLBLM_L_X62Y100_SLICE_X92Y100_AO5;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_A = CLBLM_L_X62Y100_SLICE_X93Y100_AO6;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_B = CLBLM_L_X62Y100_SLICE_X93Y100_BO6;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_C = CLBLM_L_X62Y100_SLICE_X93Y100_CO6;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_D = CLBLM_L_X62Y100_SLICE_X93Y100_DO6;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_A = CLBLM_L_X62Y101_SLICE_X92Y101_AO6;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_B = CLBLM_L_X62Y101_SLICE_X92Y101_BO6;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_C = CLBLM_L_X62Y101_SLICE_X92Y101_CO6;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_D = CLBLM_L_X62Y101_SLICE_X92Y101_DO6;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_DMUX = CLBLM_L_X62Y101_SLICE_X92Y101_DO5;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_A = CLBLM_L_X62Y101_SLICE_X93Y101_AO6;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_B = CLBLM_L_X62Y101_SLICE_X93Y101_BO6;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_C = CLBLM_L_X62Y101_SLICE_X93Y101_CO6;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_D = CLBLM_L_X62Y101_SLICE_X93Y101_DO6;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_A = CLBLM_L_X62Y102_SLICE_X92Y102_AO6;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_B = CLBLM_L_X62Y102_SLICE_X92Y102_BO6;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_C = CLBLM_L_X62Y102_SLICE_X92Y102_CO6;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_D = CLBLM_L_X62Y102_SLICE_X92Y102_DO6;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_AMUX = CLBLM_L_X62Y102_SLICE_X92Y102_AO5;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_DMUX = CLBLM_L_X62Y102_SLICE_X92Y102_DO6;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_A = CLBLM_L_X62Y102_SLICE_X93Y102_AO6;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_B = CLBLM_L_X62Y102_SLICE_X93Y102_BO6;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_C = CLBLM_L_X62Y102_SLICE_X93Y102_CO6;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_D = CLBLM_L_X62Y102_SLICE_X93Y102_DO6;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_AMUX = CLBLM_L_X62Y102_SLICE_X93Y102_AO5;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_A = CLBLM_L_X62Y103_SLICE_X92Y103_AO6;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_B = CLBLM_L_X62Y103_SLICE_X92Y103_BO6;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_C = CLBLM_L_X62Y103_SLICE_X92Y103_CO6;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_D = CLBLM_L_X62Y103_SLICE_X92Y103_DO6;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_CMUX = CLBLM_L_X62Y103_SLICE_X92Y103_CO6;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_A = CLBLM_L_X62Y103_SLICE_X93Y103_AO6;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_B = CLBLM_L_X62Y103_SLICE_X93Y103_BO6;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_C = CLBLM_L_X62Y103_SLICE_X93Y103_CO6;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_D = CLBLM_L_X62Y103_SLICE_X93Y103_DO6;
  assign CLBLM_L_X62Y104_SLICE_X92Y104_A = CLBLM_L_X62Y104_SLICE_X92Y104_AO6;
  assign CLBLM_L_X62Y104_SLICE_X92Y104_B = CLBLM_L_X62Y104_SLICE_X92Y104_BO6;
  assign CLBLM_L_X62Y104_SLICE_X92Y104_C = CLBLM_L_X62Y104_SLICE_X92Y104_CO6;
  assign CLBLM_L_X62Y104_SLICE_X92Y104_D = CLBLM_L_X62Y104_SLICE_X92Y104_DO6;
  assign CLBLM_L_X62Y104_SLICE_X92Y104_CMUX = CLBLM_L_X62Y104_SLICE_X92Y104_CO6;
  assign CLBLM_L_X62Y104_SLICE_X93Y104_A = CLBLM_L_X62Y104_SLICE_X93Y104_AO6;
  assign CLBLM_L_X62Y104_SLICE_X93Y104_B = CLBLM_L_X62Y104_SLICE_X93Y104_BO6;
  assign CLBLM_L_X62Y104_SLICE_X93Y104_C = CLBLM_L_X62Y104_SLICE_X93Y104_CO6;
  assign CLBLM_L_X62Y104_SLICE_X93Y104_D = CLBLM_L_X62Y104_SLICE_X93Y104_DO6;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_A = CLBLM_L_X62Y105_SLICE_X92Y105_AO6;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_B = CLBLM_L_X62Y105_SLICE_X92Y105_BO6;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_C = CLBLM_L_X62Y105_SLICE_X92Y105_CO6;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_D = CLBLM_L_X62Y105_SLICE_X92Y105_DO6;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_AMUX = CLBLM_L_X62Y105_SLICE_X92Y105_AO5;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_BMUX = CLBLM_L_X62Y105_SLICE_X92Y105_BO5;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_A = CLBLM_L_X62Y105_SLICE_X93Y105_AO6;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_B = CLBLM_L_X62Y105_SLICE_X93Y105_BO6;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_C = CLBLM_L_X62Y105_SLICE_X93Y105_CO6;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_D = CLBLM_L_X62Y105_SLICE_X93Y105_DO6;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_AMUX = CLBLM_L_X62Y105_SLICE_X93Y105_AO5;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_A = CLBLM_L_X62Y106_SLICE_X92Y106_AO6;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_B = CLBLM_L_X62Y106_SLICE_X92Y106_BO6;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_C = CLBLM_L_X62Y106_SLICE_X92Y106_CO6;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_D = CLBLM_L_X62Y106_SLICE_X92Y106_DO6;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_AMUX = CLBLM_L_X62Y106_SLICE_X92Y106_AO5;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_A = CLBLM_L_X62Y106_SLICE_X93Y106_AO6;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_B = CLBLM_L_X62Y106_SLICE_X93Y106_BO6;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_C = CLBLM_L_X62Y106_SLICE_X93Y106_CO6;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_D = CLBLM_L_X62Y106_SLICE_X93Y106_DO6;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_BMUX = CLBLM_L_X62Y106_SLICE_X93Y106_BO5;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_CMUX = CLBLM_L_X62Y106_SLICE_X93Y106_CO6;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_A = CLBLM_L_X62Y107_SLICE_X92Y107_AO6;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_B = CLBLM_L_X62Y107_SLICE_X92Y107_BO6;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_C = CLBLM_L_X62Y107_SLICE_X92Y107_CO6;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_D = CLBLM_L_X62Y107_SLICE_X92Y107_DO6;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_AMUX = CLBLM_L_X62Y107_SLICE_X92Y107_A5Q;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_BMUX = CLBLM_L_X62Y107_SLICE_X92Y107_BO5;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_A = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_B = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_C = CLBLM_L_X62Y107_SLICE_X93Y107_CO6;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_D = CLBLM_L_X62Y107_SLICE_X93Y107_DO6;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_BMUX = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_L_X62Y108_SLICE_X92Y108_A = CLBLM_L_X62Y108_SLICE_X92Y108_AO6;
  assign CLBLM_L_X62Y108_SLICE_X92Y108_B = CLBLM_L_X62Y108_SLICE_X92Y108_BO6;
  assign CLBLM_L_X62Y108_SLICE_X92Y108_C = CLBLM_L_X62Y108_SLICE_X92Y108_CO6;
  assign CLBLM_L_X62Y108_SLICE_X92Y108_D = CLBLM_L_X62Y108_SLICE_X92Y108_DO6;
  assign CLBLM_L_X62Y108_SLICE_X92Y108_AMUX = CLBLM_L_X62Y108_SLICE_X92Y108_A5Q;
  assign CLBLM_L_X62Y108_SLICE_X92Y108_BMUX = CLBLM_L_X62Y108_SLICE_X92Y108_BO5;
  assign CLBLM_L_X62Y108_SLICE_X93Y108_A = CLBLM_L_X62Y108_SLICE_X93Y108_AO6;
  assign CLBLM_L_X62Y108_SLICE_X93Y108_B = CLBLM_L_X62Y108_SLICE_X93Y108_BO6;
  assign CLBLM_L_X62Y108_SLICE_X93Y108_C = CLBLM_L_X62Y108_SLICE_X93Y108_CO6;
  assign CLBLM_L_X62Y108_SLICE_X93Y108_D = CLBLM_L_X62Y108_SLICE_X93Y108_DO6;
  assign CLBLM_L_X62Y109_SLICE_X92Y109_A = CLBLM_L_X62Y109_SLICE_X92Y109_AO6;
  assign CLBLM_L_X62Y109_SLICE_X92Y109_B = CLBLM_L_X62Y109_SLICE_X92Y109_BO6;
  assign CLBLM_L_X62Y109_SLICE_X92Y109_C = CLBLM_L_X62Y109_SLICE_X92Y109_CO6;
  assign CLBLM_L_X62Y109_SLICE_X92Y109_D = CLBLM_L_X62Y109_SLICE_X92Y109_DO6;
  assign CLBLM_L_X62Y109_SLICE_X93Y109_A = CLBLM_L_X62Y109_SLICE_X93Y109_AO6;
  assign CLBLM_L_X62Y109_SLICE_X93Y109_B = CLBLM_L_X62Y109_SLICE_X93Y109_BO6;
  assign CLBLM_L_X62Y109_SLICE_X93Y109_C = CLBLM_L_X62Y109_SLICE_X93Y109_CO6;
  assign CLBLM_L_X62Y109_SLICE_X93Y109_D = CLBLM_L_X62Y109_SLICE_X93Y109_DO6;
  assign CLBLM_L_X62Y110_SLICE_X92Y110_A = CLBLM_L_X62Y110_SLICE_X92Y110_AO6;
  assign CLBLM_L_X62Y110_SLICE_X92Y110_B = CLBLM_L_X62Y110_SLICE_X92Y110_BO6;
  assign CLBLM_L_X62Y110_SLICE_X92Y110_C = CLBLM_L_X62Y110_SLICE_X92Y110_CO6;
  assign CLBLM_L_X62Y110_SLICE_X92Y110_D = CLBLM_L_X62Y110_SLICE_X92Y110_DO6;
  assign CLBLM_L_X62Y110_SLICE_X93Y110_A = CLBLM_L_X62Y110_SLICE_X93Y110_AO6;
  assign CLBLM_L_X62Y110_SLICE_X93Y110_B = CLBLM_L_X62Y110_SLICE_X93Y110_BO6;
  assign CLBLM_L_X62Y110_SLICE_X93Y110_C = CLBLM_L_X62Y110_SLICE_X93Y110_CO6;
  assign CLBLM_L_X62Y110_SLICE_X93Y110_D = CLBLM_L_X62Y110_SLICE_X93Y110_DO6;
  assign CLBLM_L_X62Y110_SLICE_X93Y110_CMUX = CLBLM_L_X62Y110_SLICE_X93Y110_CO6;
  assign CLBLM_L_X62Y111_SLICE_X92Y111_A = CLBLM_L_X62Y111_SLICE_X92Y111_AO6;
  assign CLBLM_L_X62Y111_SLICE_X92Y111_B = CLBLM_L_X62Y111_SLICE_X92Y111_BO6;
  assign CLBLM_L_X62Y111_SLICE_X92Y111_C = CLBLM_L_X62Y111_SLICE_X92Y111_CO6;
  assign CLBLM_L_X62Y111_SLICE_X92Y111_D = CLBLM_L_X62Y111_SLICE_X92Y111_DO6;
  assign CLBLM_L_X62Y111_SLICE_X92Y111_AMUX = CLBLM_L_X62Y111_SLICE_X92Y111_A5Q;
  assign CLBLM_L_X62Y111_SLICE_X93Y111_A = CLBLM_L_X62Y111_SLICE_X93Y111_AO6;
  assign CLBLM_L_X62Y111_SLICE_X93Y111_B = CLBLM_L_X62Y111_SLICE_X93Y111_BO6;
  assign CLBLM_L_X62Y111_SLICE_X93Y111_C = CLBLM_L_X62Y111_SLICE_X93Y111_CO6;
  assign CLBLM_L_X62Y111_SLICE_X93Y111_D = CLBLM_L_X62Y111_SLICE_X93Y111_DO6;
  assign CLBLM_L_X62Y112_SLICE_X92Y112_A = CLBLM_L_X62Y112_SLICE_X92Y112_AO6;
  assign CLBLM_L_X62Y112_SLICE_X92Y112_B = CLBLM_L_X62Y112_SLICE_X92Y112_BO6;
  assign CLBLM_L_X62Y112_SLICE_X92Y112_C = CLBLM_L_X62Y112_SLICE_X92Y112_CO6;
  assign CLBLM_L_X62Y112_SLICE_X92Y112_D = CLBLM_L_X62Y112_SLICE_X92Y112_DO6;
  assign CLBLM_L_X62Y112_SLICE_X93Y112_A = CLBLM_L_X62Y112_SLICE_X93Y112_AO6;
  assign CLBLM_L_X62Y112_SLICE_X93Y112_B = CLBLM_L_X62Y112_SLICE_X93Y112_BO6;
  assign CLBLM_L_X62Y112_SLICE_X93Y112_C = CLBLM_L_X62Y112_SLICE_X93Y112_CO6;
  assign CLBLM_L_X62Y112_SLICE_X93Y112_D = CLBLM_L_X62Y112_SLICE_X93Y112_DO6;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_A = CLBLM_L_X64Y95_SLICE_X96Y95_AO6;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_B = CLBLM_L_X64Y95_SLICE_X96Y95_BO6;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_C = CLBLM_L_X64Y95_SLICE_X96Y95_CO6;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_D = CLBLM_L_X64Y95_SLICE_X96Y95_DO6;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_AMUX = CLBLM_L_X64Y95_SLICE_X96Y95_AO5;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_BMUX = CLBLM_L_X64Y95_SLICE_X96Y95_BO5;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_CMUX = CLBLM_L_X64Y95_SLICE_X96Y95_CO5;
  assign CLBLM_L_X64Y95_SLICE_X97Y95_A = CLBLM_L_X64Y95_SLICE_X97Y95_AO6;
  assign CLBLM_L_X64Y95_SLICE_X97Y95_B = CLBLM_L_X64Y95_SLICE_X97Y95_BO6;
  assign CLBLM_L_X64Y95_SLICE_X97Y95_C = CLBLM_L_X64Y95_SLICE_X97Y95_CO6;
  assign CLBLM_L_X64Y95_SLICE_X97Y95_D = CLBLM_L_X64Y95_SLICE_X97Y95_DO6;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_A = CLBLM_L_X64Y96_SLICE_X96Y96_AO6;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_B = CLBLM_L_X64Y96_SLICE_X96Y96_BO6;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_C = CLBLM_L_X64Y96_SLICE_X96Y96_CO6;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_D = CLBLM_L_X64Y96_SLICE_X96Y96_DO6;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_AMUX = CLBLM_L_X64Y96_SLICE_X96Y96_AO5;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_BMUX = CLBLM_L_X64Y96_SLICE_X96Y96_BO5;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_CMUX = CLBLM_L_X64Y96_SLICE_X96Y96_CO5;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_A = CLBLM_L_X64Y96_SLICE_X97Y96_AO6;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_B = CLBLM_L_X64Y96_SLICE_X97Y96_BO6;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_C = CLBLM_L_X64Y96_SLICE_X97Y96_CO6;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_D = CLBLM_L_X64Y96_SLICE_X97Y96_DO6;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_A = CLBLM_L_X64Y97_SLICE_X96Y97_AO6;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_B = CLBLM_L_X64Y97_SLICE_X96Y97_BO6;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_C = CLBLM_L_X64Y97_SLICE_X96Y97_CO6;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_D = CLBLM_L_X64Y97_SLICE_X96Y97_DO6;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_AMUX = CLBLM_L_X64Y97_SLICE_X96Y97_A5Q;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_BMUX = CLBLM_L_X64Y97_SLICE_X96Y97_B5Q;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_A = CLBLM_L_X64Y97_SLICE_X97Y97_AO6;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_B = CLBLM_L_X64Y97_SLICE_X97Y97_BO6;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_C = CLBLM_L_X64Y97_SLICE_X97Y97_CO6;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_D = CLBLM_L_X64Y97_SLICE_X97Y97_DO6;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_CMUX = CLBLM_L_X64Y97_SLICE_X97Y97_CO6;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_A = CLBLM_L_X64Y98_SLICE_X96Y98_AO6;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_B = CLBLM_L_X64Y98_SLICE_X96Y98_BO6;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_C = CLBLM_L_X64Y98_SLICE_X96Y98_CO6;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_D = CLBLM_L_X64Y98_SLICE_X96Y98_DO6;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_A = CLBLM_L_X64Y98_SLICE_X97Y98_AO6;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_B = CLBLM_L_X64Y98_SLICE_X97Y98_BO6;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_C = CLBLM_L_X64Y98_SLICE_X97Y98_CO6;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_D = CLBLM_L_X64Y98_SLICE_X97Y98_DO6;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_A = CLBLM_L_X64Y99_SLICE_X96Y99_AO6;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_B = CLBLM_L_X64Y99_SLICE_X96Y99_BO6;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_C = CLBLM_L_X64Y99_SLICE_X96Y99_CO6;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_D = CLBLM_L_X64Y99_SLICE_X96Y99_DO6;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_A = CLBLM_L_X64Y99_SLICE_X97Y99_AO6;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_B = CLBLM_L_X64Y99_SLICE_X97Y99_BO6;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_C = CLBLM_L_X64Y99_SLICE_X97Y99_CO6;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_D = CLBLM_L_X64Y99_SLICE_X97Y99_DO6;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_A = CLBLM_L_X64Y100_SLICE_X96Y100_AO6;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_B = CLBLM_L_X64Y100_SLICE_X96Y100_BO6;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_C = CLBLM_L_X64Y100_SLICE_X96Y100_CO6;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_D = CLBLM_L_X64Y100_SLICE_X96Y100_DO6;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_AMUX = CLBLM_L_X64Y100_SLICE_X96Y100_A_XOR;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_BMUX = CLBLM_L_X64Y100_SLICE_X96Y100_B_XOR;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_CMUX = CLBLM_L_X64Y100_SLICE_X96Y100_C_XOR;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_DMUX = CLBLM_L_X64Y100_SLICE_X96Y100_D_XOR;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_A = CLBLM_L_X64Y100_SLICE_X97Y100_AO6;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_B = CLBLM_L_X64Y100_SLICE_X97Y100_BO6;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_C = CLBLM_L_X64Y100_SLICE_X97Y100_CO6;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_D = CLBLM_L_X64Y100_SLICE_X97Y100_DO6;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_AMUX = CLBLM_L_X64Y100_SLICE_X97Y100_A_XOR;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_BMUX = CLBLM_L_X64Y100_SLICE_X97Y100_B_XOR;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_CMUX = CLBLM_L_X64Y100_SLICE_X97Y100_C_XOR;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_DMUX = CLBLM_L_X64Y100_SLICE_X97Y100_D_XOR;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_A = CLBLM_L_X64Y101_SLICE_X96Y101_AO6;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_B = CLBLM_L_X64Y101_SLICE_X96Y101_BO6;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_C = CLBLM_L_X64Y101_SLICE_X96Y101_CO6;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_D = CLBLM_L_X64Y101_SLICE_X96Y101_DO6;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_AMUX = CLBLM_L_X64Y101_SLICE_X96Y101_A_XOR;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_BMUX = CLBLM_L_X64Y101_SLICE_X96Y101_B_XOR;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_CMUX = CLBLM_L_X64Y101_SLICE_X96Y101_C_XOR;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_DMUX = CLBLM_L_X64Y101_SLICE_X96Y101_D_XOR;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_A = CLBLM_L_X64Y101_SLICE_X97Y101_AO6;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_B = CLBLM_L_X64Y101_SLICE_X97Y101_BO6;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_C = CLBLM_L_X64Y101_SLICE_X97Y101_CO6;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_D = CLBLM_L_X64Y101_SLICE_X97Y101_DO6;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_AMUX = CLBLM_L_X64Y101_SLICE_X97Y101_A_XOR;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_BMUX = CLBLM_L_X64Y101_SLICE_X97Y101_B_XOR;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_CMUX = CLBLM_L_X64Y101_SLICE_X97Y101_C_XOR;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_DMUX = CLBLM_L_X64Y101_SLICE_X97Y101_D_XOR;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_A = CLBLM_L_X64Y102_SLICE_X96Y102_AO6;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_B = CLBLM_L_X64Y102_SLICE_X96Y102_BO6;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_C = CLBLM_L_X64Y102_SLICE_X96Y102_CO6;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_D = CLBLM_L_X64Y102_SLICE_X96Y102_DO6;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_AMUX = CLBLM_L_X64Y102_SLICE_X96Y102_A_XOR;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_BMUX = CLBLM_L_X64Y102_SLICE_X96Y102_B_XOR;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_CMUX = CLBLM_L_X64Y102_SLICE_X96Y102_C_XOR;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_DMUX = CLBLM_L_X64Y102_SLICE_X96Y102_D_XOR;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_A = CLBLM_L_X64Y102_SLICE_X97Y102_AO6;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_B = CLBLM_L_X64Y102_SLICE_X97Y102_BO6;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_C = CLBLM_L_X64Y102_SLICE_X97Y102_CO6;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_D = CLBLM_L_X64Y102_SLICE_X97Y102_DO6;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_AMUX = CLBLM_L_X64Y102_SLICE_X97Y102_A_XOR;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_BMUX = CLBLM_L_X64Y102_SLICE_X97Y102_B_XOR;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_CMUX = CLBLM_L_X64Y102_SLICE_X97Y102_C_XOR;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_DMUX = CLBLM_L_X64Y102_SLICE_X97Y102_D_XOR;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_A = CLBLM_L_X64Y103_SLICE_X96Y103_AO6;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_B = CLBLM_L_X64Y103_SLICE_X96Y103_BO6;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_C = CLBLM_L_X64Y103_SLICE_X96Y103_CO6;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_D = CLBLM_L_X64Y103_SLICE_X96Y103_DO6;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_AMUX = CLBLM_L_X64Y103_SLICE_X96Y103_A_XOR;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_BMUX = CLBLM_L_X64Y103_SLICE_X96Y103_B_XOR;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_CMUX = CLBLM_L_X64Y103_SLICE_X96Y103_C_XOR;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_DMUX = CLBLM_L_X64Y103_SLICE_X96Y103_D_XOR;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_A = CLBLM_L_X64Y103_SLICE_X97Y103_AO6;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_B = CLBLM_L_X64Y103_SLICE_X97Y103_BO6;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_C = CLBLM_L_X64Y103_SLICE_X97Y103_CO6;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_D = CLBLM_L_X64Y103_SLICE_X97Y103_DO6;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_AMUX = CLBLM_L_X64Y103_SLICE_X97Y103_A_XOR;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_BMUX = CLBLM_L_X64Y103_SLICE_X97Y103_B_XOR;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_CMUX = CLBLM_L_X64Y103_SLICE_X97Y103_C_XOR;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_DMUX = CLBLM_L_X64Y103_SLICE_X97Y103_D_XOR;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_A = CLBLM_L_X64Y104_SLICE_X96Y104_AO6;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_B = CLBLM_L_X64Y104_SLICE_X96Y104_BO6;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_C = CLBLM_L_X64Y104_SLICE_X96Y104_CO6;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_D = CLBLM_L_X64Y104_SLICE_X96Y104_DO6;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_AMUX = CLBLM_L_X64Y104_SLICE_X96Y104_A_XOR;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_BMUX = CLBLM_L_X64Y104_SLICE_X96Y104_B_XOR;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_A = CLBLM_L_X64Y104_SLICE_X97Y104_AO6;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_B = CLBLM_L_X64Y104_SLICE_X97Y104_BO6;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_C = CLBLM_L_X64Y104_SLICE_X97Y104_CO6;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_D = CLBLM_L_X64Y104_SLICE_X97Y104_DO6;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_AMUX = CLBLM_L_X64Y104_SLICE_X97Y104_A_XOR;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_BMUX = CLBLM_L_X64Y104_SLICE_X97Y104_B_XOR;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_CMUX = CLBLM_L_X64Y104_SLICE_X97Y104_C_XOR;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_A = CLBLM_L_X64Y105_SLICE_X96Y105_AO6;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_B = CLBLM_L_X64Y105_SLICE_X96Y105_BO6;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_C = CLBLM_L_X64Y105_SLICE_X96Y105_CO6;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_D = CLBLM_L_X64Y105_SLICE_X96Y105_DO6;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_A = CLBLM_L_X64Y105_SLICE_X97Y105_AO6;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_B = CLBLM_L_X64Y105_SLICE_X97Y105_BO6;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_C = CLBLM_L_X64Y105_SLICE_X97Y105_CO6;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_D = CLBLM_L_X64Y105_SLICE_X97Y105_DO6;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_DMUX = CLBLM_L_X64Y105_SLICE_X97Y105_DO6;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_A = CLBLM_L_X64Y106_SLICE_X96Y106_AO6;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_B = CLBLM_L_X64Y106_SLICE_X96Y106_BO6;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_C = CLBLM_L_X64Y106_SLICE_X96Y106_CO6;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_D = CLBLM_L_X64Y106_SLICE_X96Y106_DO6;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_DMUX = CLBLM_L_X64Y106_SLICE_X96Y106_DO6;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_A = CLBLM_L_X64Y106_SLICE_X97Y106_AO6;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_B = CLBLM_L_X64Y106_SLICE_X97Y106_BO6;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_C = CLBLM_L_X64Y106_SLICE_X97Y106_CO6;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_D = CLBLM_L_X64Y106_SLICE_X97Y106_DO6;
  assign CLBLM_L_X64Y107_SLICE_X96Y107_A = CLBLM_L_X64Y107_SLICE_X96Y107_AO6;
  assign CLBLM_L_X64Y107_SLICE_X96Y107_B = CLBLM_L_X64Y107_SLICE_X96Y107_BO6;
  assign CLBLM_L_X64Y107_SLICE_X96Y107_C = CLBLM_L_X64Y107_SLICE_X96Y107_CO6;
  assign CLBLM_L_X64Y107_SLICE_X96Y107_D = CLBLM_L_X64Y107_SLICE_X96Y107_DO6;
  assign CLBLM_L_X64Y107_SLICE_X97Y107_A = CLBLM_L_X64Y107_SLICE_X97Y107_AO6;
  assign CLBLM_L_X64Y107_SLICE_X97Y107_B = CLBLM_L_X64Y107_SLICE_X97Y107_BO6;
  assign CLBLM_L_X64Y107_SLICE_X97Y107_C = CLBLM_L_X64Y107_SLICE_X97Y107_CO6;
  assign CLBLM_L_X64Y107_SLICE_X97Y107_D = CLBLM_L_X64Y107_SLICE_X97Y107_DO6;
  assign CLBLM_L_X64Y107_SLICE_X97Y107_DMUX = CLBLM_L_X64Y107_SLICE_X97Y107_DO6;
  assign CLBLM_L_X64Y108_SLICE_X96Y108_A = CLBLM_L_X64Y108_SLICE_X96Y108_AO6;
  assign CLBLM_L_X64Y108_SLICE_X96Y108_B = CLBLM_L_X64Y108_SLICE_X96Y108_BO6;
  assign CLBLM_L_X64Y108_SLICE_X96Y108_C = CLBLM_L_X64Y108_SLICE_X96Y108_CO6;
  assign CLBLM_L_X64Y108_SLICE_X96Y108_D = CLBLM_L_X64Y108_SLICE_X96Y108_DO6;
  assign CLBLM_L_X64Y108_SLICE_X97Y108_A = CLBLM_L_X64Y108_SLICE_X97Y108_AO6;
  assign CLBLM_L_X64Y108_SLICE_X97Y108_B = CLBLM_L_X64Y108_SLICE_X97Y108_BO6;
  assign CLBLM_L_X64Y108_SLICE_X97Y108_C = CLBLM_L_X64Y108_SLICE_X97Y108_CO6;
  assign CLBLM_L_X64Y108_SLICE_X97Y108_D = CLBLM_L_X64Y108_SLICE_X97Y108_DO6;
  assign CLBLM_L_X64Y109_SLICE_X96Y109_A = CLBLM_L_X64Y109_SLICE_X96Y109_AO6;
  assign CLBLM_L_X64Y109_SLICE_X96Y109_B = CLBLM_L_X64Y109_SLICE_X96Y109_BO6;
  assign CLBLM_L_X64Y109_SLICE_X96Y109_C = CLBLM_L_X64Y109_SLICE_X96Y109_CO6;
  assign CLBLM_L_X64Y109_SLICE_X96Y109_D = CLBLM_L_X64Y109_SLICE_X96Y109_DO6;
  assign CLBLM_L_X64Y109_SLICE_X96Y109_AMUX = CLBLM_L_X64Y109_SLICE_X96Y109_A5Q;
  assign CLBLM_L_X64Y109_SLICE_X97Y109_A = CLBLM_L_X64Y109_SLICE_X97Y109_AO6;
  assign CLBLM_L_X64Y109_SLICE_X97Y109_B = CLBLM_L_X64Y109_SLICE_X97Y109_BO6;
  assign CLBLM_L_X64Y109_SLICE_X97Y109_C = CLBLM_L_X64Y109_SLICE_X97Y109_CO6;
  assign CLBLM_L_X64Y109_SLICE_X97Y109_D = CLBLM_L_X64Y109_SLICE_X97Y109_DO6;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_A = CLBLM_R_X15Y122_SLICE_X20Y122_AO6;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_B = CLBLM_R_X15Y122_SLICE_X20Y122_BO6;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_C = CLBLM_R_X15Y122_SLICE_X20Y122_CO6;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_D = CLBLM_R_X15Y122_SLICE_X20Y122_DO6;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_A = CLBLM_R_X15Y122_SLICE_X21Y122_AO6;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_B = CLBLM_R_X15Y122_SLICE_X21Y122_BO6;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_C = CLBLM_R_X15Y122_SLICE_X21Y122_CO6;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_D = CLBLM_R_X15Y122_SLICE_X21Y122_DO6;
  assign CLBLM_R_X47Y119_SLICE_X72Y119_A = CLBLM_R_X47Y119_SLICE_X72Y119_AO6;
  assign CLBLM_R_X47Y119_SLICE_X72Y119_B = CLBLM_R_X47Y119_SLICE_X72Y119_BO6;
  assign CLBLM_R_X47Y119_SLICE_X72Y119_C = CLBLM_R_X47Y119_SLICE_X72Y119_CO6;
  assign CLBLM_R_X47Y119_SLICE_X72Y119_D = CLBLM_R_X47Y119_SLICE_X72Y119_DO6;
  assign CLBLM_R_X47Y119_SLICE_X73Y119_A = CLBLM_R_X47Y119_SLICE_X73Y119_AO6;
  assign CLBLM_R_X47Y119_SLICE_X73Y119_B = CLBLM_R_X47Y119_SLICE_X73Y119_BO6;
  assign CLBLM_R_X47Y119_SLICE_X73Y119_C = CLBLM_R_X47Y119_SLICE_X73Y119_CO6;
  assign CLBLM_R_X47Y119_SLICE_X73Y119_D = CLBLM_R_X47Y119_SLICE_X73Y119_DO6;
  assign CLBLM_R_X47Y119_SLICE_X73Y119_AMUX = CLBLM_R_X47Y119_SLICE_X73Y119_AO5;
  assign CLBLM_R_X49Y104_SLICE_X74Y104_A = CLBLM_R_X49Y104_SLICE_X74Y104_AO6;
  assign CLBLM_R_X49Y104_SLICE_X74Y104_B = CLBLM_R_X49Y104_SLICE_X74Y104_BO6;
  assign CLBLM_R_X49Y104_SLICE_X74Y104_C = CLBLM_R_X49Y104_SLICE_X74Y104_CO6;
  assign CLBLM_R_X49Y104_SLICE_X74Y104_D = CLBLM_R_X49Y104_SLICE_X74Y104_DO6;
  assign CLBLM_R_X49Y104_SLICE_X75Y104_A = CLBLM_R_X49Y104_SLICE_X75Y104_AO6;
  assign CLBLM_R_X49Y104_SLICE_X75Y104_B = CLBLM_R_X49Y104_SLICE_X75Y104_BO6;
  assign CLBLM_R_X49Y104_SLICE_X75Y104_C = CLBLM_R_X49Y104_SLICE_X75Y104_CO6;
  assign CLBLM_R_X49Y104_SLICE_X75Y104_D = CLBLM_R_X49Y104_SLICE_X75Y104_DO6;
  assign CLBLM_R_X49Y105_SLICE_X74Y105_A = CLBLM_R_X49Y105_SLICE_X74Y105_AO6;
  assign CLBLM_R_X49Y105_SLICE_X74Y105_B = CLBLM_R_X49Y105_SLICE_X74Y105_BO6;
  assign CLBLM_R_X49Y105_SLICE_X74Y105_C = CLBLM_R_X49Y105_SLICE_X74Y105_CO6;
  assign CLBLM_R_X49Y105_SLICE_X74Y105_D = CLBLM_R_X49Y105_SLICE_X74Y105_DO6;
  assign CLBLM_R_X49Y105_SLICE_X75Y105_A = CLBLM_R_X49Y105_SLICE_X75Y105_AO6;
  assign CLBLM_R_X49Y105_SLICE_X75Y105_B = CLBLM_R_X49Y105_SLICE_X75Y105_BO6;
  assign CLBLM_R_X49Y105_SLICE_X75Y105_C = CLBLM_R_X49Y105_SLICE_X75Y105_CO6;
  assign CLBLM_R_X49Y105_SLICE_X75Y105_D = CLBLM_R_X49Y105_SLICE_X75Y105_DO6;
  assign CLBLM_R_X49Y105_SLICE_X75Y105_AMUX = CLBLM_R_X49Y105_SLICE_X75Y105_F7AMUX_O;
  assign CLBLM_R_X49Y106_SLICE_X74Y106_A = CLBLM_R_X49Y106_SLICE_X74Y106_AO6;
  assign CLBLM_R_X49Y106_SLICE_X74Y106_B = CLBLM_R_X49Y106_SLICE_X74Y106_BO6;
  assign CLBLM_R_X49Y106_SLICE_X74Y106_C = CLBLM_R_X49Y106_SLICE_X74Y106_CO6;
  assign CLBLM_R_X49Y106_SLICE_X74Y106_D = CLBLM_R_X49Y106_SLICE_X74Y106_DO6;
  assign CLBLM_R_X49Y106_SLICE_X74Y106_CMUX = CLBLM_R_X49Y106_SLICE_X74Y106_CO6;
  assign CLBLM_R_X49Y106_SLICE_X75Y106_A = CLBLM_R_X49Y106_SLICE_X75Y106_AO6;
  assign CLBLM_R_X49Y106_SLICE_X75Y106_B = CLBLM_R_X49Y106_SLICE_X75Y106_BO6;
  assign CLBLM_R_X49Y106_SLICE_X75Y106_C = CLBLM_R_X49Y106_SLICE_X75Y106_CO6;
  assign CLBLM_R_X49Y106_SLICE_X75Y106_D = CLBLM_R_X49Y106_SLICE_X75Y106_DO6;
  assign CLBLM_R_X49Y106_SLICE_X75Y106_AMUX = CLBLM_R_X49Y106_SLICE_X75Y106_F7AMUX_O;
  assign CLBLM_R_X49Y106_SLICE_X75Y106_DMUX = CLBLM_R_X49Y106_SLICE_X75Y106_DO6;
  assign CLBLM_R_X49Y107_SLICE_X74Y107_A = CLBLM_R_X49Y107_SLICE_X74Y107_AO6;
  assign CLBLM_R_X49Y107_SLICE_X74Y107_B = CLBLM_R_X49Y107_SLICE_X74Y107_BO6;
  assign CLBLM_R_X49Y107_SLICE_X74Y107_C = CLBLM_R_X49Y107_SLICE_X74Y107_CO6;
  assign CLBLM_R_X49Y107_SLICE_X74Y107_D = CLBLM_R_X49Y107_SLICE_X74Y107_DO6;
  assign CLBLM_R_X49Y107_SLICE_X75Y107_A = CLBLM_R_X49Y107_SLICE_X75Y107_AO6;
  assign CLBLM_R_X49Y107_SLICE_X75Y107_B = CLBLM_R_X49Y107_SLICE_X75Y107_BO6;
  assign CLBLM_R_X49Y107_SLICE_X75Y107_C = CLBLM_R_X49Y107_SLICE_X75Y107_CO6;
  assign CLBLM_R_X49Y107_SLICE_X75Y107_D = CLBLM_R_X49Y107_SLICE_X75Y107_DO6;
  assign CLBLM_R_X49Y107_SLICE_X75Y107_AMUX = CLBLM_R_X49Y107_SLICE_X75Y107_F7AMUX_O;
  assign CLBLM_R_X49Y107_SLICE_X75Y107_CMUX = CLBLM_R_X49Y107_SLICE_X75Y107_CO5;
  assign CLBLM_R_X49Y108_SLICE_X74Y108_A = CLBLM_R_X49Y108_SLICE_X74Y108_AO6;
  assign CLBLM_R_X49Y108_SLICE_X74Y108_B = CLBLM_R_X49Y108_SLICE_X74Y108_BO6;
  assign CLBLM_R_X49Y108_SLICE_X74Y108_C = CLBLM_R_X49Y108_SLICE_X74Y108_CO6;
  assign CLBLM_R_X49Y108_SLICE_X74Y108_D = CLBLM_R_X49Y108_SLICE_X74Y108_DO6;
  assign CLBLM_R_X49Y108_SLICE_X74Y108_AMUX = CLBLM_R_X49Y108_SLICE_X74Y108_A5Q;
  assign CLBLM_R_X49Y108_SLICE_X74Y108_BMUX = CLBLM_R_X49Y108_SLICE_X74Y108_B5Q;
  assign CLBLM_R_X49Y108_SLICE_X74Y108_CMUX = CLBLM_R_X49Y108_SLICE_X74Y108_C5Q;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_A = CLBLM_R_X49Y108_SLICE_X75Y108_AO6;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_B = CLBLM_R_X49Y108_SLICE_X75Y108_BO6;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_C = CLBLM_R_X49Y108_SLICE_X75Y108_CO6;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_D = CLBLM_R_X49Y108_SLICE_X75Y108_DO6;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_AMUX = CLBLM_R_X49Y108_SLICE_X75Y108_A_XOR;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_BMUX = CLBLM_R_X49Y108_SLICE_X75Y108_B_XOR;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_CMUX = CLBLM_R_X49Y108_SLICE_X75Y108_C_XOR;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_DMUX = CLBLM_R_X49Y108_SLICE_X75Y108_D_XOR;
  assign CLBLM_R_X49Y109_SLICE_X74Y109_A = CLBLM_R_X49Y109_SLICE_X74Y109_AO6;
  assign CLBLM_R_X49Y109_SLICE_X74Y109_B = CLBLM_R_X49Y109_SLICE_X74Y109_BO6;
  assign CLBLM_R_X49Y109_SLICE_X74Y109_C = CLBLM_R_X49Y109_SLICE_X74Y109_CO6;
  assign CLBLM_R_X49Y109_SLICE_X74Y109_D = CLBLM_R_X49Y109_SLICE_X74Y109_DO6;
  assign CLBLM_R_X49Y109_SLICE_X75Y109_A = CLBLM_R_X49Y109_SLICE_X75Y109_AO6;
  assign CLBLM_R_X49Y109_SLICE_X75Y109_B = CLBLM_R_X49Y109_SLICE_X75Y109_BO6;
  assign CLBLM_R_X49Y109_SLICE_X75Y109_C = CLBLM_R_X49Y109_SLICE_X75Y109_CO6;
  assign CLBLM_R_X49Y109_SLICE_X75Y109_D = CLBLM_R_X49Y109_SLICE_X75Y109_DO6;
  assign CLBLM_R_X49Y109_SLICE_X75Y109_AMUX = CLBLM_R_X49Y109_SLICE_X75Y109_A_XOR;
  assign CLBLM_R_X49Y109_SLICE_X75Y109_BMUX = CLBLM_R_X49Y109_SLICE_X75Y109_B_XOR;
  assign CLBLM_R_X49Y109_SLICE_X75Y109_CMUX = CLBLM_R_X49Y109_SLICE_X75Y109_C_XOR;
  assign CLBLM_R_X49Y109_SLICE_X75Y109_DMUX = CLBLM_R_X49Y109_SLICE_X75Y109_D_XOR;
  assign CLBLM_R_X49Y110_SLICE_X74Y110_A = CLBLM_R_X49Y110_SLICE_X74Y110_AO6;
  assign CLBLM_R_X49Y110_SLICE_X74Y110_B = CLBLM_R_X49Y110_SLICE_X74Y110_BO6;
  assign CLBLM_R_X49Y110_SLICE_X74Y110_C = CLBLM_R_X49Y110_SLICE_X74Y110_CO6;
  assign CLBLM_R_X49Y110_SLICE_X74Y110_D = CLBLM_R_X49Y110_SLICE_X74Y110_DO6;
  assign CLBLM_R_X49Y110_SLICE_X74Y110_AMUX = CLBLM_R_X49Y110_SLICE_X74Y110_A5Q;
  assign CLBLM_R_X49Y110_SLICE_X75Y110_A = CLBLM_R_X49Y110_SLICE_X75Y110_AO6;
  assign CLBLM_R_X49Y110_SLICE_X75Y110_B = CLBLM_R_X49Y110_SLICE_X75Y110_BO6;
  assign CLBLM_R_X49Y110_SLICE_X75Y110_C = CLBLM_R_X49Y110_SLICE_X75Y110_CO6;
  assign CLBLM_R_X49Y110_SLICE_X75Y110_D = CLBLM_R_X49Y110_SLICE_X75Y110_DO6;
  assign CLBLM_R_X49Y110_SLICE_X75Y110_AMUX = CLBLM_R_X49Y110_SLICE_X75Y110_A_CY;
  assign CLBLM_R_X49Y111_SLICE_X74Y111_A = CLBLM_R_X49Y111_SLICE_X74Y111_AO6;
  assign CLBLM_R_X49Y111_SLICE_X74Y111_B = CLBLM_R_X49Y111_SLICE_X74Y111_BO6;
  assign CLBLM_R_X49Y111_SLICE_X74Y111_C = CLBLM_R_X49Y111_SLICE_X74Y111_CO6;
  assign CLBLM_R_X49Y111_SLICE_X74Y111_D = CLBLM_R_X49Y111_SLICE_X74Y111_DO6;
  assign CLBLM_R_X49Y111_SLICE_X75Y111_A = CLBLM_R_X49Y111_SLICE_X75Y111_AO6;
  assign CLBLM_R_X49Y111_SLICE_X75Y111_B = CLBLM_R_X49Y111_SLICE_X75Y111_BO6;
  assign CLBLM_R_X49Y111_SLICE_X75Y111_C = CLBLM_R_X49Y111_SLICE_X75Y111_CO6;
  assign CLBLM_R_X49Y111_SLICE_X75Y111_D = CLBLM_R_X49Y111_SLICE_X75Y111_DO6;
  assign CLBLM_R_X49Y111_SLICE_X75Y111_AMUX = CLBLM_R_X49Y111_SLICE_X75Y111_A5Q;
  assign CLBLM_R_X49Y111_SLICE_X75Y111_BMUX = CLBLM_R_X49Y111_SLICE_X75Y111_BO6;
  assign CLBLM_R_X49Y119_SLICE_X74Y119_A = CLBLM_R_X49Y119_SLICE_X74Y119_AO6;
  assign CLBLM_R_X49Y119_SLICE_X74Y119_B = CLBLM_R_X49Y119_SLICE_X74Y119_BO6;
  assign CLBLM_R_X49Y119_SLICE_X74Y119_C = CLBLM_R_X49Y119_SLICE_X74Y119_CO6;
  assign CLBLM_R_X49Y119_SLICE_X74Y119_D = CLBLM_R_X49Y119_SLICE_X74Y119_DO6;
  assign CLBLM_R_X49Y119_SLICE_X75Y119_A = CLBLM_R_X49Y119_SLICE_X75Y119_AO6;
  assign CLBLM_R_X49Y119_SLICE_X75Y119_B = CLBLM_R_X49Y119_SLICE_X75Y119_BO6;
  assign CLBLM_R_X49Y119_SLICE_X75Y119_C = CLBLM_R_X49Y119_SLICE_X75Y119_CO6;
  assign CLBLM_R_X49Y119_SLICE_X75Y119_D = CLBLM_R_X49Y119_SLICE_X75Y119_DO6;
  assign CLBLM_R_X53Y98_SLICE_X80Y98_A = CLBLM_R_X53Y98_SLICE_X80Y98_AO6;
  assign CLBLM_R_X53Y98_SLICE_X80Y98_B = CLBLM_R_X53Y98_SLICE_X80Y98_BO6;
  assign CLBLM_R_X53Y98_SLICE_X80Y98_C = CLBLM_R_X53Y98_SLICE_X80Y98_CO6;
  assign CLBLM_R_X53Y98_SLICE_X80Y98_D = CLBLM_R_X53Y98_SLICE_X80Y98_DO6;
  assign CLBLM_R_X53Y98_SLICE_X81Y98_A = CLBLM_R_X53Y98_SLICE_X81Y98_AO6;
  assign CLBLM_R_X53Y98_SLICE_X81Y98_B = CLBLM_R_X53Y98_SLICE_X81Y98_BO6;
  assign CLBLM_R_X53Y98_SLICE_X81Y98_C = CLBLM_R_X53Y98_SLICE_X81Y98_CO6;
  assign CLBLM_R_X53Y98_SLICE_X81Y98_D = CLBLM_R_X53Y98_SLICE_X81Y98_DO6;
  assign CLBLM_R_X53Y99_SLICE_X80Y99_A = CLBLM_R_X53Y99_SLICE_X80Y99_AO6;
  assign CLBLM_R_X53Y99_SLICE_X80Y99_B = CLBLM_R_X53Y99_SLICE_X80Y99_BO6;
  assign CLBLM_R_X53Y99_SLICE_X80Y99_C = CLBLM_R_X53Y99_SLICE_X80Y99_CO6;
  assign CLBLM_R_X53Y99_SLICE_X80Y99_D = CLBLM_R_X53Y99_SLICE_X80Y99_DO6;
  assign CLBLM_R_X53Y99_SLICE_X80Y99_AMUX = CLBLM_R_X53Y99_SLICE_X80Y99_AO5;
  assign CLBLM_R_X53Y99_SLICE_X80Y99_BMUX = CLBLM_R_X53Y99_SLICE_X80Y99_BO5;
  assign CLBLM_R_X53Y99_SLICE_X80Y99_DMUX = CLBLM_R_X53Y99_SLICE_X80Y99_DO6;
  assign CLBLM_R_X53Y99_SLICE_X81Y99_A = CLBLM_R_X53Y99_SLICE_X81Y99_AO6;
  assign CLBLM_R_X53Y99_SLICE_X81Y99_B = CLBLM_R_X53Y99_SLICE_X81Y99_BO6;
  assign CLBLM_R_X53Y99_SLICE_X81Y99_C = CLBLM_R_X53Y99_SLICE_X81Y99_CO6;
  assign CLBLM_R_X53Y99_SLICE_X81Y99_D = CLBLM_R_X53Y99_SLICE_X81Y99_DO6;
  assign CLBLM_R_X53Y99_SLICE_X81Y99_AMUX = CLBLM_R_X53Y99_SLICE_X81Y99_AO5;
  assign CLBLM_R_X53Y100_SLICE_X80Y100_A = CLBLM_R_X53Y100_SLICE_X80Y100_AO6;
  assign CLBLM_R_X53Y100_SLICE_X80Y100_B = CLBLM_R_X53Y100_SLICE_X80Y100_BO6;
  assign CLBLM_R_X53Y100_SLICE_X80Y100_C = CLBLM_R_X53Y100_SLICE_X80Y100_CO6;
  assign CLBLM_R_X53Y100_SLICE_X80Y100_D = CLBLM_R_X53Y100_SLICE_X80Y100_DO6;
  assign CLBLM_R_X53Y100_SLICE_X80Y100_AMUX = CLBLM_R_X53Y100_SLICE_X80Y100_A5Q;
  assign CLBLM_R_X53Y100_SLICE_X80Y100_BMUX = CLBLM_R_X53Y100_SLICE_X80Y100_BO5;
  assign CLBLM_R_X53Y100_SLICE_X80Y100_CMUX = CLBLM_R_X53Y100_SLICE_X80Y100_CO6;
  assign CLBLM_R_X53Y100_SLICE_X81Y100_A = CLBLM_R_X53Y100_SLICE_X81Y100_AO6;
  assign CLBLM_R_X53Y100_SLICE_X81Y100_B = CLBLM_R_X53Y100_SLICE_X81Y100_BO6;
  assign CLBLM_R_X53Y100_SLICE_X81Y100_C = CLBLM_R_X53Y100_SLICE_X81Y100_CO6;
  assign CLBLM_R_X53Y100_SLICE_X81Y100_D = CLBLM_R_X53Y100_SLICE_X81Y100_DO6;
  assign CLBLM_R_X53Y100_SLICE_X81Y100_AMUX = CLBLM_R_X53Y100_SLICE_X81Y100_AO5;
  assign CLBLM_R_X53Y101_SLICE_X80Y101_A = CLBLM_R_X53Y101_SLICE_X80Y101_AO6;
  assign CLBLM_R_X53Y101_SLICE_X80Y101_B = CLBLM_R_X53Y101_SLICE_X80Y101_BO6;
  assign CLBLM_R_X53Y101_SLICE_X80Y101_C = CLBLM_R_X53Y101_SLICE_X80Y101_CO6;
  assign CLBLM_R_X53Y101_SLICE_X80Y101_D = CLBLM_R_X53Y101_SLICE_X80Y101_DO6;
  assign CLBLM_R_X53Y101_SLICE_X80Y101_AMUX = CLBLM_R_X53Y101_SLICE_X80Y101_AO5;
  assign CLBLM_R_X53Y101_SLICE_X81Y101_A = CLBLM_R_X53Y101_SLICE_X81Y101_AO6;
  assign CLBLM_R_X53Y101_SLICE_X81Y101_B = CLBLM_R_X53Y101_SLICE_X81Y101_BO6;
  assign CLBLM_R_X53Y101_SLICE_X81Y101_C = CLBLM_R_X53Y101_SLICE_X81Y101_CO6;
  assign CLBLM_R_X53Y101_SLICE_X81Y101_D = CLBLM_R_X53Y101_SLICE_X81Y101_DO6;
  assign CLBLM_R_X53Y101_SLICE_X81Y101_BMUX = CLBLM_R_X53Y101_SLICE_X81Y101_BO6;
  assign CLBLM_R_X53Y102_SLICE_X80Y102_A = CLBLM_R_X53Y102_SLICE_X80Y102_AO6;
  assign CLBLM_R_X53Y102_SLICE_X80Y102_B = CLBLM_R_X53Y102_SLICE_X80Y102_BO6;
  assign CLBLM_R_X53Y102_SLICE_X80Y102_C = CLBLM_R_X53Y102_SLICE_X80Y102_CO6;
  assign CLBLM_R_X53Y102_SLICE_X80Y102_D = CLBLM_R_X53Y102_SLICE_X80Y102_DO6;
  assign CLBLM_R_X53Y102_SLICE_X81Y102_A = CLBLM_R_X53Y102_SLICE_X81Y102_AO6;
  assign CLBLM_R_X53Y102_SLICE_X81Y102_B = CLBLM_R_X53Y102_SLICE_X81Y102_BO6;
  assign CLBLM_R_X53Y102_SLICE_X81Y102_C = CLBLM_R_X53Y102_SLICE_X81Y102_CO6;
  assign CLBLM_R_X53Y102_SLICE_X81Y102_D = CLBLM_R_X53Y102_SLICE_X81Y102_DO6;
  assign CLBLM_R_X53Y103_SLICE_X80Y103_A = CLBLM_R_X53Y103_SLICE_X80Y103_AO6;
  assign CLBLM_R_X53Y103_SLICE_X80Y103_B = CLBLM_R_X53Y103_SLICE_X80Y103_BO6;
  assign CLBLM_R_X53Y103_SLICE_X80Y103_C = CLBLM_R_X53Y103_SLICE_X80Y103_CO6;
  assign CLBLM_R_X53Y103_SLICE_X80Y103_D = CLBLM_R_X53Y103_SLICE_X80Y103_DO6;
  assign CLBLM_R_X53Y103_SLICE_X81Y103_A = CLBLM_R_X53Y103_SLICE_X81Y103_AO6;
  assign CLBLM_R_X53Y103_SLICE_X81Y103_B = CLBLM_R_X53Y103_SLICE_X81Y103_BO6;
  assign CLBLM_R_X53Y103_SLICE_X81Y103_C = CLBLM_R_X53Y103_SLICE_X81Y103_CO6;
  assign CLBLM_R_X53Y103_SLICE_X81Y103_D = CLBLM_R_X53Y103_SLICE_X81Y103_DO6;
  assign CLBLM_R_X53Y103_SLICE_X81Y103_AMUX = CLBLM_R_X53Y103_SLICE_X81Y103_A_XOR;
  assign CLBLM_R_X53Y103_SLICE_X81Y103_BMUX = CLBLM_R_X53Y103_SLICE_X81Y103_B_XOR;
  assign CLBLM_R_X53Y103_SLICE_X81Y103_CMUX = CLBLM_R_X53Y103_SLICE_X81Y103_C_XOR;
  assign CLBLM_R_X53Y103_SLICE_X81Y103_DMUX = CLBLM_R_X53Y103_SLICE_X81Y103_D_XOR;
  assign CLBLM_R_X53Y104_SLICE_X80Y104_A = CLBLM_R_X53Y104_SLICE_X80Y104_AO6;
  assign CLBLM_R_X53Y104_SLICE_X80Y104_B = CLBLM_R_X53Y104_SLICE_X80Y104_BO6;
  assign CLBLM_R_X53Y104_SLICE_X80Y104_C = CLBLM_R_X53Y104_SLICE_X80Y104_CO6;
  assign CLBLM_R_X53Y104_SLICE_X80Y104_D = CLBLM_R_X53Y104_SLICE_X80Y104_DO6;
  assign CLBLM_R_X53Y104_SLICE_X80Y104_AMUX = CLBLM_R_X53Y104_SLICE_X80Y104_AO5;
  assign CLBLM_R_X53Y104_SLICE_X80Y104_CMUX = CLBLM_R_X53Y104_SLICE_X80Y104_CO6;
  assign CLBLM_R_X53Y104_SLICE_X80Y104_DMUX = CLBLM_R_X53Y104_SLICE_X80Y104_DO5;
  assign CLBLM_R_X53Y104_SLICE_X81Y104_A = CLBLM_R_X53Y104_SLICE_X81Y104_AO6;
  assign CLBLM_R_X53Y104_SLICE_X81Y104_B = CLBLM_R_X53Y104_SLICE_X81Y104_BO6;
  assign CLBLM_R_X53Y104_SLICE_X81Y104_C = CLBLM_R_X53Y104_SLICE_X81Y104_CO6;
  assign CLBLM_R_X53Y104_SLICE_X81Y104_D = CLBLM_R_X53Y104_SLICE_X81Y104_DO6;
  assign CLBLM_R_X53Y104_SLICE_X81Y104_AMUX = CLBLM_R_X53Y104_SLICE_X81Y104_A_XOR;
  assign CLBLM_R_X53Y104_SLICE_X81Y104_BMUX = CLBLM_R_X53Y104_SLICE_X81Y104_B_XOR;
  assign CLBLM_R_X53Y104_SLICE_X81Y104_CMUX = CLBLM_R_X53Y104_SLICE_X81Y104_C_XOR;
  assign CLBLM_R_X53Y104_SLICE_X81Y104_DMUX = CLBLM_R_X53Y104_SLICE_X81Y104_D_XOR;
  assign CLBLM_R_X53Y105_SLICE_X80Y105_A = CLBLM_R_X53Y105_SLICE_X80Y105_AO6;
  assign CLBLM_R_X53Y105_SLICE_X80Y105_B = CLBLM_R_X53Y105_SLICE_X80Y105_BO6;
  assign CLBLM_R_X53Y105_SLICE_X80Y105_C = CLBLM_R_X53Y105_SLICE_X80Y105_CO6;
  assign CLBLM_R_X53Y105_SLICE_X80Y105_D = CLBLM_R_X53Y105_SLICE_X80Y105_DO6;
  assign CLBLM_R_X53Y105_SLICE_X81Y105_A = CLBLM_R_X53Y105_SLICE_X81Y105_AO6;
  assign CLBLM_R_X53Y105_SLICE_X81Y105_B = CLBLM_R_X53Y105_SLICE_X81Y105_BO6;
  assign CLBLM_R_X53Y105_SLICE_X81Y105_C = CLBLM_R_X53Y105_SLICE_X81Y105_CO6;
  assign CLBLM_R_X53Y105_SLICE_X81Y105_D = CLBLM_R_X53Y105_SLICE_X81Y105_DO6;
  assign CLBLM_R_X53Y105_SLICE_X81Y105_AMUX = CLBLM_R_X53Y105_SLICE_X81Y105_A_XOR;
  assign CLBLM_R_X53Y105_SLICE_X81Y105_BMUX = CLBLM_R_X53Y105_SLICE_X81Y105_B_XOR;
  assign CLBLM_R_X53Y105_SLICE_X81Y105_CMUX = CLBLM_R_X53Y105_SLICE_X81Y105_C_CY;
  assign CLBLM_R_X53Y106_SLICE_X80Y106_A = CLBLM_R_X53Y106_SLICE_X80Y106_AO6;
  assign CLBLM_R_X53Y106_SLICE_X80Y106_B = CLBLM_R_X53Y106_SLICE_X80Y106_BO6;
  assign CLBLM_R_X53Y106_SLICE_X80Y106_C = CLBLM_R_X53Y106_SLICE_X80Y106_CO6;
  assign CLBLM_R_X53Y106_SLICE_X80Y106_D = CLBLM_R_X53Y106_SLICE_X80Y106_DO6;
  assign CLBLM_R_X53Y106_SLICE_X80Y106_AMUX = CLBLM_R_X53Y106_SLICE_X80Y106_AO5;
  assign CLBLM_R_X53Y106_SLICE_X81Y106_A = CLBLM_R_X53Y106_SLICE_X81Y106_AO6;
  assign CLBLM_R_X53Y106_SLICE_X81Y106_B = CLBLM_R_X53Y106_SLICE_X81Y106_BO6;
  assign CLBLM_R_X53Y106_SLICE_X81Y106_C = CLBLM_R_X53Y106_SLICE_X81Y106_CO6;
  assign CLBLM_R_X53Y106_SLICE_X81Y106_D = CLBLM_R_X53Y106_SLICE_X81Y106_DO6;
  assign CLBLM_R_X53Y106_SLICE_X81Y106_AMUX = CLBLM_R_X53Y106_SLICE_X81Y106_A_XOR;
  assign CLBLM_R_X53Y106_SLICE_X81Y106_BMUX = CLBLM_R_X53Y106_SLICE_X81Y106_B_XOR;
  assign CLBLM_R_X53Y106_SLICE_X81Y106_CMUX = CLBLM_R_X53Y106_SLICE_X81Y106_C_XOR;
  assign CLBLM_R_X53Y106_SLICE_X81Y106_DMUX = CLBLM_R_X53Y106_SLICE_X81Y106_D_XOR;
  assign CLBLM_R_X53Y107_SLICE_X80Y107_A = CLBLM_R_X53Y107_SLICE_X80Y107_AO6;
  assign CLBLM_R_X53Y107_SLICE_X80Y107_B = CLBLM_R_X53Y107_SLICE_X80Y107_BO6;
  assign CLBLM_R_X53Y107_SLICE_X80Y107_C = CLBLM_R_X53Y107_SLICE_X80Y107_CO6;
  assign CLBLM_R_X53Y107_SLICE_X80Y107_D = CLBLM_R_X53Y107_SLICE_X80Y107_DO6;
  assign CLBLM_R_X53Y107_SLICE_X80Y107_AMUX = CLBLM_R_X53Y107_SLICE_X80Y107_AO5;
  assign CLBLM_R_X53Y107_SLICE_X80Y107_BMUX = CLBLM_R_X53Y107_SLICE_X80Y107_BO5;
  assign CLBLM_R_X53Y107_SLICE_X81Y107_A = CLBLM_R_X53Y107_SLICE_X81Y107_AO6;
  assign CLBLM_R_X53Y107_SLICE_X81Y107_B = CLBLM_R_X53Y107_SLICE_X81Y107_BO6;
  assign CLBLM_R_X53Y107_SLICE_X81Y107_C = CLBLM_R_X53Y107_SLICE_X81Y107_CO6;
  assign CLBLM_R_X53Y107_SLICE_X81Y107_D = CLBLM_R_X53Y107_SLICE_X81Y107_DO6;
  assign CLBLM_R_X53Y107_SLICE_X81Y107_AMUX = CLBLM_R_X53Y107_SLICE_X81Y107_A_XOR;
  assign CLBLM_R_X53Y107_SLICE_X81Y107_BMUX = CLBLM_R_X53Y107_SLICE_X81Y107_B_XOR;
  assign CLBLM_R_X53Y107_SLICE_X81Y107_CMUX = CLBLM_R_X53Y107_SLICE_X81Y107_C_XOR;
  assign CLBLM_R_X53Y107_SLICE_X81Y107_DMUX = CLBLM_R_X53Y107_SLICE_X81Y107_D_XOR;
  assign CLBLM_R_X53Y108_SLICE_X80Y108_A = CLBLM_R_X53Y108_SLICE_X80Y108_AO6;
  assign CLBLM_R_X53Y108_SLICE_X80Y108_B = CLBLM_R_X53Y108_SLICE_X80Y108_BO6;
  assign CLBLM_R_X53Y108_SLICE_X80Y108_C = CLBLM_R_X53Y108_SLICE_X80Y108_CO6;
  assign CLBLM_R_X53Y108_SLICE_X80Y108_D = CLBLM_R_X53Y108_SLICE_X80Y108_DO6;
  assign CLBLM_R_X53Y108_SLICE_X80Y108_CMUX = CLBLM_R_X53Y108_SLICE_X80Y108_CO6;
  assign CLBLM_R_X53Y108_SLICE_X81Y108_A = CLBLM_R_X53Y108_SLICE_X81Y108_AO6;
  assign CLBLM_R_X53Y108_SLICE_X81Y108_B = CLBLM_R_X53Y108_SLICE_X81Y108_BO6;
  assign CLBLM_R_X53Y108_SLICE_X81Y108_C = CLBLM_R_X53Y108_SLICE_X81Y108_CO6;
  assign CLBLM_R_X53Y108_SLICE_X81Y108_D = CLBLM_R_X53Y108_SLICE_X81Y108_DO6;
  assign CLBLM_R_X53Y108_SLICE_X81Y108_AMUX = CLBLM_R_X53Y108_SLICE_X81Y108_A_XOR;
  assign CLBLM_R_X53Y108_SLICE_X81Y108_BMUX = CLBLM_R_X53Y108_SLICE_X81Y108_B_XOR;
  assign CLBLM_R_X53Y108_SLICE_X81Y108_CMUX = CLBLM_R_X53Y108_SLICE_X81Y108_C_CY;
  assign CLBLM_R_X59Y96_SLICE_X88Y96_A = CLBLM_R_X59Y96_SLICE_X88Y96_AO6;
  assign CLBLM_R_X59Y96_SLICE_X88Y96_B = CLBLM_R_X59Y96_SLICE_X88Y96_BO6;
  assign CLBLM_R_X59Y96_SLICE_X88Y96_C = CLBLM_R_X59Y96_SLICE_X88Y96_CO6;
  assign CLBLM_R_X59Y96_SLICE_X88Y96_D = CLBLM_R_X59Y96_SLICE_X88Y96_DO6;
  assign CLBLM_R_X59Y96_SLICE_X88Y96_DMUX = CLBLM_R_X59Y96_SLICE_X88Y96_DO6;
  assign CLBLM_R_X59Y96_SLICE_X89Y96_A = CLBLM_R_X59Y96_SLICE_X89Y96_AO6;
  assign CLBLM_R_X59Y96_SLICE_X89Y96_B = CLBLM_R_X59Y96_SLICE_X89Y96_BO6;
  assign CLBLM_R_X59Y96_SLICE_X89Y96_C = CLBLM_R_X59Y96_SLICE_X89Y96_CO6;
  assign CLBLM_R_X59Y96_SLICE_X89Y96_D = CLBLM_R_X59Y96_SLICE_X89Y96_DO6;
  assign CLBLM_R_X59Y96_SLICE_X89Y96_AMUX = CLBLM_R_X59Y96_SLICE_X89Y96_A5Q;
  assign CLBLM_R_X59Y97_SLICE_X88Y97_A = CLBLM_R_X59Y97_SLICE_X88Y97_AO6;
  assign CLBLM_R_X59Y97_SLICE_X88Y97_B = CLBLM_R_X59Y97_SLICE_X88Y97_BO6;
  assign CLBLM_R_X59Y97_SLICE_X88Y97_C = CLBLM_R_X59Y97_SLICE_X88Y97_CO6;
  assign CLBLM_R_X59Y97_SLICE_X88Y97_D = CLBLM_R_X59Y97_SLICE_X88Y97_DO6;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_A = CLBLM_R_X59Y97_SLICE_X89Y97_AO6;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_B = CLBLM_R_X59Y97_SLICE_X89Y97_BO6;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_C = CLBLM_R_X59Y97_SLICE_X89Y97_CO6;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_D = CLBLM_R_X59Y97_SLICE_X89Y97_DO6;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_AMUX = CLBLM_R_X59Y97_SLICE_X89Y97_A5Q;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_BMUX = CLBLM_R_X59Y97_SLICE_X89Y97_B5Q;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_CMUX = CLBLM_R_X59Y97_SLICE_X89Y97_C5Q;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_DMUX = CLBLM_R_X59Y97_SLICE_X89Y97_D5Q;
  assign CLBLM_R_X59Y98_SLICE_X88Y98_A = CLBLM_R_X59Y98_SLICE_X88Y98_AO6;
  assign CLBLM_R_X59Y98_SLICE_X88Y98_B = CLBLM_R_X59Y98_SLICE_X88Y98_BO6;
  assign CLBLM_R_X59Y98_SLICE_X88Y98_C = CLBLM_R_X59Y98_SLICE_X88Y98_CO6;
  assign CLBLM_R_X59Y98_SLICE_X88Y98_D = CLBLM_R_X59Y98_SLICE_X88Y98_DO6;
  assign CLBLM_R_X59Y98_SLICE_X89Y98_A = CLBLM_R_X59Y98_SLICE_X89Y98_AO6;
  assign CLBLM_R_X59Y98_SLICE_X89Y98_B = CLBLM_R_X59Y98_SLICE_X89Y98_BO6;
  assign CLBLM_R_X59Y98_SLICE_X89Y98_C = CLBLM_R_X59Y98_SLICE_X89Y98_CO6;
  assign CLBLM_R_X59Y98_SLICE_X89Y98_D = CLBLM_R_X59Y98_SLICE_X89Y98_DO6;
  assign CLBLM_R_X59Y98_SLICE_X89Y98_AMUX = CLBLM_R_X59Y98_SLICE_X89Y98_A5Q;
  assign CLBLM_R_X59Y98_SLICE_X89Y98_BMUX = CLBLM_R_X59Y98_SLICE_X89Y98_B5Q;
  assign CLBLM_R_X59Y98_SLICE_X89Y98_CMUX = CLBLM_R_X59Y98_SLICE_X89Y98_C5Q;
  assign CLBLM_R_X59Y98_SLICE_X89Y98_DMUX = CLBLM_R_X59Y98_SLICE_X89Y98_DO6;
  assign CLBLM_R_X59Y99_SLICE_X88Y99_A = CLBLM_R_X59Y99_SLICE_X88Y99_AO6;
  assign CLBLM_R_X59Y99_SLICE_X88Y99_B = CLBLM_R_X59Y99_SLICE_X88Y99_BO6;
  assign CLBLM_R_X59Y99_SLICE_X88Y99_C = CLBLM_R_X59Y99_SLICE_X88Y99_CO6;
  assign CLBLM_R_X59Y99_SLICE_X88Y99_D = CLBLM_R_X59Y99_SLICE_X88Y99_DO6;
  assign CLBLM_R_X59Y99_SLICE_X88Y99_BMUX = CLBLM_R_X59Y99_SLICE_X88Y99_B5Q;
  assign CLBLM_R_X59Y99_SLICE_X89Y99_A = CLBLM_R_X59Y99_SLICE_X89Y99_AO6;
  assign CLBLM_R_X59Y99_SLICE_X89Y99_B = CLBLM_R_X59Y99_SLICE_X89Y99_BO6;
  assign CLBLM_R_X59Y99_SLICE_X89Y99_C = CLBLM_R_X59Y99_SLICE_X89Y99_CO6;
  assign CLBLM_R_X59Y99_SLICE_X89Y99_D = CLBLM_R_X59Y99_SLICE_X89Y99_DO6;
  assign CLBLM_R_X59Y99_SLICE_X89Y99_AMUX = CLBLM_R_X59Y99_SLICE_X89Y99_A5Q;
  assign CLBLM_R_X59Y100_SLICE_X88Y100_A = CLBLM_R_X59Y100_SLICE_X88Y100_AO6;
  assign CLBLM_R_X59Y100_SLICE_X88Y100_B = CLBLM_R_X59Y100_SLICE_X88Y100_BO6;
  assign CLBLM_R_X59Y100_SLICE_X88Y100_C = CLBLM_R_X59Y100_SLICE_X88Y100_CO6;
  assign CLBLM_R_X59Y100_SLICE_X88Y100_D = CLBLM_R_X59Y100_SLICE_X88Y100_DO6;
  assign CLBLM_R_X59Y100_SLICE_X88Y100_AMUX = CLBLM_R_X59Y100_SLICE_X88Y100_AO5;
  assign CLBLM_R_X59Y100_SLICE_X88Y100_BMUX = CLBLM_R_X59Y100_SLICE_X88Y100_B5Q;
  assign CLBLM_R_X59Y100_SLICE_X88Y100_CMUX = CLBLM_R_X59Y100_SLICE_X88Y100_C5Q;
  assign CLBLM_R_X59Y100_SLICE_X89Y100_A = CLBLM_R_X59Y100_SLICE_X89Y100_AO6;
  assign CLBLM_R_X59Y100_SLICE_X89Y100_B = CLBLM_R_X59Y100_SLICE_X89Y100_BO6;
  assign CLBLM_R_X59Y100_SLICE_X89Y100_C = CLBLM_R_X59Y100_SLICE_X89Y100_CO6;
  assign CLBLM_R_X59Y100_SLICE_X89Y100_D = CLBLM_R_X59Y100_SLICE_X89Y100_DO6;
  assign CLBLM_R_X59Y101_SLICE_X88Y101_A = CLBLM_R_X59Y101_SLICE_X88Y101_AO6;
  assign CLBLM_R_X59Y101_SLICE_X88Y101_B = CLBLM_R_X59Y101_SLICE_X88Y101_BO6;
  assign CLBLM_R_X59Y101_SLICE_X88Y101_C = CLBLM_R_X59Y101_SLICE_X88Y101_CO6;
  assign CLBLM_R_X59Y101_SLICE_X88Y101_D = CLBLM_R_X59Y101_SLICE_X88Y101_DO6;
  assign CLBLM_R_X59Y101_SLICE_X88Y101_DMUX = CLBLM_R_X59Y101_SLICE_X88Y101_DO6;
  assign CLBLM_R_X59Y101_SLICE_X89Y101_A = CLBLM_R_X59Y101_SLICE_X89Y101_AO6;
  assign CLBLM_R_X59Y101_SLICE_X89Y101_B = CLBLM_R_X59Y101_SLICE_X89Y101_BO6;
  assign CLBLM_R_X59Y101_SLICE_X89Y101_C = CLBLM_R_X59Y101_SLICE_X89Y101_CO6;
  assign CLBLM_R_X59Y101_SLICE_X89Y101_D = CLBLM_R_X59Y101_SLICE_X89Y101_DO6;
  assign CLBLM_R_X59Y101_SLICE_X89Y101_BMUX = CLBLM_R_X59Y101_SLICE_X89Y101_BO6;
  assign CLBLM_R_X59Y102_SLICE_X88Y102_A = CLBLM_R_X59Y102_SLICE_X88Y102_AO6;
  assign CLBLM_R_X59Y102_SLICE_X88Y102_B = CLBLM_R_X59Y102_SLICE_X88Y102_BO6;
  assign CLBLM_R_X59Y102_SLICE_X88Y102_C = CLBLM_R_X59Y102_SLICE_X88Y102_CO6;
  assign CLBLM_R_X59Y102_SLICE_X88Y102_D = CLBLM_R_X59Y102_SLICE_X88Y102_DO6;
  assign CLBLM_R_X59Y102_SLICE_X89Y102_A = CLBLM_R_X59Y102_SLICE_X89Y102_AO6;
  assign CLBLM_R_X59Y102_SLICE_X89Y102_B = CLBLM_R_X59Y102_SLICE_X89Y102_BO6;
  assign CLBLM_R_X59Y102_SLICE_X89Y102_C = CLBLM_R_X59Y102_SLICE_X89Y102_CO6;
  assign CLBLM_R_X59Y102_SLICE_X89Y102_D = CLBLM_R_X59Y102_SLICE_X89Y102_DO6;
  assign CLBLM_R_X59Y102_SLICE_X89Y102_DMUX = CLBLM_R_X59Y102_SLICE_X89Y102_DO6;
  assign CLBLM_R_X59Y103_SLICE_X88Y103_A = CLBLM_R_X59Y103_SLICE_X88Y103_AO6;
  assign CLBLM_R_X59Y103_SLICE_X88Y103_B = CLBLM_R_X59Y103_SLICE_X88Y103_BO6;
  assign CLBLM_R_X59Y103_SLICE_X88Y103_C = CLBLM_R_X59Y103_SLICE_X88Y103_CO6;
  assign CLBLM_R_X59Y103_SLICE_X88Y103_D = CLBLM_R_X59Y103_SLICE_X88Y103_DO6;
  assign CLBLM_R_X59Y103_SLICE_X88Y103_AMUX = CLBLM_R_X59Y103_SLICE_X88Y103_F7AMUX_O;
  assign CLBLM_R_X59Y103_SLICE_X89Y103_A = CLBLM_R_X59Y103_SLICE_X89Y103_AO6;
  assign CLBLM_R_X59Y103_SLICE_X89Y103_B = CLBLM_R_X59Y103_SLICE_X89Y103_BO6;
  assign CLBLM_R_X59Y103_SLICE_X89Y103_C = CLBLM_R_X59Y103_SLICE_X89Y103_CO6;
  assign CLBLM_R_X59Y103_SLICE_X89Y103_D = CLBLM_R_X59Y103_SLICE_X89Y103_DO6;
  assign CLBLM_R_X59Y103_SLICE_X89Y103_AMUX = CLBLM_R_X59Y103_SLICE_X89Y103_A5Q;
  assign CLBLM_R_X59Y104_SLICE_X88Y104_A = CLBLM_R_X59Y104_SLICE_X88Y104_AO6;
  assign CLBLM_R_X59Y104_SLICE_X88Y104_B = CLBLM_R_X59Y104_SLICE_X88Y104_BO6;
  assign CLBLM_R_X59Y104_SLICE_X88Y104_C = CLBLM_R_X59Y104_SLICE_X88Y104_CO6;
  assign CLBLM_R_X59Y104_SLICE_X88Y104_D = CLBLM_R_X59Y104_SLICE_X88Y104_DO6;
  assign CLBLM_R_X59Y104_SLICE_X88Y104_AMUX = CLBLM_R_X59Y104_SLICE_X88Y104_AO5;
  assign CLBLM_R_X59Y104_SLICE_X88Y104_BMUX = CLBLM_R_X59Y104_SLICE_X88Y104_BO6;
  assign CLBLM_R_X59Y104_SLICE_X88Y104_CMUX = CLBLM_R_X59Y104_SLICE_X88Y104_CO6;
  assign CLBLM_R_X59Y104_SLICE_X89Y104_A = CLBLM_R_X59Y104_SLICE_X89Y104_AO6;
  assign CLBLM_R_X59Y104_SLICE_X89Y104_B = CLBLM_R_X59Y104_SLICE_X89Y104_BO6;
  assign CLBLM_R_X59Y104_SLICE_X89Y104_C = CLBLM_R_X59Y104_SLICE_X89Y104_CO6;
  assign CLBLM_R_X59Y104_SLICE_X89Y104_D = CLBLM_R_X59Y104_SLICE_X89Y104_DO6;
  assign CLBLM_R_X59Y104_SLICE_X89Y104_AMUX = CLBLM_R_X59Y104_SLICE_X89Y104_F7AMUX_O;
  assign CLBLM_R_X59Y105_SLICE_X88Y105_A = CLBLM_R_X59Y105_SLICE_X88Y105_AO6;
  assign CLBLM_R_X59Y105_SLICE_X88Y105_B = CLBLM_R_X59Y105_SLICE_X88Y105_BO6;
  assign CLBLM_R_X59Y105_SLICE_X88Y105_C = CLBLM_R_X59Y105_SLICE_X88Y105_CO6;
  assign CLBLM_R_X59Y105_SLICE_X88Y105_D = CLBLM_R_X59Y105_SLICE_X88Y105_DO6;
  assign CLBLM_R_X59Y105_SLICE_X88Y105_AMUX = CLBLM_R_X59Y105_SLICE_X88Y105_F7AMUX_O;
  assign CLBLM_R_X59Y105_SLICE_X89Y105_A = CLBLM_R_X59Y105_SLICE_X89Y105_AO6;
  assign CLBLM_R_X59Y105_SLICE_X89Y105_B = CLBLM_R_X59Y105_SLICE_X89Y105_BO6;
  assign CLBLM_R_X59Y105_SLICE_X89Y105_C = CLBLM_R_X59Y105_SLICE_X89Y105_CO6;
  assign CLBLM_R_X59Y105_SLICE_X89Y105_D = CLBLM_R_X59Y105_SLICE_X89Y105_DO6;
  assign CLBLM_R_X59Y105_SLICE_X89Y105_AMUX = CLBLM_R_X59Y105_SLICE_X89Y105_F7AMUX_O;
  assign CLBLM_R_X59Y106_SLICE_X88Y106_A = CLBLM_R_X59Y106_SLICE_X88Y106_AO6;
  assign CLBLM_R_X59Y106_SLICE_X88Y106_B = CLBLM_R_X59Y106_SLICE_X88Y106_BO6;
  assign CLBLM_R_X59Y106_SLICE_X88Y106_C = CLBLM_R_X59Y106_SLICE_X88Y106_CO6;
  assign CLBLM_R_X59Y106_SLICE_X88Y106_D = CLBLM_R_X59Y106_SLICE_X88Y106_DO6;
  assign CLBLM_R_X59Y106_SLICE_X89Y106_A = CLBLM_R_X59Y106_SLICE_X89Y106_AO6;
  assign CLBLM_R_X59Y106_SLICE_X89Y106_B = CLBLM_R_X59Y106_SLICE_X89Y106_BO6;
  assign CLBLM_R_X59Y106_SLICE_X89Y106_C = CLBLM_R_X59Y106_SLICE_X89Y106_CO6;
  assign CLBLM_R_X59Y106_SLICE_X89Y106_D = CLBLM_R_X59Y106_SLICE_X89Y106_DO6;
  assign CLBLM_R_X59Y106_SLICE_X89Y106_AMUX = CLBLM_R_X59Y106_SLICE_X89Y106_AO5;
  assign CLBLM_R_X59Y107_SLICE_X88Y107_A = CLBLM_R_X59Y107_SLICE_X88Y107_AO6;
  assign CLBLM_R_X59Y107_SLICE_X88Y107_B = CLBLM_R_X59Y107_SLICE_X88Y107_BO6;
  assign CLBLM_R_X59Y107_SLICE_X88Y107_C = CLBLM_R_X59Y107_SLICE_X88Y107_CO6;
  assign CLBLM_R_X59Y107_SLICE_X88Y107_D = CLBLM_R_X59Y107_SLICE_X88Y107_DO6;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_A = CLBLM_R_X59Y107_SLICE_X89Y107_AO6;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_B = CLBLM_R_X59Y107_SLICE_X89Y107_BO6;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_C = CLBLM_R_X59Y107_SLICE_X89Y107_CO6;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_D = CLBLM_R_X59Y107_SLICE_X89Y107_DO6;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_AMUX = CLBLM_R_X59Y107_SLICE_X89Y107_A_XOR;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_BMUX = CLBLM_R_X59Y107_SLICE_X89Y107_B_XOR;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_CMUX = CLBLM_R_X59Y107_SLICE_X89Y107_C_XOR;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_DMUX = CLBLM_R_X59Y107_SLICE_X89Y107_D_XOR;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_A = CLBLM_R_X59Y108_SLICE_X88Y108_AO6;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_B = CLBLM_R_X59Y108_SLICE_X88Y108_BO6;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_C = CLBLM_R_X59Y108_SLICE_X88Y108_CO6;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_D = CLBLM_R_X59Y108_SLICE_X88Y108_DO6;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_AMUX = CLBLM_R_X59Y108_SLICE_X88Y108_A_XOR;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_BMUX = CLBLM_R_X59Y108_SLICE_X88Y108_B_XOR;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_CMUX = CLBLM_R_X59Y108_SLICE_X88Y108_C_XOR;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_DMUX = CLBLM_R_X59Y108_SLICE_X88Y108_D_XOR;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_A = CLBLM_R_X59Y108_SLICE_X89Y108_AO6;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_B = CLBLM_R_X59Y108_SLICE_X89Y108_BO6;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_C = CLBLM_R_X59Y108_SLICE_X89Y108_CO6;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_D = CLBLM_R_X59Y108_SLICE_X89Y108_DO6;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_AMUX = CLBLM_R_X59Y108_SLICE_X89Y108_A_XOR;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_BMUX = CLBLM_R_X59Y108_SLICE_X89Y108_B_XOR;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_CMUX = CLBLM_R_X59Y108_SLICE_X89Y108_C_XOR;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_DMUX = CLBLM_R_X59Y108_SLICE_X89Y108_D_XOR;
  assign CLBLM_R_X59Y109_SLICE_X88Y109_A = CLBLM_R_X59Y109_SLICE_X88Y109_AO6;
  assign CLBLM_R_X59Y109_SLICE_X88Y109_B = CLBLM_R_X59Y109_SLICE_X88Y109_BO6;
  assign CLBLM_R_X59Y109_SLICE_X88Y109_C = CLBLM_R_X59Y109_SLICE_X88Y109_CO6;
  assign CLBLM_R_X59Y109_SLICE_X88Y109_D = CLBLM_R_X59Y109_SLICE_X88Y109_DO6;
  assign CLBLM_R_X59Y109_SLICE_X88Y109_AMUX = CLBLM_R_X59Y109_SLICE_X88Y109_A_XOR;
  assign CLBLM_R_X59Y109_SLICE_X88Y109_BMUX = CLBLM_R_X59Y109_SLICE_X88Y109_B_XOR;
  assign CLBLM_R_X59Y109_SLICE_X88Y109_CMUX = CLBLM_R_X59Y109_SLICE_X88Y109_C_XOR;
  assign CLBLM_R_X59Y109_SLICE_X88Y109_DMUX = CLBLM_R_X59Y109_SLICE_X88Y109_D_XOR;
  assign CLBLM_R_X59Y109_SLICE_X89Y109_A = CLBLM_R_X59Y109_SLICE_X89Y109_AO6;
  assign CLBLM_R_X59Y109_SLICE_X89Y109_B = CLBLM_R_X59Y109_SLICE_X89Y109_BO6;
  assign CLBLM_R_X59Y109_SLICE_X89Y109_C = CLBLM_R_X59Y109_SLICE_X89Y109_CO6;
  assign CLBLM_R_X59Y109_SLICE_X89Y109_D = CLBLM_R_X59Y109_SLICE_X89Y109_DO6;
  assign CLBLM_R_X59Y109_SLICE_X89Y109_AMUX = CLBLM_R_X59Y109_SLICE_X89Y109_A_XOR;
  assign CLBLM_R_X59Y109_SLICE_X89Y109_BMUX = CLBLM_R_X59Y109_SLICE_X89Y109_B_XOR;
  assign CLBLM_R_X59Y109_SLICE_X89Y109_CMUX = CLBLM_R_X59Y109_SLICE_X89Y109_C_XOR;
  assign CLBLM_R_X59Y110_SLICE_X88Y110_A = CLBLM_R_X59Y110_SLICE_X88Y110_AO6;
  assign CLBLM_R_X59Y110_SLICE_X88Y110_B = CLBLM_R_X59Y110_SLICE_X88Y110_BO6;
  assign CLBLM_R_X59Y110_SLICE_X88Y110_C = CLBLM_R_X59Y110_SLICE_X88Y110_CO6;
  assign CLBLM_R_X59Y110_SLICE_X88Y110_D = CLBLM_R_X59Y110_SLICE_X88Y110_DO6;
  assign CLBLM_R_X59Y110_SLICE_X88Y110_AMUX = CLBLM_R_X59Y110_SLICE_X88Y110_A_XOR;
  assign CLBLM_R_X59Y110_SLICE_X88Y110_BMUX = CLBLM_R_X59Y110_SLICE_X88Y110_B_XOR;
  assign CLBLM_R_X59Y110_SLICE_X88Y110_CMUX = CLBLM_R_X59Y110_SLICE_X88Y110_C_XOR;
  assign CLBLM_R_X59Y110_SLICE_X88Y110_DMUX = CLBLM_R_X59Y110_SLICE_X88Y110_D_XOR;
  assign CLBLM_R_X59Y110_SLICE_X89Y110_A = CLBLM_R_X59Y110_SLICE_X89Y110_AO6;
  assign CLBLM_R_X59Y110_SLICE_X89Y110_B = CLBLM_R_X59Y110_SLICE_X89Y110_BO6;
  assign CLBLM_R_X59Y110_SLICE_X89Y110_C = CLBLM_R_X59Y110_SLICE_X89Y110_CO6;
  assign CLBLM_R_X59Y110_SLICE_X89Y110_D = CLBLM_R_X59Y110_SLICE_X89Y110_DO6;
  assign CLBLM_R_X59Y110_SLICE_X89Y110_DMUX = CLBLM_R_X59Y110_SLICE_X89Y110_DO6;
  assign CLBLM_R_X59Y111_SLICE_X88Y111_A = CLBLM_R_X59Y111_SLICE_X88Y111_AO6;
  assign CLBLM_R_X59Y111_SLICE_X88Y111_B = CLBLM_R_X59Y111_SLICE_X88Y111_BO6;
  assign CLBLM_R_X59Y111_SLICE_X88Y111_C = CLBLM_R_X59Y111_SLICE_X88Y111_CO6;
  assign CLBLM_R_X59Y111_SLICE_X88Y111_D = CLBLM_R_X59Y111_SLICE_X88Y111_DO6;
  assign CLBLM_R_X59Y111_SLICE_X88Y111_AMUX = CLBLM_R_X59Y111_SLICE_X88Y111_AO6;
  assign CLBLM_R_X59Y111_SLICE_X89Y111_A = CLBLM_R_X59Y111_SLICE_X89Y111_AO6;
  assign CLBLM_R_X59Y111_SLICE_X89Y111_B = CLBLM_R_X59Y111_SLICE_X89Y111_BO6;
  assign CLBLM_R_X59Y111_SLICE_X89Y111_C = CLBLM_R_X59Y111_SLICE_X89Y111_CO6;
  assign CLBLM_R_X59Y111_SLICE_X89Y111_D = CLBLM_R_X59Y111_SLICE_X89Y111_DO6;
  assign CLBLM_R_X59Y112_SLICE_X88Y112_A = CLBLM_R_X59Y112_SLICE_X88Y112_AO6;
  assign CLBLM_R_X59Y112_SLICE_X88Y112_B = CLBLM_R_X59Y112_SLICE_X88Y112_BO6;
  assign CLBLM_R_X59Y112_SLICE_X88Y112_C = CLBLM_R_X59Y112_SLICE_X88Y112_CO6;
  assign CLBLM_R_X59Y112_SLICE_X88Y112_D = CLBLM_R_X59Y112_SLICE_X88Y112_DO6;
  assign CLBLM_R_X59Y112_SLICE_X89Y112_A = CLBLM_R_X59Y112_SLICE_X89Y112_AO6;
  assign CLBLM_R_X59Y112_SLICE_X89Y112_B = CLBLM_R_X59Y112_SLICE_X89Y112_BO6;
  assign CLBLM_R_X59Y112_SLICE_X89Y112_C = CLBLM_R_X59Y112_SLICE_X89Y112_CO6;
  assign CLBLM_R_X59Y112_SLICE_X89Y112_D = CLBLM_R_X59Y112_SLICE_X89Y112_DO6;
  assign CLBLM_R_X63Y94_SLICE_X94Y94_A = CLBLM_R_X63Y94_SLICE_X94Y94_AO6;
  assign CLBLM_R_X63Y94_SLICE_X94Y94_B = CLBLM_R_X63Y94_SLICE_X94Y94_BO6;
  assign CLBLM_R_X63Y94_SLICE_X94Y94_C = CLBLM_R_X63Y94_SLICE_X94Y94_CO6;
  assign CLBLM_R_X63Y94_SLICE_X94Y94_D = CLBLM_R_X63Y94_SLICE_X94Y94_DO6;
  assign CLBLM_R_X63Y94_SLICE_X95Y94_A = CLBLM_R_X63Y94_SLICE_X95Y94_AO6;
  assign CLBLM_R_X63Y94_SLICE_X95Y94_B = CLBLM_R_X63Y94_SLICE_X95Y94_BO6;
  assign CLBLM_R_X63Y94_SLICE_X95Y94_C = CLBLM_R_X63Y94_SLICE_X95Y94_CO6;
  assign CLBLM_R_X63Y94_SLICE_X95Y94_D = CLBLM_R_X63Y94_SLICE_X95Y94_DO6;
  assign CLBLM_R_X63Y95_SLICE_X94Y95_A = CLBLM_R_X63Y95_SLICE_X94Y95_AO6;
  assign CLBLM_R_X63Y95_SLICE_X94Y95_B = CLBLM_R_X63Y95_SLICE_X94Y95_BO6;
  assign CLBLM_R_X63Y95_SLICE_X94Y95_C = CLBLM_R_X63Y95_SLICE_X94Y95_CO6;
  assign CLBLM_R_X63Y95_SLICE_X94Y95_D = CLBLM_R_X63Y95_SLICE_X94Y95_DO6;
  assign CLBLM_R_X63Y95_SLICE_X94Y95_AMUX = CLBLM_R_X63Y95_SLICE_X94Y95_AO5;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_A = CLBLM_R_X63Y95_SLICE_X95Y95_AO6;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_B = CLBLM_R_X63Y95_SLICE_X95Y95_BO6;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_C = CLBLM_R_X63Y95_SLICE_X95Y95_CO6;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_D = CLBLM_R_X63Y95_SLICE_X95Y95_DO6;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_AMUX = CLBLM_R_X63Y95_SLICE_X95Y95_AO5;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_BMUX = CLBLM_R_X63Y95_SLICE_X95Y95_B5Q;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_CMUX = CLBLM_R_X63Y95_SLICE_X95Y95_C5Q;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_DMUX = CLBLM_R_X63Y95_SLICE_X95Y95_D5Q;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_A = CLBLM_R_X63Y96_SLICE_X94Y96_AO6;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_B = CLBLM_R_X63Y96_SLICE_X94Y96_BO6;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_C = CLBLM_R_X63Y96_SLICE_X94Y96_CO6;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_D = CLBLM_R_X63Y96_SLICE_X94Y96_DO6;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_AMUX = CLBLM_R_X63Y96_SLICE_X94Y96_AO5;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_BMUX = CLBLM_R_X63Y96_SLICE_X94Y96_BO5;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_CMUX = CLBLM_R_X63Y96_SLICE_X94Y96_CO5;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_A = CLBLM_R_X63Y96_SLICE_X95Y96_AO6;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_B = CLBLM_R_X63Y96_SLICE_X95Y96_BO6;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_C = CLBLM_R_X63Y96_SLICE_X95Y96_CO6;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_D = CLBLM_R_X63Y96_SLICE_X95Y96_DO6;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_AMUX = CLBLM_R_X63Y96_SLICE_X95Y96_AO5;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_A = CLBLM_R_X63Y97_SLICE_X94Y97_AO6;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_B = CLBLM_R_X63Y97_SLICE_X94Y97_BO6;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_C = CLBLM_R_X63Y97_SLICE_X94Y97_CO6;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_D = CLBLM_R_X63Y97_SLICE_X94Y97_DO6;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_AMUX = CLBLM_R_X63Y97_SLICE_X94Y97_F7AMUX_O;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_CMUX = CLBLM_R_X63Y97_SLICE_X94Y97_CO5;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_A = CLBLM_R_X63Y97_SLICE_X95Y97_AO6;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_B = CLBLM_R_X63Y97_SLICE_X95Y97_BO6;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_C = CLBLM_R_X63Y97_SLICE_X95Y97_CO6;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_D = CLBLM_R_X63Y97_SLICE_X95Y97_DO6;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_AMUX = CLBLM_R_X63Y97_SLICE_X95Y97_F7AMUX_O;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_CMUX = CLBLM_R_X63Y97_SLICE_X95Y97_C5Q;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_DMUX = CLBLM_R_X63Y97_SLICE_X95Y97_D5Q;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_A = CLBLM_R_X63Y98_SLICE_X94Y98_AO6;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_B = CLBLM_R_X63Y98_SLICE_X94Y98_BO6;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_C = CLBLM_R_X63Y98_SLICE_X94Y98_CO6;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_D = CLBLM_R_X63Y98_SLICE_X94Y98_DO6;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_AMUX = CLBLM_R_X63Y98_SLICE_X94Y98_F7AMUX_O;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_CMUX = CLBLM_R_X63Y98_SLICE_X94Y98_C5Q;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_A = CLBLM_R_X63Y98_SLICE_X95Y98_AO6;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_B = CLBLM_R_X63Y98_SLICE_X95Y98_BO6;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_C = CLBLM_R_X63Y98_SLICE_X95Y98_CO6;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_D = CLBLM_R_X63Y98_SLICE_X95Y98_DO6;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_AMUX = CLBLM_R_X63Y98_SLICE_X95Y98_A5Q;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_BMUX = CLBLM_R_X63Y98_SLICE_X95Y98_B5Q;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_CMUX = CLBLM_R_X63Y98_SLICE_X95Y98_C5Q;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_DMUX = CLBLM_R_X63Y98_SLICE_X95Y98_D5Q;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_A = CLBLM_R_X63Y99_SLICE_X94Y99_AO6;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_B = CLBLM_R_X63Y99_SLICE_X94Y99_BO6;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_C = CLBLM_R_X63Y99_SLICE_X94Y99_CO6;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_D = CLBLM_R_X63Y99_SLICE_X94Y99_DO6;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_AMUX = CLBLM_R_X63Y99_SLICE_X94Y99_F7AMUX_O;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_CMUX = CLBLM_R_X63Y99_SLICE_X94Y99_C5Q;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_DMUX = CLBLM_R_X63Y99_SLICE_X94Y99_DO5;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_A = CLBLM_R_X63Y99_SLICE_X95Y99_AO6;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_B = CLBLM_R_X63Y99_SLICE_X95Y99_BO6;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_C = CLBLM_R_X63Y99_SLICE_X95Y99_CO6;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_D = CLBLM_R_X63Y99_SLICE_X95Y99_DO6;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_AMUX = CLBLM_R_X63Y99_SLICE_X95Y99_A5Q;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_BMUX = CLBLM_R_X63Y99_SLICE_X95Y99_B5Q;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_CMUX = CLBLM_R_X63Y99_SLICE_X95Y99_C5Q;
  assign CLBLM_R_X63Y100_SLICE_X94Y100_A = CLBLM_R_X63Y100_SLICE_X94Y100_AO6;
  assign CLBLM_R_X63Y100_SLICE_X94Y100_B = CLBLM_R_X63Y100_SLICE_X94Y100_BO6;
  assign CLBLM_R_X63Y100_SLICE_X94Y100_C = CLBLM_R_X63Y100_SLICE_X94Y100_CO6;
  assign CLBLM_R_X63Y100_SLICE_X94Y100_D = CLBLM_R_X63Y100_SLICE_X94Y100_DO6;
  assign CLBLM_R_X63Y100_SLICE_X95Y100_A = CLBLM_R_X63Y100_SLICE_X95Y100_AO6;
  assign CLBLM_R_X63Y100_SLICE_X95Y100_B = CLBLM_R_X63Y100_SLICE_X95Y100_BO6;
  assign CLBLM_R_X63Y100_SLICE_X95Y100_C = CLBLM_R_X63Y100_SLICE_X95Y100_CO6;
  assign CLBLM_R_X63Y100_SLICE_X95Y100_D = CLBLM_R_X63Y100_SLICE_X95Y100_DO6;
  assign CLBLM_R_X63Y100_SLICE_X95Y100_AMUX = CLBLM_R_X63Y100_SLICE_X95Y100_A5Q;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_A = CLBLM_R_X63Y101_SLICE_X94Y101_AO6;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_B = CLBLM_R_X63Y101_SLICE_X94Y101_BO6;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_C = CLBLM_R_X63Y101_SLICE_X94Y101_CO6;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_D = CLBLM_R_X63Y101_SLICE_X94Y101_DO6;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_A = CLBLM_R_X63Y101_SLICE_X95Y101_AO6;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_B = CLBLM_R_X63Y101_SLICE_X95Y101_BO6;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_C = CLBLM_R_X63Y101_SLICE_X95Y101_CO6;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_D = CLBLM_R_X63Y101_SLICE_X95Y101_DO6;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_A = CLBLM_R_X63Y102_SLICE_X94Y102_AO6;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_B = CLBLM_R_X63Y102_SLICE_X94Y102_BO6;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_C = CLBLM_R_X63Y102_SLICE_X94Y102_CO6;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_D = CLBLM_R_X63Y102_SLICE_X94Y102_DO6;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_A = CLBLM_R_X63Y102_SLICE_X95Y102_AO6;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_B = CLBLM_R_X63Y102_SLICE_X95Y102_BO6;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_C = CLBLM_R_X63Y102_SLICE_X95Y102_CO6;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_D = CLBLM_R_X63Y102_SLICE_X95Y102_DO6;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_A = CLBLM_R_X63Y103_SLICE_X94Y103_AO6;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_B = CLBLM_R_X63Y103_SLICE_X94Y103_BO6;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_C = CLBLM_R_X63Y103_SLICE_X94Y103_CO6;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_D = CLBLM_R_X63Y103_SLICE_X94Y103_DO6;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_A = CLBLM_R_X63Y103_SLICE_X95Y103_AO6;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_B = CLBLM_R_X63Y103_SLICE_X95Y103_BO6;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_C = CLBLM_R_X63Y103_SLICE_X95Y103_CO6;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_D = CLBLM_R_X63Y103_SLICE_X95Y103_DO6;
  assign CLBLM_R_X63Y104_SLICE_X94Y104_A = CLBLM_R_X63Y104_SLICE_X94Y104_AO6;
  assign CLBLM_R_X63Y104_SLICE_X94Y104_B = CLBLM_R_X63Y104_SLICE_X94Y104_BO6;
  assign CLBLM_R_X63Y104_SLICE_X94Y104_C = CLBLM_R_X63Y104_SLICE_X94Y104_CO6;
  assign CLBLM_R_X63Y104_SLICE_X94Y104_D = CLBLM_R_X63Y104_SLICE_X94Y104_DO6;
  assign CLBLM_R_X63Y104_SLICE_X94Y104_CMUX = CLBLM_R_X63Y104_SLICE_X94Y104_CO6;
  assign CLBLM_R_X63Y104_SLICE_X95Y104_A = CLBLM_R_X63Y104_SLICE_X95Y104_AO6;
  assign CLBLM_R_X63Y104_SLICE_X95Y104_B = CLBLM_R_X63Y104_SLICE_X95Y104_BO6;
  assign CLBLM_R_X63Y104_SLICE_X95Y104_C = CLBLM_R_X63Y104_SLICE_X95Y104_CO6;
  assign CLBLM_R_X63Y104_SLICE_X95Y104_D = CLBLM_R_X63Y104_SLICE_X95Y104_DO6;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_A = CLBLM_R_X63Y105_SLICE_X94Y105_AO6;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_B = CLBLM_R_X63Y105_SLICE_X94Y105_BO6;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_C = CLBLM_R_X63Y105_SLICE_X94Y105_CO6;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_D = CLBLM_R_X63Y105_SLICE_X94Y105_DO6;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_AMUX = CLBLM_R_X63Y105_SLICE_X94Y105_A_XOR;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_BMUX = CLBLM_R_X63Y105_SLICE_X94Y105_B_XOR;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_CMUX = CLBLM_R_X63Y105_SLICE_X94Y105_C_XOR;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_DMUX = CLBLM_R_X63Y105_SLICE_X94Y105_D_XOR;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_A = CLBLM_R_X63Y105_SLICE_X95Y105_AO6;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_B = CLBLM_R_X63Y105_SLICE_X95Y105_BO6;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_C = CLBLM_R_X63Y105_SLICE_X95Y105_CO6;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_D = CLBLM_R_X63Y105_SLICE_X95Y105_DO6;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_AMUX = CLBLM_R_X63Y105_SLICE_X95Y105_A_XOR;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_BMUX = CLBLM_R_X63Y105_SLICE_X95Y105_B_XOR;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_CMUX = CLBLM_R_X63Y105_SLICE_X95Y105_C_XOR;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_DMUX = CLBLM_R_X63Y105_SLICE_X95Y105_D_XOR;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_A = CLBLM_R_X63Y106_SLICE_X94Y106_AO6;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_B = CLBLM_R_X63Y106_SLICE_X94Y106_BO6;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_C = CLBLM_R_X63Y106_SLICE_X94Y106_CO6;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_D = CLBLM_R_X63Y106_SLICE_X94Y106_DO6;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_AMUX = CLBLM_R_X63Y106_SLICE_X94Y106_A_XOR;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_BMUX = CLBLM_R_X63Y106_SLICE_X94Y106_B_XOR;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_CMUX = CLBLM_R_X63Y106_SLICE_X94Y106_C_XOR;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_DMUX = CLBLM_R_X63Y106_SLICE_X94Y106_D_XOR;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_A = CLBLM_R_X63Y106_SLICE_X95Y106_AO6;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_B = CLBLM_R_X63Y106_SLICE_X95Y106_BO6;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_C = CLBLM_R_X63Y106_SLICE_X95Y106_CO6;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_D = CLBLM_R_X63Y106_SLICE_X95Y106_DO6;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_AMUX = CLBLM_R_X63Y106_SLICE_X95Y106_A_XOR;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_BMUX = CLBLM_R_X63Y106_SLICE_X95Y106_B_XOR;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_CMUX = CLBLM_R_X63Y106_SLICE_X95Y106_C_XOR;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_DMUX = CLBLM_R_X63Y106_SLICE_X95Y106_D_XOR;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_A = CLBLM_R_X63Y107_SLICE_X94Y107_AO6;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_B = CLBLM_R_X63Y107_SLICE_X94Y107_BO6;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_C = CLBLM_R_X63Y107_SLICE_X94Y107_CO6;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_D = CLBLM_R_X63Y107_SLICE_X94Y107_DO6;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_AMUX = CLBLM_R_X63Y107_SLICE_X94Y107_A_XOR;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_BMUX = CLBLM_R_X63Y107_SLICE_X94Y107_B_XOR;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_CMUX = CLBLM_R_X63Y107_SLICE_X94Y107_C_XOR;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_DMUX = CLBLM_R_X63Y107_SLICE_X94Y107_D_XOR;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_A = CLBLM_R_X63Y107_SLICE_X95Y107_AO6;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_B = CLBLM_R_X63Y107_SLICE_X95Y107_BO6;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_C = CLBLM_R_X63Y107_SLICE_X95Y107_CO6;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_D = CLBLM_R_X63Y107_SLICE_X95Y107_DO6;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_AMUX = CLBLM_R_X63Y107_SLICE_X95Y107_A_XOR;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_BMUX = CLBLM_R_X63Y107_SLICE_X95Y107_B_XOR;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_CMUX = CLBLM_R_X63Y107_SLICE_X95Y107_C_XOR;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_DMUX = CLBLM_R_X63Y107_SLICE_X95Y107_D_XOR;
  assign CLBLM_R_X63Y108_SLICE_X94Y108_A = CLBLM_R_X63Y108_SLICE_X94Y108_AO6;
  assign CLBLM_R_X63Y108_SLICE_X94Y108_B = CLBLM_R_X63Y108_SLICE_X94Y108_BO6;
  assign CLBLM_R_X63Y108_SLICE_X94Y108_C = CLBLM_R_X63Y108_SLICE_X94Y108_CO6;
  assign CLBLM_R_X63Y108_SLICE_X94Y108_D = CLBLM_R_X63Y108_SLICE_X94Y108_DO6;
  assign CLBLM_R_X63Y108_SLICE_X94Y108_AMUX = CLBLM_R_X63Y108_SLICE_X94Y108_A_XOR;
  assign CLBLM_R_X63Y108_SLICE_X94Y108_BMUX = CLBLM_R_X63Y108_SLICE_X94Y108_B_XOR;
  assign CLBLM_R_X63Y108_SLICE_X94Y108_CMUX = CLBLM_R_X63Y108_SLICE_X94Y108_C_XOR;
  assign CLBLM_R_X63Y108_SLICE_X94Y108_DMUX = CLBLM_R_X63Y108_SLICE_X94Y108_D_XOR;
  assign CLBLM_R_X63Y108_SLICE_X95Y108_A = CLBLM_R_X63Y108_SLICE_X95Y108_AO6;
  assign CLBLM_R_X63Y108_SLICE_X95Y108_B = CLBLM_R_X63Y108_SLICE_X95Y108_BO6;
  assign CLBLM_R_X63Y108_SLICE_X95Y108_C = CLBLM_R_X63Y108_SLICE_X95Y108_CO6;
  assign CLBLM_R_X63Y108_SLICE_X95Y108_D = CLBLM_R_X63Y108_SLICE_X95Y108_DO6;
  assign CLBLM_R_X63Y108_SLICE_X95Y108_AMUX = CLBLM_R_X63Y108_SLICE_X95Y108_A_XOR;
  assign CLBLM_R_X63Y108_SLICE_X95Y108_BMUX = CLBLM_R_X63Y108_SLICE_X95Y108_B_XOR;
  assign CLBLM_R_X63Y108_SLICE_X95Y108_CMUX = CLBLM_R_X63Y108_SLICE_X95Y108_C_XOR;
  assign CLBLM_R_X63Y108_SLICE_X95Y108_DMUX = CLBLM_R_X63Y108_SLICE_X95Y108_D_XOR;
  assign CLBLM_R_X63Y109_SLICE_X94Y109_A = CLBLM_R_X63Y109_SLICE_X94Y109_AO6;
  assign CLBLM_R_X63Y109_SLICE_X94Y109_B = CLBLM_R_X63Y109_SLICE_X94Y109_BO6;
  assign CLBLM_R_X63Y109_SLICE_X94Y109_C = CLBLM_R_X63Y109_SLICE_X94Y109_CO6;
  assign CLBLM_R_X63Y109_SLICE_X94Y109_D = CLBLM_R_X63Y109_SLICE_X94Y109_DO6;
  assign CLBLM_R_X63Y109_SLICE_X94Y109_AMUX = CLBLM_R_X63Y109_SLICE_X94Y109_A_XOR;
  assign CLBLM_R_X63Y109_SLICE_X94Y109_BMUX = CLBLM_R_X63Y109_SLICE_X94Y109_B_XOR;
  assign CLBLM_R_X63Y109_SLICE_X94Y109_CMUX = CLBLM_R_X63Y109_SLICE_X94Y109_C_XOR;
  assign CLBLM_R_X63Y109_SLICE_X94Y109_DMUX = CLBLM_R_X63Y109_SLICE_X94Y109_D_XOR;
  assign CLBLM_R_X63Y109_SLICE_X95Y109_A = CLBLM_R_X63Y109_SLICE_X95Y109_AO6;
  assign CLBLM_R_X63Y109_SLICE_X95Y109_B = CLBLM_R_X63Y109_SLICE_X95Y109_BO6;
  assign CLBLM_R_X63Y109_SLICE_X95Y109_C = CLBLM_R_X63Y109_SLICE_X95Y109_CO6;
  assign CLBLM_R_X63Y109_SLICE_X95Y109_D = CLBLM_R_X63Y109_SLICE_X95Y109_DO6;
  assign CLBLM_R_X63Y109_SLICE_X95Y109_AMUX = CLBLM_R_X63Y109_SLICE_X95Y109_A_XOR;
  assign CLBLM_R_X63Y109_SLICE_X95Y109_BMUX = CLBLM_R_X63Y109_SLICE_X95Y109_B_XOR;
  assign CLBLM_R_X63Y109_SLICE_X95Y109_CMUX = CLBLM_R_X63Y109_SLICE_X95Y109_C_XOR;
  assign CLBLM_R_X63Y110_SLICE_X94Y110_A = CLBLM_R_X63Y110_SLICE_X94Y110_AO6;
  assign CLBLM_R_X63Y110_SLICE_X94Y110_B = CLBLM_R_X63Y110_SLICE_X94Y110_BO6;
  assign CLBLM_R_X63Y110_SLICE_X94Y110_C = CLBLM_R_X63Y110_SLICE_X94Y110_CO6;
  assign CLBLM_R_X63Y110_SLICE_X94Y110_D = CLBLM_R_X63Y110_SLICE_X94Y110_DO6;
  assign CLBLM_R_X63Y110_SLICE_X95Y110_A = CLBLM_R_X63Y110_SLICE_X95Y110_AO6;
  assign CLBLM_R_X63Y110_SLICE_X95Y110_B = CLBLM_R_X63Y110_SLICE_X95Y110_BO6;
  assign CLBLM_R_X63Y110_SLICE_X95Y110_C = CLBLM_R_X63Y110_SLICE_X95Y110_CO6;
  assign CLBLM_R_X63Y110_SLICE_X95Y110_D = CLBLM_R_X63Y110_SLICE_X95Y110_DO6;
  assign CLBLM_R_X65Y96_SLICE_X98Y96_A = CLBLM_R_X65Y96_SLICE_X98Y96_AO6;
  assign CLBLM_R_X65Y96_SLICE_X98Y96_B = CLBLM_R_X65Y96_SLICE_X98Y96_BO6;
  assign CLBLM_R_X65Y96_SLICE_X98Y96_C = CLBLM_R_X65Y96_SLICE_X98Y96_CO6;
  assign CLBLM_R_X65Y96_SLICE_X98Y96_D = CLBLM_R_X65Y96_SLICE_X98Y96_DO6;
  assign CLBLM_R_X65Y96_SLICE_X99Y96_A = CLBLM_R_X65Y96_SLICE_X99Y96_AO6;
  assign CLBLM_R_X65Y96_SLICE_X99Y96_B = CLBLM_R_X65Y96_SLICE_X99Y96_BO6;
  assign CLBLM_R_X65Y96_SLICE_X99Y96_C = CLBLM_R_X65Y96_SLICE_X99Y96_CO6;
  assign CLBLM_R_X65Y96_SLICE_X99Y96_D = CLBLM_R_X65Y96_SLICE_X99Y96_DO6;
  assign CLBLM_R_X65Y97_SLICE_X98Y97_A = CLBLM_R_X65Y97_SLICE_X98Y97_AO6;
  assign CLBLM_R_X65Y97_SLICE_X98Y97_B = CLBLM_R_X65Y97_SLICE_X98Y97_BO6;
  assign CLBLM_R_X65Y97_SLICE_X98Y97_C = CLBLM_R_X65Y97_SLICE_X98Y97_CO6;
  assign CLBLM_R_X65Y97_SLICE_X98Y97_D = CLBLM_R_X65Y97_SLICE_X98Y97_DO6;
  assign CLBLM_R_X65Y97_SLICE_X98Y97_AMUX = CLBLM_R_X65Y97_SLICE_X98Y97_AO5;
  assign CLBLM_R_X65Y97_SLICE_X99Y97_A = CLBLM_R_X65Y97_SLICE_X99Y97_AO6;
  assign CLBLM_R_X65Y97_SLICE_X99Y97_B = CLBLM_R_X65Y97_SLICE_X99Y97_BO6;
  assign CLBLM_R_X65Y97_SLICE_X99Y97_C = CLBLM_R_X65Y97_SLICE_X99Y97_CO6;
  assign CLBLM_R_X65Y97_SLICE_X99Y97_D = CLBLM_R_X65Y97_SLICE_X99Y97_DO6;
  assign CLBLM_R_X65Y98_SLICE_X98Y98_A = CLBLM_R_X65Y98_SLICE_X98Y98_AO6;
  assign CLBLM_R_X65Y98_SLICE_X98Y98_B = CLBLM_R_X65Y98_SLICE_X98Y98_BO6;
  assign CLBLM_R_X65Y98_SLICE_X98Y98_C = CLBLM_R_X65Y98_SLICE_X98Y98_CO6;
  assign CLBLM_R_X65Y98_SLICE_X98Y98_D = CLBLM_R_X65Y98_SLICE_X98Y98_DO6;
  assign CLBLM_R_X65Y98_SLICE_X98Y98_CMUX = CLBLM_R_X65Y98_SLICE_X98Y98_CO6;
  assign CLBLM_R_X65Y98_SLICE_X99Y98_A = CLBLM_R_X65Y98_SLICE_X99Y98_AO6;
  assign CLBLM_R_X65Y98_SLICE_X99Y98_B = CLBLM_R_X65Y98_SLICE_X99Y98_BO6;
  assign CLBLM_R_X65Y98_SLICE_X99Y98_C = CLBLM_R_X65Y98_SLICE_X99Y98_CO6;
  assign CLBLM_R_X65Y98_SLICE_X99Y98_D = CLBLM_R_X65Y98_SLICE_X99Y98_DO6;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_A = CLBLM_R_X65Y99_SLICE_X98Y99_AO6;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_B = CLBLM_R_X65Y99_SLICE_X98Y99_BO6;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_C = CLBLM_R_X65Y99_SLICE_X98Y99_CO6;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_D = CLBLM_R_X65Y99_SLICE_X98Y99_DO6;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_A = CLBLM_R_X65Y99_SLICE_X99Y99_AO6;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_B = CLBLM_R_X65Y99_SLICE_X99Y99_BO6;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_C = CLBLM_R_X65Y99_SLICE_X99Y99_CO6;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_D = CLBLM_R_X65Y99_SLICE_X99Y99_DO6;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_A = CLBLM_R_X65Y100_SLICE_X98Y100_AO6;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_B = CLBLM_R_X65Y100_SLICE_X98Y100_BO6;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_C = CLBLM_R_X65Y100_SLICE_X98Y100_CO6;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_D = CLBLM_R_X65Y100_SLICE_X98Y100_DO6;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_BMUX = CLBLM_R_X65Y100_SLICE_X98Y100_B_XOR;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_CMUX = CLBLM_R_X65Y100_SLICE_X98Y100_C_XOR;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_DMUX = CLBLM_R_X65Y100_SLICE_X98Y100_D_XOR;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_A = CLBLM_R_X65Y100_SLICE_X99Y100_AO6;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_B = CLBLM_R_X65Y100_SLICE_X99Y100_BO6;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_C = CLBLM_R_X65Y100_SLICE_X99Y100_CO6;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_D = CLBLM_R_X65Y100_SLICE_X99Y100_DO6;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_A = CLBLM_R_X65Y101_SLICE_X98Y101_AO6;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_B = CLBLM_R_X65Y101_SLICE_X98Y101_BO6;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_C = CLBLM_R_X65Y101_SLICE_X98Y101_CO6;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_D = CLBLM_R_X65Y101_SLICE_X98Y101_DO6;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_AMUX = CLBLM_R_X65Y101_SLICE_X98Y101_A_XOR;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_BMUX = CLBLM_R_X65Y101_SLICE_X98Y101_B_XOR;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_CMUX = CLBLM_R_X65Y101_SLICE_X98Y101_C_XOR;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_DMUX = CLBLM_R_X65Y101_SLICE_X98Y101_D_XOR;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_A = CLBLM_R_X65Y101_SLICE_X99Y101_AO6;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_B = CLBLM_R_X65Y101_SLICE_X99Y101_BO6;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_C = CLBLM_R_X65Y101_SLICE_X99Y101_CO6;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_D = CLBLM_R_X65Y101_SLICE_X99Y101_DO6;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_A = CLBLM_R_X65Y102_SLICE_X98Y102_AO6;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_B = CLBLM_R_X65Y102_SLICE_X98Y102_BO6;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_C = CLBLM_R_X65Y102_SLICE_X98Y102_CO6;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_D = CLBLM_R_X65Y102_SLICE_X98Y102_DO6;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_AMUX = CLBLM_R_X65Y102_SLICE_X98Y102_A_XOR;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_BMUX = CLBLM_R_X65Y102_SLICE_X98Y102_B_XOR;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_CMUX = CLBLM_R_X65Y102_SLICE_X98Y102_C_XOR;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_DMUX = CLBLM_R_X65Y102_SLICE_X98Y102_D_XOR;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_A = CLBLM_R_X65Y102_SLICE_X99Y102_AO6;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_B = CLBLM_R_X65Y102_SLICE_X99Y102_BO6;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_C = CLBLM_R_X65Y102_SLICE_X99Y102_CO6;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_D = CLBLM_R_X65Y102_SLICE_X99Y102_DO6;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_A = CLBLM_R_X65Y103_SLICE_X98Y103_AO6;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_B = CLBLM_R_X65Y103_SLICE_X98Y103_BO6;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_C = CLBLM_R_X65Y103_SLICE_X98Y103_CO6;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_D = CLBLM_R_X65Y103_SLICE_X98Y103_DO6;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_AMUX = CLBLM_R_X65Y103_SLICE_X98Y103_A_XOR;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_BMUX = CLBLM_R_X65Y103_SLICE_X98Y103_B_XOR;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_CMUX = CLBLM_R_X65Y103_SLICE_X98Y103_C_XOR;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_DMUX = CLBLM_R_X65Y103_SLICE_X98Y103_D_XOR;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_A = CLBLM_R_X65Y103_SLICE_X99Y103_AO6;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_B = CLBLM_R_X65Y103_SLICE_X99Y103_BO6;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_C = CLBLM_R_X65Y103_SLICE_X99Y103_CO6;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_D = CLBLM_R_X65Y103_SLICE_X99Y103_DO6;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_CMUX = CLBLM_R_X65Y103_SLICE_X99Y103_CO6;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_A = CLBLM_R_X65Y104_SLICE_X98Y104_AO6;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_B = CLBLM_R_X65Y104_SLICE_X98Y104_BO6;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_C = CLBLM_R_X65Y104_SLICE_X98Y104_CO6;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_D = CLBLM_R_X65Y104_SLICE_X98Y104_DO6;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_AMUX = CLBLM_R_X65Y104_SLICE_X98Y104_A_XOR;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_BMUX = CLBLM_R_X65Y104_SLICE_X98Y104_B_XOR;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_CMUX = CLBLM_R_X65Y104_SLICE_X98Y104_C_XOR;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_A = CLBLM_R_X65Y104_SLICE_X99Y104_AO6;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_B = CLBLM_R_X65Y104_SLICE_X99Y104_BO6;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_C = CLBLM_R_X65Y104_SLICE_X99Y104_CO6;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_D = CLBLM_R_X65Y104_SLICE_X99Y104_DO6;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_A = CLBLM_R_X65Y105_SLICE_X98Y105_AO6;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_B = CLBLM_R_X65Y105_SLICE_X98Y105_BO6;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_C = CLBLM_R_X65Y105_SLICE_X98Y105_CO6;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_D = CLBLM_R_X65Y105_SLICE_X98Y105_DO6;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_A = CLBLM_R_X65Y105_SLICE_X99Y105_AO6;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_B = CLBLM_R_X65Y105_SLICE_X99Y105_BO6;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_C = CLBLM_R_X65Y105_SLICE_X99Y105_CO6;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_D = CLBLM_R_X65Y105_SLICE_X99Y105_DO6;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_A = CLBLM_R_X65Y106_SLICE_X98Y106_AO6;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_B = CLBLM_R_X65Y106_SLICE_X98Y106_BO6;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_C = CLBLM_R_X65Y106_SLICE_X98Y106_CO6;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_D = CLBLM_R_X65Y106_SLICE_X98Y106_DO6;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_A = CLBLM_R_X65Y106_SLICE_X99Y106_AO6;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_B = CLBLM_R_X65Y106_SLICE_X99Y106_BO6;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_C = CLBLM_R_X65Y106_SLICE_X99Y106_CO6;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_D = CLBLM_R_X65Y106_SLICE_X99Y106_DO6;
  assign CLBLM_R_X65Y107_SLICE_X98Y107_A = CLBLM_R_X65Y107_SLICE_X98Y107_AO6;
  assign CLBLM_R_X65Y107_SLICE_X98Y107_B = CLBLM_R_X65Y107_SLICE_X98Y107_BO6;
  assign CLBLM_R_X65Y107_SLICE_X98Y107_C = CLBLM_R_X65Y107_SLICE_X98Y107_CO6;
  assign CLBLM_R_X65Y107_SLICE_X98Y107_D = CLBLM_R_X65Y107_SLICE_X98Y107_DO6;
  assign CLBLM_R_X65Y107_SLICE_X99Y107_A = CLBLM_R_X65Y107_SLICE_X99Y107_AO6;
  assign CLBLM_R_X65Y107_SLICE_X99Y107_B = CLBLM_R_X65Y107_SLICE_X99Y107_BO6;
  assign CLBLM_R_X65Y107_SLICE_X99Y107_C = CLBLM_R_X65Y107_SLICE_X99Y107_CO6;
  assign CLBLM_R_X65Y107_SLICE_X99Y107_D = CLBLM_R_X65Y107_SLICE_X99Y107_DO6;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_O = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_O = LIOB33_X0Y101_IOB_X0Y101_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_O = LIOB33_X0Y103_IOB_X0Y104_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_O = LIOB33_X0Y103_IOB_X0Y103_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_O = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_O = LIOB33_X0Y105_IOB_X0Y105_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_O = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_O = LIOB33_X0Y109_IOB_X0Y109_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_O = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_O = LIOB33_X0Y111_IOB_X0Y111_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_O = LIOB33_X0Y115_IOB_X0Y116_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_O = LIOB33_X0Y115_IOB_X0Y115_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y118_O = LIOB33_X0Y117_IOB_X0Y118_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_O = LIOB33_X0Y117_IOB_X0Y117_I;
  assign LIOI3_X0Y121_ILOGIC_X0Y122_O = LIOB33_X0Y121_IOB_X0Y122_I;
  assign LIOI3_X0Y121_ILOGIC_X0Y121_O = LIOB33_X0Y121_IOB_X0Y121_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y123_O = LIOB33_X0Y123_IOB_X0Y123_I;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_OQ = CLBLM_R_X49Y109_SLICE_X74Y109_DQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_OQ = CLBLM_R_X49Y111_SLICE_X74Y111_AQ;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_OQ = CLBLM_R_X49Y107_SLICE_X74Y107_AQ;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_OQ = CLBLM_R_X49Y109_SLICE_X74Y109_AQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_OQ = CLBLM_R_X49Y111_SLICE_X74Y111_BQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_OQ = CLBLM_R_X49Y111_SLICE_X74Y111_CQ;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_OQ = CLBLM_R_X49Y109_SLICE_X74Y109_BQ;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_OQ = CLBLM_R_X49Y111_SLICE_X74Y111_AQ;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_OQ = CLBLM_R_X49Y107_SLICE_X74Y107_AQ;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_OQ = CLBLM_R_X49Y109_SLICE_X74Y109_AQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_OQ = CLBLM_R_X49Y111_SLICE_X74Y111_BQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_OQ = CLBLM_L_X50Y104_SLICE_X76Y104_AQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_OQ = CLBLM_R_X49Y109_SLICE_X74Y109_CQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_OQ = CLBLM_R_X49Y105_SLICE_X75Y105_CQ;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_OQ = CLBLM_L_X50Y105_SLICE_X77Y105_AQ;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_OQ = CLBLM_L_X50Y107_SLICE_X76Y107_BQ;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_OQ = CLBLM_L_X50Y106_SLICE_X76Y106_CQ;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_OQ = CLBLM_R_X49Y111_SLICE_X75Y111_AQ;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_OQ = CLBLM_L_X50Y107_SLICE_X77Y107_AQ;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_TQ = 1'b1;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_O = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ = CLBLM_R_X49Y111_SLICE_X75Y111_A5Q;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O = LIOB33_X0Y107_IOB_X0Y107_I;
  assign LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_O = LIOB33_X0Y119_IOB_X0Y120_I;
  assign LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y119_O = LIOB33_X0Y119_IOB_X0Y119_I;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ = CLBLM_R_X49Y109_SLICE_X74Y109_DQ;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ = CLBLM_R_X49Y109_SLICE_X74Y109_CQ;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ = CLBLM_L_X50Y106_SLICE_X76Y106_AQ;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ = CLBLM_R_X49Y106_SLICE_X74Y106_AQ;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O = LIOB33_X0Y113_IOB_X0Y114_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O = LIOB33_X0Y113_IOB_X0Y113_I;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ = CLBLM_R_X49Y111_SLICE_X74Y111_CQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ = CLBLM_R_X49Y109_SLICE_X74Y109_BQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_O = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y109_OLOGIC_X1Y110_OQ = CLBLM_R_X65Y106_SLICE_X98Y106_CQ;
  assign RIOI3_X105Y109_OLOGIC_X1Y110_TQ = 1'b1;
  assign RIOI3_X105Y109_OLOGIC_X1Y109_OQ = CLBLM_R_X65Y100_SLICE_X99Y100_AQ;
  assign RIOI3_X105Y109_OLOGIC_X1Y109_TQ = 1'b1;
  assign RIOI3_X105Y111_OLOGIC_X1Y112_OQ = CLBLM_R_X65Y100_SLICE_X99Y100_BQ;
  assign RIOI3_X105Y111_OLOGIC_X1Y112_TQ = 1'b1;
  assign RIOI3_X105Y111_OLOGIC_X1Y111_OQ = CLBLM_L_X64Y106_SLICE_X97Y106_DQ;
  assign RIOI3_X105Y111_OLOGIC_X1Y111_TQ = 1'b1;
  assign RIOI3_X105Y115_OLOGIC_X1Y116_OQ = CLBLM_R_X63Y103_SLICE_X95Y103_CQ;
  assign RIOI3_X105Y115_OLOGIC_X1Y116_TQ = 1'b1;
  assign RIOI3_X105Y115_OLOGIC_X1Y115_OQ = CLBLM_R_X63Y101_SLICE_X95Y101_AQ;
  assign RIOI3_X105Y115_OLOGIC_X1Y115_TQ = 1'b1;
  assign RIOI3_X105Y117_OLOGIC_X1Y118_OQ = CLBLM_R_X65Y107_SLICE_X98Y107_AQ;
  assign RIOI3_X105Y117_OLOGIC_X1Y118_TQ = 1'b1;
  assign RIOI3_X105Y117_OLOGIC_X1Y117_OQ = CLBLM_R_X65Y107_SLICE_X98Y107_DQ;
  assign RIOI3_X105Y117_OLOGIC_X1Y117_TQ = 1'b1;
  assign RIOI3_X105Y121_OLOGIC_X1Y122_OQ = CLBLM_L_X64Y106_SLICE_X97Y106_AQ;
  assign RIOI3_X105Y121_OLOGIC_X1Y122_TQ = 1'b1;
  assign RIOI3_X105Y121_OLOGIC_X1Y121_OQ = CLBLM_R_X65Y106_SLICE_X98Y106_AQ;
  assign RIOI3_X105Y121_OLOGIC_X1Y121_TQ = 1'b1;
  assign RIOI3_X105Y123_OLOGIC_X1Y124_OQ = CLBLM_R_X65Y106_SLICE_X98Y106_BQ;
  assign RIOI3_X105Y123_OLOGIC_X1Y124_TQ = 1'b1;
  assign RIOI3_X105Y123_OLOGIC_X1Y123_OQ = CLBLM_R_X63Y103_SLICE_X95Y103_AQ;
  assign RIOI3_X105Y123_OLOGIC_X1Y123_TQ = 1'b1;
  assign RIOI3_X105Y125_OLOGIC_X1Y126_OQ = CLBLM_L_X64Y106_SLICE_X97Y106_CQ;
  assign RIOI3_X105Y125_OLOGIC_X1Y126_TQ = 1'b1;
  assign RIOI3_X105Y125_OLOGIC_X1Y125_OQ = CLBLM_L_X64Y106_SLICE_X97Y106_BQ;
  assign RIOI3_X105Y125_OLOGIC_X1Y125_TQ = 1'b1;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_OQ = CLBLM_R_X59Y102_SLICE_X88Y102_AQ;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_TQ = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_OQ = CLBLM_L_X62Y103_SLICE_X92Y103_AQ;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_TQ = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_OQ = CLBLM_L_X62Y104_SLICE_X93Y104_AQ;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_TQ = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_OQ = CLBLM_L_X62Y110_SLICE_X92Y110_AQ;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_TQ = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_OQ = CLBLM_L_X62Y106_SLICE_X93Y106_AQ;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_TQ = 1'b1;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_OQ = CLBLM_L_X60Y111_SLICE_X91Y111_BQ;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_TQ = 1'b1;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_OQ = CLBLM_L_X62Y108_SLICE_X93Y108_AQ;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_TQ = 1'b1;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_OQ = CLBLL_R_X57Y99_SLICE_X87Y99_AQ;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_TQ = 1'b1;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_OQ = CLBLM_L_X60Y111_SLICE_X91Y111_AQ;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_TQ = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_OQ = CLBLM_L_X62Y110_SLICE_X93Y110_AQ;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_TQ = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_OQ = CLBLM_L_X60Y98_SLICE_X90Y98_BQ;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_TQ = 1'b1;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_OQ = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_TQ = 1'b1;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_OQ = CLBLM_R_X65Y100_SLICE_X99Y100_CQ;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_OQ = 1'b0;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_OQ = CLBLM_R_X65Y107_SLICE_X98Y107_CQ;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_OQ = CLBLM_R_X65Y107_SLICE_X98Y107_BQ;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_OQ = CLBLM_L_X60Y110_SLICE_X91Y110_AQ;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_OQ = CLBLM_R_X59Y102_SLICE_X89Y102_AQ;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_OQ = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_OQ = CLBLM_L_X56Y111_SLICE_X84Y111_AQ;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_OQ = CLBLM_R_X63Y103_SLICE_X95Y103_BQ;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_OQ = CLBLM_R_X65Y106_SLICE_X98Y106_DQ;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_OQ = CLBLM_L_X62Y110_SLICE_X92Y110_BQ;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_OQ = CLBLM_L_X60Y111_SLICE_X90Y111_AQ;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_TQ = 1'b1;
  assign LIOB33_X0Y147_IOB_X0Y148_O = CLBLM_R_X49Y111_SLICE_X75Y111_AQ;
  assign LIOB33_X0Y147_IOB_X0Y147_O = CLBLM_L_X50Y107_SLICE_X77Y107_AQ;
  assign CLBLL_L_X52Y101_SLICE_X78Y101_A1 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X78Y101_A2 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X78Y101_A3 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X78Y101_A4 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X78Y101_A5 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X78Y101_A6 = 1'b1;
  assign CLBLM_R_X59Y100_SLICE_X89Y100_C4 = CLBLM_L_X62Y101_SLICE_X93Y101_BQ;
  assign CLBLL_L_X52Y101_SLICE_X78Y101_B1 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X78Y101_B2 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X78Y101_B3 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X78Y101_B4 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X78Y101_B5 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X78Y101_B6 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X78Y101_C1 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X78Y101_C2 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X78Y101_C3 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X78Y101_C4 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X78Y101_C5 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X78Y101_C6 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X78Y101_D1 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X78Y101_D2 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X78Y101_D3 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X78Y101_D4 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X78Y101_D5 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X78Y101_D6 = 1'b1;
  assign CLBLL_R_X57Y100_SLICE_X86Y100_A2 = CLBLM_R_X59Y98_SLICE_X89Y98_AQ;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_D1 = CLBLL_R_X57Y99_SLICE_X87Y99_AQ;
  assign CLBLL_L_X52Y101_SLICE_X79Y101_A1 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign CLBLL_L_X52Y101_SLICE_X79Y101_A2 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLL_L_X52Y101_SLICE_X79Y101_A3 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLL_L_X52Y101_SLICE_X79Y101_A4 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLL_L_X52Y101_SLICE_X79Y101_A5 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLL_L_X52Y101_SLICE_X79Y101_A6 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLM_R_X59Y100_SLICE_X89Y100_D4 = CLBLM_L_X62Y101_SLICE_X93Y101_CQ;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_T1 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X79Y101_B1 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X79Y101_B2 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X79Y101_B3 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X79Y101_B4 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X79Y101_B5 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X79Y101_B6 = 1'b1;
  assign CLBLL_R_X57Y100_SLICE_X86Y100_A3 = CLBLM_L_X60Y100_SLICE_X90Y100_AO6;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_D1 = CLBLM_L_X60Y111_SLICE_X91Y111_AQ;
  assign CLBLL_L_X52Y101_SLICE_X79Y101_C1 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X79Y101_C2 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X79Y101_C3 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X79Y101_C4 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X79Y101_C5 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X79Y101_C6 = 1'b1;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_T1 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X79Y101_D1 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X79Y101_D2 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X79Y101_D3 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X79Y101_D4 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X79Y101_D5 = 1'b1;
  assign CLBLL_L_X52Y101_SLICE_X79Y101_D6 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X81Y102_A1 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X81Y102_A2 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X81Y102_A3 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X81Y102_A4 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X81Y102_A5 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X81Y102_A6 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X81Y102_B1 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X81Y102_B2 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X81Y102_B3 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X81Y102_B4 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X81Y102_B5 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X81Y102_B6 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X81Y102_C1 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X81Y102_C2 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X81Y102_C3 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X81Y102_C4 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X81Y102_C5 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X81Y102_C6 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X81Y102_D1 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X81Y102_D2 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X81Y102_D3 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X81Y102_D4 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X81Y102_D5 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X81Y102_D6 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X80Y102_A1 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLM_R_X53Y102_SLICE_X80Y102_A2 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLM_R_X53Y102_SLICE_X80Y102_A3 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLM_R_X53Y102_SLICE_X80Y102_A4 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLM_R_X53Y102_SLICE_X80Y102_A5 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign CLBLM_R_X53Y102_SLICE_X80Y102_A6 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLM_R_X53Y102_SLICE_X80Y102_B1 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X80Y102_B2 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X80Y102_B3 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X80Y102_B4 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X80Y102_B5 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X80Y102_B6 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X80Y102_C1 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X80Y102_C2 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X80Y102_C3 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X80Y102_C4 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X80Y102_C5 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X80Y102_C6 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X80Y102_D1 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X80Y102_D2 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X80Y102_D3 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X80Y102_D4 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X80Y102_D5 = 1'b1;
  assign CLBLM_R_X53Y102_SLICE_X80Y102_D6 = 1'b1;
  assign CLBLL_R_X57Y100_SLICE_X86Y100_B1 = CLBLL_L_X54Y99_SLICE_X82Y99_AQ;
  assign CLBLL_R_X57Y100_SLICE_X86Y100_B2 = 1'b1;
  assign CLBLL_R_X57Y100_SLICE_X86Y100_B3 = CLBLL_L_X54Y98_SLICE_X83Y98_BQ;
  assign CLBLM_R_X53Y103_SLICE_X81Y103_A1 = 1'b1;
  assign CLBLM_R_X53Y103_SLICE_X81Y103_A2 = CLBLL_R_X57Y100_SLICE_X86Y100_DQ;
  assign CLBLM_R_X53Y103_SLICE_X81Y103_A3 = 1'b1;
  assign CLBLM_R_X53Y103_SLICE_X81Y103_A4 = 1'b1;
  assign CLBLM_R_X53Y103_SLICE_X81Y103_A5 = 1'b1;
  assign CLBLM_R_X53Y103_SLICE_X81Y103_A6 = CLBLL_R_X57Y100_SLICE_X86Y100_AQ;
  assign CLBLM_R_X53Y103_SLICE_X81Y103_AX = 1'b0;
  assign CLBLM_R_X53Y103_SLICE_X81Y103_B1 = CLBLL_R_X57Y100_SLICE_X86Y100_BQ;
  assign CLBLM_R_X53Y103_SLICE_X81Y103_B2 = CLBLL_R_X57Y100_SLICE_X86Y100_AQ;
  assign CLBLM_R_X53Y103_SLICE_X81Y103_B3 = 1'b1;
  assign CLBLM_R_X53Y103_SLICE_X81Y103_B4 = CLBLL_R_X57Y100_SLICE_X86Y100_DQ;
  assign CLBLM_R_X53Y103_SLICE_X81Y103_B5 = CLBLL_R_X57Y100_SLICE_X86Y100_CQ;
  assign CLBLM_R_X53Y103_SLICE_X81Y103_B6 = 1'b1;
  assign CLBLM_R_X53Y103_SLICE_X81Y103_C1 = CLBLL_R_X57Y100_SLICE_X86Y100_CQ;
  assign CLBLM_R_X53Y103_SLICE_X81Y103_C2 = CLBLL_R_X57Y100_SLICE_X86Y100_DQ;
  assign CLBLM_R_X53Y103_SLICE_X81Y103_C3 = CLBLM_L_X56Y101_SLICE_X85Y101_AQ;
  assign CLBLM_R_X53Y103_SLICE_X81Y103_C4 = CLBLL_R_X57Y100_SLICE_X86Y100_BQ;
  assign CLBLM_R_X53Y103_SLICE_X81Y103_C5 = CLBLL_R_X57Y100_SLICE_X86Y100_AQ;
  assign CLBLM_R_X53Y103_SLICE_X81Y103_C6 = CLBLM_L_X56Y101_SLICE_X85Y101_CQ;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_CX = CLBLM_L_X62Y97_SLICE_X93Y97_CO5;
  assign CLBLM_R_X53Y103_SLICE_X81Y103_CX = CLBLM_R_X53Y103_SLICE_X80Y103_BO6;
  assign CLBLM_R_X53Y103_SLICE_X81Y103_D1 = CLBLL_R_X57Y100_SLICE_X86Y100_CQ;
  assign CLBLM_R_X53Y103_SLICE_X81Y103_D2 = CLBLL_R_X57Y100_SLICE_X87Y100_AQ;
  assign CLBLM_R_X53Y103_SLICE_X81Y103_D3 = CLBLM_L_X56Y101_SLICE_X85Y101_AQ;
  assign CLBLM_R_X53Y103_SLICE_X81Y103_D4 = CLBLL_L_X52Y105_SLICE_X78Y105_BO6;
  assign CLBLM_R_X53Y103_SLICE_X81Y103_D5 = CLBLL_R_X57Y100_SLICE_X86Y100_AQ;
  assign CLBLM_R_X53Y103_SLICE_X81Y103_D6 = CLBLL_R_X57Y100_SLICE_X86Y100_DQ;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_D1 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X53Y103_SLICE_X81Y103_DX = CLBLM_R_X53Y103_SLICE_X80Y103_AO6;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_D2 = CLBLM_R_X63Y99_SLICE_X95Y99_B5Q;
  assign CLBLM_R_X53Y103_SLICE_X80Y103_A1 = CLBLM_L_X56Y101_SLICE_X85Y101_AQ;
  assign CLBLM_R_X53Y103_SLICE_X80Y103_A2 = CLBLM_L_X56Y101_SLICE_X85Y101_CQ;
  assign CLBLM_R_X53Y103_SLICE_X80Y103_A3 = CLBLL_R_X57Y100_SLICE_X86Y100_CQ;
  assign CLBLM_R_X53Y103_SLICE_X80Y103_A4 = CLBLL_R_X57Y100_SLICE_X86Y100_DQ;
  assign CLBLM_R_X53Y103_SLICE_X80Y103_A5 = CLBLL_R_X57Y100_SLICE_X87Y100_AQ;
  assign CLBLM_R_X53Y103_SLICE_X80Y103_A6 = CLBLL_R_X57Y100_SLICE_X86Y100_BQ;
  assign CLBLM_R_X53Y103_SLICE_X80Y103_B1 = CLBLL_R_X57Y100_SLICE_X86Y100_AQ;
  assign CLBLM_R_X53Y103_SLICE_X80Y103_B2 = CLBLM_L_X56Y101_SLICE_X85Y101_CQ;
  assign CLBLM_R_X53Y103_SLICE_X80Y103_B3 = CLBLL_R_X57Y100_SLICE_X86Y100_CQ;
  assign CLBLM_R_X53Y103_SLICE_X80Y103_B4 = CLBLL_R_X57Y100_SLICE_X86Y100_BQ;
  assign CLBLM_R_X53Y103_SLICE_X80Y103_B5 = 1'b1;
  assign CLBLM_R_X53Y103_SLICE_X80Y103_B6 = 1'b1;
  assign CLBLM_R_X53Y103_SLICE_X80Y103_C1 = 1'b1;
  assign CLBLM_R_X53Y103_SLICE_X80Y103_C2 = 1'b1;
  assign CLBLM_R_X53Y103_SLICE_X80Y103_C3 = 1'b1;
  assign CLBLM_R_X53Y103_SLICE_X80Y103_C4 = 1'b1;
  assign CLBLM_R_X53Y103_SLICE_X80Y103_C5 = 1'b1;
  assign CLBLM_R_X53Y103_SLICE_X80Y103_C6 = 1'b1;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_DX = CLBLM_R_X63Y96_SLICE_X95Y96_AO5;
  assign CLBLM_R_X53Y103_SLICE_X80Y103_D1 = 1'b1;
  assign CLBLM_R_X53Y103_SLICE_X80Y103_D2 = 1'b1;
  assign CLBLM_R_X53Y103_SLICE_X80Y103_D3 = 1'b1;
  assign CLBLM_R_X53Y103_SLICE_X80Y103_D4 = 1'b1;
  assign CLBLM_R_X53Y103_SLICE_X80Y103_D5 = 1'b1;
  assign CLBLM_R_X53Y103_SLICE_X80Y103_D6 = 1'b1;
  assign CLBLM_R_X63Y95_SLICE_X94Y95_A1 = CLBLM_L_X62Y95_SLICE_X92Y95_AQ;
  assign CLBLM_R_X63Y95_SLICE_X94Y95_A2 = CLBLM_L_X62Y98_SLICE_X92Y98_CQ;
  assign CLBLM_R_X63Y95_SLICE_X94Y95_A4 = CLBLM_L_X62Y98_SLICE_X92Y98_AQ;
  assign CLBLM_R_X63Y95_SLICE_X94Y95_A5 = CLBLM_L_X62Y95_SLICE_X92Y95_A5Q;
  assign CLBLM_R_X53Y104_SLICE_X81Y104_A1 = CLBLL_R_X57Y101_SLICE_X87Y101_AQ;
  assign CLBLM_R_X53Y104_SLICE_X81Y104_A2 = CLBLM_R_X53Y104_SLICE_X80Y104_DO5;
  assign CLBLM_R_X53Y104_SLICE_X81Y104_A3 = CLBLM_R_X53Y104_SLICE_X80Y104_CO6;
  assign CLBLM_R_X53Y104_SLICE_X81Y104_A4 = CLBLL_R_X57Y100_SLICE_X86Y100_DQ;
  assign CLBLM_R_X53Y104_SLICE_X81Y104_A5 = CLBLL_R_X57Y100_SLICE_X86Y100_CQ;
  assign CLBLM_R_X53Y104_SLICE_X81Y104_A6 = CLBLL_R_X57Y100_SLICE_X87Y100_AQ;
  assign CLBLM_R_X53Y104_SLICE_X81Y104_AX = CLBLM_R_X53Y104_SLICE_X80Y104_CO6;
  assign CLBLM_R_X53Y104_SLICE_X81Y104_B1 = CLBLM_L_X56Y101_SLICE_X85Y101_BQ;
  assign CLBLM_R_X53Y104_SLICE_X81Y104_B2 = CLBLM_R_X53Y104_SLICE_X80Y104_BO6;
  assign CLBLM_R_X53Y104_SLICE_X81Y104_B3 = CLBLM_R_X53Y104_SLICE_X80Y104_AO5;
  assign CLBLM_R_X53Y104_SLICE_X81Y104_B4 = CLBLM_L_X56Y101_SLICE_X85Y101_CQ;
  assign CLBLM_R_X53Y104_SLICE_X81Y104_B5 = CLBLL_R_X57Y100_SLICE_X86Y100_DQ;
  assign CLBLM_R_X53Y104_SLICE_X81Y104_B6 = CLBLL_R_X57Y100_SLICE_X87Y100_AQ;
  assign CLBLM_R_X53Y104_SLICE_X81Y104_BX = CLBLM_R_X53Y104_SLICE_X80Y104_BO6;
  assign CLBLM_R_X53Y104_SLICE_X81Y104_C1 = CLBLL_R_X57Y100_SLICE_X86Y100_DQ;
  assign CLBLM_R_X53Y104_SLICE_X81Y104_C2 = CLBLM_L_X56Y101_SLICE_X85Y101_CQ;
  assign CLBLM_R_X53Y104_SLICE_X81Y104_C3 = CLBLL_R_X57Y101_SLICE_X87Y101_AQ;
  assign CLBLM_R_X53Y104_SLICE_X81Y104_C4 = CLBLL_L_X54Y104_SLICE_X82Y104_AO6;
  assign CLBLM_R_X53Y104_SLICE_X81Y104_C5 = CLBLM_R_X53Y104_SLICE_X80Y104_AO6;
  assign CLBLM_R_X53Y104_SLICE_X81Y104_C6 = CLBLL_R_X57Y100_SLICE_X87Y100_BQ;
  assign CLBLM_R_X53Y104_SLICE_X81Y104_CIN = CLBLM_R_X53Y103_SLICE_X81Y103_COUT;
  assign CLBLM_R_X53Y104_SLICE_X81Y104_CX = CLBLL_L_X54Y104_SLICE_X82Y104_AO6;
  assign CLBLM_R_X53Y104_SLICE_X81Y104_D1 = CLBLL_R_X57Y100_SLICE_X86Y100_DQ;
  assign CLBLM_R_X53Y104_SLICE_X81Y104_D2 = CLBLM_L_X56Y101_SLICE_X85Y101_CQ;
  assign CLBLM_R_X53Y104_SLICE_X81Y104_D3 = CLBLM_R_X53Y104_SLICE_X80Y104_DO6;
  assign CLBLM_R_X53Y104_SLICE_X81Y104_D4 = CLBLM_L_X56Y101_SLICE_X85Y101_BQ;
  assign CLBLM_R_X53Y104_SLICE_X81Y104_D5 = CLBLL_L_X54Y104_SLICE_X82Y104_BO6;
  assign CLBLM_R_X53Y104_SLICE_X81Y104_D6 = CLBLL_R_X57Y99_SLICE_X86Y99_AQ;
  assign CLBLM_R_X53Y104_SLICE_X81Y104_DX = CLBLL_L_X54Y104_SLICE_X82Y104_BO6;
  assign CLBLM_R_X53Y104_SLICE_X80Y104_A1 = CLBLL_R_X57Y101_SLICE_X87Y101_AQ;
  assign CLBLM_R_X53Y104_SLICE_X80Y104_A2 = CLBLM_L_X56Y101_SLICE_X85Y101_BQ;
  assign CLBLM_R_X53Y104_SLICE_X80Y104_A3 = 1'b1;
  assign CLBLM_R_X53Y104_SLICE_X80Y104_A4 = CLBLL_R_X57Y100_SLICE_X86Y100_CQ;
  assign CLBLM_R_X53Y104_SLICE_X80Y104_A5 = 1'b1;
  assign CLBLM_R_X53Y104_SLICE_X80Y104_A6 = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_D1 = CLBLM_L_X62Y110_SLICE_X93Y110_AQ;
  assign CLBLM_R_X53Y104_SLICE_X80Y104_B1 = CLBLL_R_X57Y101_SLICE_X87Y101_AQ;
  assign CLBLM_R_X53Y104_SLICE_X80Y104_B2 = CLBLL_R_X57Y100_SLICE_X86Y100_DQ;
  assign CLBLM_R_X53Y104_SLICE_X80Y104_B3 = CLBLL_R_X57Y100_SLICE_X86Y100_CQ;
  assign CLBLM_R_X53Y104_SLICE_X80Y104_B4 = CLBLM_L_X56Y101_SLICE_X85Y101_CQ;
  assign CLBLM_R_X53Y104_SLICE_X80Y104_B5 = CLBLM_L_X56Y101_SLICE_X85Y101_AQ;
  assign CLBLM_R_X53Y104_SLICE_X80Y104_B6 = CLBLL_R_X57Y100_SLICE_X87Y100_AQ;
  assign CLBLM_R_X63Y94_SLICE_X95Y94_D4 = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_T1 = 1'b1;
  assign CLBLM_R_X53Y104_SLICE_X80Y104_C1 = CLBLM_L_X56Y101_SLICE_X85Y101_AQ;
  assign CLBLM_R_X53Y104_SLICE_X80Y104_C2 = CLBLL_R_X57Y100_SLICE_X87Y100_AQ;
  assign CLBLM_R_X53Y104_SLICE_X80Y104_C3 = CLBLL_R_X57Y100_SLICE_X86Y100_DQ;
  assign CLBLM_R_X53Y104_SLICE_X80Y104_C4 = CLBLL_R_X57Y100_SLICE_X86Y100_CQ;
  assign CLBLM_R_X53Y104_SLICE_X80Y104_C5 = CLBLM_L_X56Y101_SLICE_X85Y101_CQ;
  assign CLBLM_R_X53Y104_SLICE_X80Y104_C6 = CLBLL_R_X57Y100_SLICE_X86Y100_BQ;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_D1 = CLBLM_L_X60Y98_SLICE_X90Y98_BQ;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_T1 = 1'b1;
  assign CLBLM_R_X53Y104_SLICE_X80Y104_D1 = CLBLM_L_X56Y101_SLICE_X85Y101_AQ;
  assign CLBLM_R_X53Y104_SLICE_X80Y104_D2 = 1'b1;
  assign CLBLM_R_X53Y104_SLICE_X80Y104_D3 = CLBLM_L_X56Y101_SLICE_X85Y101_CQ;
  assign CLBLM_R_X53Y104_SLICE_X80Y104_D4 = CLBLL_R_X57Y100_SLICE_X86Y100_CQ;
  assign CLBLM_R_X53Y104_SLICE_X80Y104_D5 = CLBLL_R_X57Y100_SLICE_X87Y100_BQ;
  assign CLBLM_R_X53Y104_SLICE_X80Y104_D6 = 1'b1;
  assign CLBLM_R_X53Y105_SLICE_X81Y105_A1 = CLBLM_L_X56Y101_SLICE_X85Y101_CQ;
  assign CLBLM_R_X53Y105_SLICE_X81Y105_A2 = CLBLL_R_X57Y100_SLICE_X87Y100_BQ;
  assign CLBLM_R_X53Y105_SLICE_X81Y105_A3 = CLBLL_R_X57Y99_SLICE_X86Y99_AQ;
  assign CLBLM_R_X53Y105_SLICE_X81Y105_A4 = CLBLL_R_X57Y100_SLICE_X86Y100_DQ;
  assign CLBLM_R_X53Y105_SLICE_X81Y105_A5 = CLBLL_R_X57Y100_SLICE_X86Y100_CQ;
  assign CLBLM_R_X53Y105_SLICE_X81Y105_A6 = CLBLM_L_X56Y101_SLICE_X85Y101_BQ;
  assign CLBLM_R_X53Y105_SLICE_X81Y105_AX = CLBLM_R_X53Y105_SLICE_X80Y105_BO6;
  assign CLBLM_R_X53Y105_SLICE_X81Y105_B1 = 1'b1;
  assign CLBLM_R_X53Y105_SLICE_X81Y105_B2 = CLBLL_R_X57Y100_SLICE_X87Y100_BQ;
  assign CLBLM_R_X53Y105_SLICE_X81Y105_B3 = CLBLL_R_X57Y99_SLICE_X86Y99_AQ;
  assign CLBLM_R_X53Y105_SLICE_X81Y105_B4 = CLBLL_R_X57Y100_SLICE_X86Y100_CQ;
  assign CLBLM_R_X53Y105_SLICE_X81Y105_B5 = CLBLM_L_X56Y101_SLICE_X85Y101_CQ;
  assign CLBLM_R_X53Y105_SLICE_X81Y105_B6 = 1'b1;
  assign CLBLM_R_X53Y105_SLICE_X81Y105_C1 = 1'b1;
  assign CLBLM_R_X53Y105_SLICE_X81Y105_C2 = 1'b1;
  assign CLBLM_R_X53Y105_SLICE_X81Y105_C3 = 1'b1;
  assign CLBLM_R_X53Y105_SLICE_X81Y105_C4 = 1'b1;
  assign CLBLM_R_X53Y105_SLICE_X81Y105_C5 = 1'b1;
  assign CLBLM_R_X53Y105_SLICE_X81Y105_C6 = 1'b1;
  assign CLBLM_R_X53Y105_SLICE_X81Y105_CIN = CLBLM_R_X53Y104_SLICE_X81Y104_COUT;
  assign CLBLM_R_X53Y105_SLICE_X81Y105_CX = 1'b0;
  assign CLBLM_R_X53Y105_SLICE_X81Y105_D1 = 1'b1;
  assign CLBLM_R_X53Y105_SLICE_X81Y105_D2 = 1'b1;
  assign CLBLM_R_X53Y105_SLICE_X81Y105_D3 = 1'b1;
  assign CLBLM_R_X53Y105_SLICE_X81Y105_D4 = 1'b1;
  assign CLBLM_R_X53Y105_SLICE_X81Y105_D5 = 1'b1;
  assign CLBLM_R_X53Y105_SLICE_X81Y105_D6 = 1'b1;
  assign CLBLM_R_X53Y105_SLICE_X81Y105_DX = 1'b0;
  assign CLBLM_R_X53Y105_SLICE_X80Y105_A1 = CLBLM_L_X56Y101_SLICE_X85Y101_AQ;
  assign CLBLM_R_X53Y105_SLICE_X80Y105_A2 = CLBLM_R_X53Y106_SLICE_X81Y106_D_XOR;
  assign CLBLM_R_X53Y105_SLICE_X80Y105_A3 = CLBLM_R_X53Y106_SLICE_X80Y106_AO5;
  assign CLBLM_R_X53Y105_SLICE_X80Y105_A4 = CLBLL_R_X57Y101_SLICE_X87Y101_DQ;
  assign CLBLM_R_X53Y105_SLICE_X80Y105_A5 = CLBLM_R_X53Y104_SLICE_X81Y104_C_XOR;
  assign CLBLM_R_X53Y105_SLICE_X80Y105_A6 = CLBLL_R_X57Y100_SLICE_X86Y100_BQ;
  assign CLBLM_R_X53Y105_SLICE_X80Y105_B1 = CLBLM_L_X56Y101_SLICE_X85Y101_CQ;
  assign CLBLM_R_X53Y105_SLICE_X80Y105_B2 = CLBLL_R_X57Y100_SLICE_X86Y100_DQ;
  assign CLBLM_R_X53Y105_SLICE_X80Y105_B3 = CLBLL_R_X57Y100_SLICE_X86Y100_CQ;
  assign CLBLM_R_X53Y105_SLICE_X80Y105_B4 = CLBLM_L_X56Y101_SLICE_X85Y101_BQ;
  assign CLBLM_R_X53Y105_SLICE_X80Y105_B5 = CLBLL_R_X57Y99_SLICE_X86Y99_AQ;
  assign CLBLM_R_X53Y105_SLICE_X80Y105_B6 = CLBLL_R_X57Y100_SLICE_X87Y100_BQ;
  assign CLBLM_R_X53Y105_SLICE_X80Y105_C1 = 1'b1;
  assign CLBLM_R_X53Y105_SLICE_X80Y105_C2 = 1'b1;
  assign CLBLM_R_X53Y105_SLICE_X80Y105_C3 = 1'b1;
  assign CLBLM_R_X53Y105_SLICE_X80Y105_C4 = 1'b1;
  assign CLBLM_R_X53Y105_SLICE_X80Y105_C5 = 1'b1;
  assign CLBLM_R_X53Y105_SLICE_X80Y105_C6 = 1'b1;
  assign CLBLM_R_X53Y105_SLICE_X80Y105_D1 = 1'b1;
  assign CLBLM_R_X53Y105_SLICE_X80Y105_D2 = 1'b1;
  assign CLBLM_R_X53Y105_SLICE_X80Y105_D3 = 1'b1;
  assign CLBLM_R_X53Y105_SLICE_X80Y105_D4 = 1'b1;
  assign CLBLM_R_X53Y105_SLICE_X80Y105_D5 = 1'b1;
  assign CLBLM_R_X53Y105_SLICE_X80Y105_D6 = 1'b1;
  assign CLBLM_L_X64Y95_SLICE_X97Y95_D1 = 1'b1;
  assign CLBLM_L_X64Y95_SLICE_X97Y95_D3 = 1'b1;
  assign CLBLL_L_X52Y105_SLICE_X78Y105_A1 = CLBLM_R_X53Y100_SLICE_X81Y100_AQ;
  assign CLBLL_L_X52Y105_SLICE_X78Y105_A2 = CLBLL_R_X57Y100_SLICE_X86Y100_DQ;
  assign CLBLL_L_X52Y105_SLICE_X78Y105_A3 = CLBLM_R_X53Y101_SLICE_X80Y101_BQ;
  assign CLBLL_L_X52Y105_SLICE_X78Y105_A4 = CLBLL_R_X57Y99_SLICE_X86Y99_BQ;
  assign CLBLL_L_X52Y105_SLICE_X78Y105_A5 = CLBLL_L_X54Y100_SLICE_X82Y100_BQ;
  assign CLBLL_L_X52Y105_SLICE_X78Y105_A6 = 1'b1;
  assign CLBLL_L_X52Y105_SLICE_X78Y105_B1 = CLBLL_R_X57Y100_SLICE_X86Y100_BQ;
  assign CLBLL_L_X52Y105_SLICE_X78Y105_B2 = 1'b1;
  assign CLBLL_L_X52Y105_SLICE_X78Y105_B3 = CLBLL_R_X57Y100_SLICE_X86Y100_DQ;
  assign CLBLL_L_X52Y105_SLICE_X78Y105_B4 = CLBLM_L_X56Y101_SLICE_X85Y101_CQ;
  assign CLBLL_L_X52Y105_SLICE_X78Y105_B5 = CLBLL_L_X54Y100_SLICE_X82Y100_BQ;
  assign CLBLL_L_X52Y105_SLICE_X78Y105_B6 = 1'b1;
  assign CLBLL_L_X52Y105_SLICE_X78Y105_C1 = CLBLM_R_X53Y101_SLICE_X80Y101_BQ;
  assign CLBLL_L_X52Y105_SLICE_X78Y105_C2 = CLBLL_L_X52Y106_SLICE_X78Y106_AO5;
  assign CLBLL_L_X52Y105_SLICE_X78Y105_C3 = CLBLL_R_X57Y97_SLICE_X86Y97_AQ;
  assign CLBLL_L_X52Y105_SLICE_X78Y105_C4 = CLBLL_L_X52Y105_SLICE_X78Y105_AO5;
  assign CLBLL_L_X52Y105_SLICE_X78Y105_C5 = CLBLM_R_X53Y101_SLICE_X81Y101_AQ;
  assign CLBLL_L_X52Y105_SLICE_X78Y105_C6 = CLBLL_R_X57Y99_SLICE_X86Y99_BQ;
  assign CLBLL_L_X52Y105_SLICE_X78Y105_D1 = 1'b1;
  assign CLBLL_L_X52Y105_SLICE_X78Y105_D2 = 1'b1;
  assign CLBLL_L_X52Y105_SLICE_X78Y105_D3 = 1'b1;
  assign CLBLL_L_X52Y105_SLICE_X78Y105_D4 = 1'b1;
  assign CLBLL_L_X52Y105_SLICE_X78Y105_D5 = 1'b1;
  assign CLBLL_L_X52Y105_SLICE_X78Y105_D6 = 1'b1;
  assign CLBLL_L_X52Y105_SLICE_X79Y105_A1 = 1'b1;
  assign CLBLL_L_X52Y105_SLICE_X79Y105_A2 = 1'b1;
  assign CLBLL_L_X52Y105_SLICE_X79Y105_A3 = 1'b1;
  assign CLBLL_L_X52Y105_SLICE_X79Y105_A4 = 1'b1;
  assign CLBLL_L_X52Y105_SLICE_X79Y105_A5 = 1'b1;
  assign CLBLL_L_X52Y105_SLICE_X79Y105_A6 = 1'b1;
  assign CLBLL_L_X52Y105_SLICE_X79Y105_B1 = 1'b1;
  assign CLBLL_L_X52Y105_SLICE_X79Y105_B2 = 1'b1;
  assign CLBLL_L_X52Y105_SLICE_X79Y105_B3 = 1'b1;
  assign CLBLL_L_X52Y105_SLICE_X79Y105_B4 = 1'b1;
  assign CLBLL_L_X52Y105_SLICE_X79Y105_B5 = 1'b1;
  assign CLBLL_L_X52Y105_SLICE_X79Y105_B6 = 1'b1;
  assign CLBLL_L_X52Y105_SLICE_X79Y105_C1 = 1'b1;
  assign CLBLL_L_X52Y105_SLICE_X79Y105_C2 = 1'b1;
  assign CLBLL_L_X52Y105_SLICE_X79Y105_C3 = 1'b1;
  assign CLBLL_L_X52Y105_SLICE_X79Y105_C4 = 1'b1;
  assign CLBLL_L_X52Y105_SLICE_X79Y105_C5 = 1'b1;
  assign CLBLL_L_X52Y105_SLICE_X79Y105_C6 = 1'b1;
  assign CLBLL_L_X52Y105_SLICE_X79Y105_D1 = 1'b1;
  assign CLBLL_L_X52Y105_SLICE_X79Y105_D2 = 1'b1;
  assign CLBLL_L_X52Y105_SLICE_X79Y105_D3 = 1'b1;
  assign CLBLL_L_X52Y105_SLICE_X79Y105_D4 = 1'b1;
  assign CLBLL_L_X52Y105_SLICE_X79Y105_D5 = 1'b1;
  assign CLBLL_L_X52Y105_SLICE_X79Y105_D6 = 1'b1;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_B1 = CLBLM_L_X62Y95_SLICE_X92Y95_AQ;
  assign CLBLM_R_X53Y106_SLICE_X81Y106_A1 = 1'b1;
  assign CLBLM_R_X53Y106_SLICE_X81Y106_A2 = CLBLL_R_X57Y100_SLICE_X87Y100_CQ;
  assign CLBLM_R_X53Y106_SLICE_X81Y106_A3 = CLBLL_R_X57Y100_SLICE_X86Y100_AQ;
  assign CLBLM_R_X53Y106_SLICE_X81Y106_A4 = 1'b1;
  assign CLBLM_R_X53Y106_SLICE_X81Y106_A5 = 1'b1;
  assign CLBLM_R_X53Y106_SLICE_X81Y106_A6 = 1'b1;
  assign CLBLM_R_X53Y106_SLICE_X81Y106_AX = 1'b0;
  assign CLBLM_R_X53Y106_SLICE_X81Y106_B1 = 1'b1;
  assign CLBLM_R_X53Y106_SLICE_X81Y106_B2 = CLBLL_R_X57Y100_SLICE_X87Y100_CQ;
  assign CLBLM_R_X53Y106_SLICE_X81Y106_B3 = CLBLL_R_X57Y100_SLICE_X86Y100_AQ;
  assign CLBLM_R_X53Y106_SLICE_X81Y106_B4 = CLBLL_R_X57Y101_SLICE_X87Y101_CQ;
  assign CLBLM_R_X53Y106_SLICE_X81Y106_B5 = CLBLL_R_X57Y100_SLICE_X86Y100_BQ;
  assign CLBLM_R_X53Y106_SLICE_X81Y106_B6 = 1'b1;
  assign CLBLM_R_X53Y106_SLICE_X81Y106_C1 = CLBLL_R_X57Y100_SLICE_X86Y100_BQ;
  assign CLBLM_R_X53Y106_SLICE_X81Y106_C2 = CLBLL_R_X57Y100_SLICE_X87Y100_CQ;
  assign CLBLM_R_X53Y106_SLICE_X81Y106_C3 = CLBLL_R_X57Y101_SLICE_X87Y101_CQ;
  assign CLBLM_R_X53Y106_SLICE_X81Y106_C4 = CLBLM_L_X56Y101_SLICE_X85Y101_DQ;
  assign CLBLM_R_X53Y106_SLICE_X81Y106_C5 = CLBLL_R_X57Y100_SLICE_X86Y100_AQ;
  assign CLBLM_R_X53Y106_SLICE_X81Y106_C6 = CLBLM_L_X56Y101_SLICE_X85Y101_AQ;
  assign CLBLM_R_X53Y106_SLICE_X81Y106_CX = CLBLL_L_X52Y106_SLICE_X79Y106_BO6;
  assign CLBLM_R_X53Y106_SLICE_X81Y106_D1 = CLBLL_R_X57Y100_SLICE_X87Y100_CQ;
  assign CLBLM_R_X53Y106_SLICE_X81Y106_D2 = CLBLL_R_X57Y100_SLICE_X87Y100_AQ;
  assign CLBLM_R_X53Y106_SLICE_X81Y106_D3 = CLBLM_R_X53Y106_SLICE_X80Y106_DO6;
  assign CLBLM_R_X53Y106_SLICE_X81Y106_D4 = CLBLL_R_X57Y100_SLICE_X86Y100_AQ;
  assign CLBLM_R_X53Y106_SLICE_X81Y106_D5 = CLBLL_R_X57Y101_SLICE_X87Y101_CQ;
  assign CLBLM_R_X53Y106_SLICE_X81Y106_D6 = CLBLM_L_X56Y101_SLICE_X85Y101_AQ;
  assign CLBLM_R_X53Y106_SLICE_X81Y106_DX = CLBLM_R_X53Y106_SLICE_X80Y106_CO6;
  assign CLBLM_R_X53Y106_SLICE_X80Y106_A1 = CLBLM_R_X53Y107_SLICE_X81Y107_B_XOR;
  assign CLBLM_R_X53Y106_SLICE_X80Y106_A2 = CLBLM_R_X53Y105_SLICE_X81Y105_A_XOR;
  assign CLBLM_R_X53Y106_SLICE_X80Y106_A3 = CLBLL_R_X57Y100_SLICE_X86Y100_BQ;
  assign CLBLM_R_X53Y106_SLICE_X80Y106_A4 = CLBLL_R_X57Y99_SLICE_X86Y99_BQ;
  assign CLBLM_R_X53Y106_SLICE_X80Y106_A5 = 1'b1;
  assign CLBLM_R_X53Y106_SLICE_X80Y106_A6 = 1'b1;
  assign CLBLM_R_X53Y106_SLICE_X80Y106_B1 = CLBLL_R_X57Y100_SLICE_X86Y100_BQ;
  assign CLBLM_R_X53Y106_SLICE_X80Y106_B2 = CLBLM_R_X53Y106_SLICE_X81Y106_D_XOR;
  assign CLBLM_R_X53Y106_SLICE_X80Y106_B3 = CLBLM_R_X53Y104_SLICE_X81Y104_C_XOR;
  assign CLBLM_R_X53Y106_SLICE_X80Y106_B4 = CLBLL_R_X57Y101_SLICE_X87Y101_DQ;
  assign CLBLM_R_X53Y106_SLICE_X80Y106_B5 = CLBLM_L_X56Y101_SLICE_X85Y101_AQ;
  assign CLBLM_R_X53Y106_SLICE_X80Y106_B6 = CLBLM_R_X53Y106_SLICE_X80Y106_AO5;
  assign CLBLM_R_X53Y106_SLICE_X80Y106_C1 = CLBLL_R_X57Y100_SLICE_X86Y100_BQ;
  assign CLBLM_R_X53Y106_SLICE_X80Y106_C2 = CLBLM_L_X56Y101_SLICE_X85Y101_DQ;
  assign CLBLM_R_X53Y106_SLICE_X80Y106_C3 = CLBLL_R_X57Y100_SLICE_X87Y100_AQ;
  assign CLBLM_R_X53Y106_SLICE_X80Y106_C4 = CLBLL_R_X57Y100_SLICE_X87Y100_CQ;
  assign CLBLM_R_X53Y106_SLICE_X80Y106_C5 = CLBLL_R_X57Y101_SLICE_X87Y101_CQ;
  assign CLBLM_R_X53Y106_SLICE_X80Y106_C6 = CLBLM_L_X56Y101_SLICE_X85Y101_AQ;
  assign CLBLM_R_X53Y106_SLICE_X80Y106_D1 = CLBLL_R_X57Y100_SLICE_X86Y100_BQ;
  assign CLBLM_R_X53Y106_SLICE_X80Y106_D2 = 1'b1;
  assign CLBLM_R_X53Y106_SLICE_X80Y106_D3 = 1'b1;
  assign CLBLM_R_X53Y106_SLICE_X80Y106_D4 = CLBLM_L_X56Y101_SLICE_X85Y101_DQ;
  assign CLBLM_R_X53Y106_SLICE_X80Y106_D5 = 1'b1;
  assign CLBLM_R_X53Y106_SLICE_X80Y106_D6 = 1'b1;
  assign CLBLM_R_X59Y101_SLICE_X89Y101_B4 = CLBLM_R_X59Y103_SLICE_X89Y103_DQ;
  assign CLBLM_R_X59Y101_SLICE_X89Y101_B5 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLL_L_X52Y106_SLICE_X78Y106_A1 = CLBLM_L_X50Y106_SLICE_X76Y106_BO5;
  assign CLBLL_L_X52Y106_SLICE_X78Y106_A2 = 1'b1;
  assign CLBLL_L_X52Y106_SLICE_X78Y106_A3 = CLBLL_R_X57Y101_SLICE_X87Y101_DQ;
  assign CLBLL_L_X52Y106_SLICE_X78Y106_A4 = CLBLM_L_X56Y101_SLICE_X85Y101_DQ;
  assign CLBLL_L_X52Y106_SLICE_X78Y106_A5 = CLBLL_R_X57Y99_SLICE_X86Y99_AQ;
  assign CLBLL_L_X52Y106_SLICE_X78Y106_A6 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_A1 = 1'b1;
  assign CLBLL_L_X52Y106_SLICE_X78Y106_B1 = 1'b1;
  assign CLBLL_L_X52Y106_SLICE_X78Y106_B2 = 1'b1;
  assign CLBLL_L_X52Y106_SLICE_X78Y106_B3 = 1'b1;
  assign CLBLL_L_X52Y106_SLICE_X78Y106_B4 = 1'b1;
  assign CLBLL_L_X52Y106_SLICE_X78Y106_B5 = 1'b1;
  assign CLBLL_L_X52Y106_SLICE_X78Y106_B6 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_A2 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_A3 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_A4 = 1'b1;
  assign CLBLL_L_X52Y106_SLICE_X78Y106_C1 = 1'b1;
  assign CLBLL_L_X52Y106_SLICE_X78Y106_C2 = 1'b1;
  assign CLBLL_L_X52Y106_SLICE_X78Y106_C3 = 1'b1;
  assign CLBLL_L_X52Y106_SLICE_X78Y106_C4 = 1'b1;
  assign CLBLL_L_X52Y106_SLICE_X78Y106_C5 = 1'b1;
  assign CLBLL_L_X52Y106_SLICE_X78Y106_C6 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_B1 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_B2 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_B3 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_B4 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_B5 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_B6 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_C1 = 1'b1;
  assign CLBLL_L_X52Y106_SLICE_X78Y106_D1 = 1'b1;
  assign CLBLL_L_X52Y106_SLICE_X78Y106_D2 = 1'b1;
  assign CLBLL_L_X52Y106_SLICE_X78Y106_D3 = 1'b1;
  assign CLBLL_L_X52Y106_SLICE_X78Y106_D4 = 1'b1;
  assign CLBLL_L_X52Y106_SLICE_X78Y106_D5 = 1'b1;
  assign CLBLL_L_X52Y106_SLICE_X78Y106_D6 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_C5 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_C6 = 1'b1;
  assign CLBLM_L_X64Y95_SLICE_X97Y95_A1 = 1'b1;
  assign CLBLM_L_X64Y95_SLICE_X97Y95_A2 = 1'b1;
  assign CLBLM_L_X64Y95_SLICE_X97Y95_A3 = 1'b1;
  assign CLBLM_L_X64Y95_SLICE_X97Y95_A4 = 1'b1;
  assign CLBLM_L_X64Y95_SLICE_X97Y95_A5 = 1'b1;
  assign CLBLM_L_X64Y95_SLICE_X97Y95_A6 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_D1 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_D2 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_D3 = 1'b1;
  assign CLBLM_L_X64Y95_SLICE_X97Y95_B1 = 1'b1;
  assign CLBLM_L_X64Y95_SLICE_X97Y95_B2 = 1'b1;
  assign CLBLM_L_X64Y95_SLICE_X97Y95_B3 = 1'b1;
  assign CLBLM_L_X64Y95_SLICE_X97Y95_B4 = 1'b1;
  assign CLBLM_L_X64Y95_SLICE_X97Y95_B5 = 1'b1;
  assign CLBLM_L_X64Y95_SLICE_X97Y95_B6 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_A1 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_A2 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_A3 = 1'b1;
  assign CLBLM_L_X64Y95_SLICE_X97Y95_C1 = 1'b1;
  assign CLBLM_L_X64Y95_SLICE_X97Y95_C2 = 1'b1;
  assign CLBLM_L_X64Y95_SLICE_X97Y95_C3 = 1'b1;
  assign CLBLM_L_X64Y95_SLICE_X97Y95_C4 = 1'b1;
  assign CLBLM_L_X64Y95_SLICE_X97Y95_C5 = 1'b1;
  assign CLBLL_L_X52Y106_SLICE_X79Y106_A1 = CLBLL_R_X57Y101_SLICE_X87Y101_CQ;
  assign CLBLL_L_X52Y106_SLICE_X79Y106_A2 = CLBLL_L_X54Y100_SLICE_X82Y100_BQ;
  assign CLBLL_L_X52Y106_SLICE_X79Y106_A3 = CLBLL_R_X57Y101_SLICE_X87Y101_AQ;
  assign CLBLL_L_X52Y106_SLICE_X79Y106_A4 = CLBLL_R_X57Y100_SLICE_X86Y100_DQ;
  assign CLBLL_L_X52Y106_SLICE_X79Y106_A5 = CLBLM_R_X53Y101_SLICE_X80Y101_BQ;
  assign CLBLL_L_X52Y106_SLICE_X79Y106_A6 = 1'b1;
  assign CLBLM_L_X64Y95_SLICE_X97Y95_C6 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_B2 = 1'b1;
  assign CLBLL_L_X52Y106_SLICE_X79Y106_B1 = CLBLL_R_X57Y101_SLICE_X87Y101_CQ;
  assign CLBLL_L_X52Y106_SLICE_X79Y106_B2 = 1'b1;
  assign CLBLL_L_X52Y106_SLICE_X79Y106_B3 = 1'b1;
  assign CLBLM_L_X64Y95_SLICE_X97Y95_D4 = 1'b1;
  assign CLBLM_L_X64Y95_SLICE_X97Y95_D5 = 1'b1;
  assign CLBLM_L_X64Y95_SLICE_X97Y95_D6 = 1'b1;
  assign CLBLL_L_X52Y106_SLICE_X79Y106_B4 = CLBLM_L_X56Y101_SLICE_X85Y101_DQ;
  assign CLBLL_L_X52Y106_SLICE_X79Y106_B5 = CLBLL_R_X57Y100_SLICE_X86Y100_AQ;
  assign CLBLL_L_X52Y106_SLICE_X79Y106_B6 = CLBLL_R_X57Y100_SLICE_X86Y100_BQ;
  assign CLBLM_L_X64Y95_SLICE_X97Y95_D2 = 1'b1;
  assign CLBLL_L_X52Y106_SLICE_X79Y106_C1 = 1'b1;
  assign CLBLL_L_X52Y106_SLICE_X79Y106_C2 = 1'b1;
  assign CLBLL_L_X52Y106_SLICE_X79Y106_C3 = 1'b1;
  assign CLBLL_L_X52Y106_SLICE_X79Y106_C4 = 1'b1;
  assign CLBLL_L_X52Y106_SLICE_X79Y106_C5 = 1'b1;
  assign CLBLL_L_X52Y106_SLICE_X79Y106_C6 = 1'b1;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_A1 = CLBLM_L_X62Y95_SLICE_X92Y95_AQ;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_AI = CLBLM_R_X63Y94_SLICE_X95Y94_AQ;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_A2 = CLBLM_L_X62Y98_SLICE_X92Y98_CQ;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_A3 = CLBLM_L_X62Y98_SLICE_X92Y98_DQ;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_AX = CLBLM_R_X63Y95_SLICE_X95Y95_DQ;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_A4 = CLBLM_L_X62Y98_SLICE_X92Y98_AQ;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_A5 = CLBLM_L_X62Y95_SLICE_X92Y95_A5Q;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_B2 = CLBLM_L_X62Y98_SLICE_X92Y98_CQ;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_A6 = 1'b1;
  assign CLBLL_L_X52Y106_SLICE_X79Y106_D1 = 1'b1;
  assign CLBLL_L_X52Y106_SLICE_X79Y106_D2 = 1'b1;
  assign CLBLL_L_X52Y106_SLICE_X79Y106_D3 = 1'b1;
  assign CLBLL_L_X52Y106_SLICE_X79Y106_D4 = 1'b1;
  assign CLBLL_L_X52Y106_SLICE_X79Y106_D5 = 1'b1;
  assign CLBLL_L_X52Y106_SLICE_X79Y106_D6 = 1'b1;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_B3 = CLBLM_L_X62Y98_SLICE_X92Y98_DQ;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_B4 = CLBLM_L_X62Y98_SLICE_X92Y98_AQ;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_B5 = CLBLM_L_X62Y95_SLICE_X92Y95_A5Q;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_B6 = 1'b1;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_BI = CLBLM_R_X63Y95_SLICE_X95Y95_BQ;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_BX = CLBLM_R_X63Y95_SLICE_X95Y95_CQ;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_C1 = CLBLM_L_X62Y95_SLICE_X92Y95_AQ;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_C2 = CLBLM_L_X62Y98_SLICE_X92Y98_CQ;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_C3 = CLBLM_L_X62Y98_SLICE_X92Y98_DQ;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_C4 = CLBLM_L_X62Y98_SLICE_X92Y98_AQ;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_C5 = CLBLM_L_X62Y95_SLICE_X92Y95_A5Q;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_C6 = 1'b1;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_CE = CLBLM_L_X60Y98_SLICE_X91Y98_BQ;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_CI = CLBLM_R_X63Y95_SLICE_X95Y95_AQ;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_CX = CLBLM_R_X63Y95_SLICE_X95Y95_B5Q;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_D1 = CLBLM_L_X62Y95_SLICE_X93Y95_DQ;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_D2 = CLBLM_L_X62Y95_SLICE_X93Y95_D5Q;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_D3 = CLBLM_L_X62Y95_SLICE_X93Y95_AQ;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_D4 = CLBLM_L_X62Y95_SLICE_X93Y95_BQ;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_D5 = CLBLM_L_X62Y95_SLICE_X93Y95_CQ;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_D6 = 1'b1;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_DI = 1'b0;
  assign CLBLM_L_X56Y111_SLICE_X84Y111_B6 = 1'b1;
  assign CLBLM_L_X64Y95_SLICE_X96Y95_DX = 1'b0;
  assign CLBLM_R_X53Y107_SLICE_X81Y107_A1 = CLBLL_R_X57Y101_SLICE_X87Y101_AQ;
  assign CLBLM_R_X53Y107_SLICE_X81Y107_A2 = CLBLM_L_X56Y101_SLICE_X85Y101_DQ;
  assign CLBLM_R_X53Y107_SLICE_X81Y107_A3 = CLBLM_R_X53Y107_SLICE_X80Y107_AO5;
  assign CLBLM_R_X53Y107_SLICE_X81Y107_A4 = CLBLL_R_X57Y100_SLICE_X87Y100_CQ;
  assign CLBLM_R_X53Y107_SLICE_X81Y107_A5 = CLBLM_L_X56Y101_SLICE_X85Y101_AQ;
  assign CLBLM_R_X53Y107_SLICE_X81Y107_A6 = CLBLM_R_X53Y108_SLICE_X80Y108_BO6;
  assign CLBLM_R_X53Y107_SLICE_X81Y107_AX = CLBLM_R_X53Y108_SLICE_X80Y108_BO6;
  assign CLBLM_R_X53Y107_SLICE_X81Y107_B1 = CLBLM_L_X56Y101_SLICE_X85Y101_BQ;
  assign CLBLM_R_X53Y107_SLICE_X81Y107_B2 = CLBLM_R_X53Y108_SLICE_X80Y108_AO6;
  assign CLBLM_R_X53Y107_SLICE_X81Y107_B3 = CLBLL_L_X52Y106_SLICE_X79Y106_AO6;
  assign CLBLM_R_X53Y107_SLICE_X81Y107_B4 = CLBLM_L_X56Y101_SLICE_X85Y101_DQ;
  assign CLBLM_R_X53Y107_SLICE_X81Y107_B5 = CLBLL_R_X57Y100_SLICE_X87Y100_AQ;
  assign CLBLM_R_X53Y107_SLICE_X81Y107_B6 = CLBLL_R_X57Y100_SLICE_X87Y100_CQ;
  assign CLBLM_R_X53Y107_SLICE_X81Y107_BX = CLBLM_R_X53Y108_SLICE_X80Y108_AO6;
  assign CLBLM_R_X53Y107_SLICE_X81Y107_C1 = CLBLL_R_X57Y100_SLICE_X87Y100_CQ;
  assign CLBLM_R_X53Y107_SLICE_X81Y107_C2 = CLBLM_L_X56Y101_SLICE_X85Y101_DQ;
  assign CLBLM_R_X53Y107_SLICE_X81Y107_C3 = CLBLL_R_X57Y101_SLICE_X87Y101_AQ;
  assign CLBLM_R_X53Y107_SLICE_X81Y107_C4 = CLBLM_R_X53Y107_SLICE_X80Y107_DO6;
  assign CLBLM_R_X53Y107_SLICE_X81Y107_C5 = CLBLM_R_X53Y107_SLICE_X80Y107_AO6;
  assign CLBLM_R_X53Y107_SLICE_X81Y107_C6 = CLBLL_R_X57Y100_SLICE_X87Y100_BQ;
  assign CLBLM_L_X56Y111_SLICE_X84Y111_C5 = 1'b1;
  assign CLBLM_R_X53Y107_SLICE_X81Y107_CIN = CLBLM_R_X53Y106_SLICE_X81Y106_COUT;
  assign RIOI3_X105Y123_OLOGIC_X1Y123_D1 = CLBLM_R_X63Y103_SLICE_X95Y103_AQ;
  assign CLBLM_R_X53Y107_SLICE_X81Y107_CX = CLBLM_R_X53Y107_SLICE_X80Y107_DO6;
  assign CLBLM_R_X53Y107_SLICE_X81Y107_D1 = CLBLL_R_X57Y100_SLICE_X87Y100_CQ;
  assign CLBLM_R_X53Y107_SLICE_X81Y107_D2 = CLBLL_R_X57Y101_SLICE_X87Y101_CQ;
  assign CLBLM_R_X53Y107_SLICE_X81Y107_D3 = CLBLM_R_X53Y107_SLICE_X80Y107_CO6;
  assign CLBLM_R_X53Y107_SLICE_X81Y107_D4 = CLBLL_R_X57Y100_SLICE_X87Y100_BQ;
  assign CLBLM_R_X53Y107_SLICE_X81Y107_D5 = CLBLL_R_X57Y99_SLICE_X86Y99_AQ;
  assign CLBLM_R_X53Y107_SLICE_X81Y107_D6 = CLBLL_L_X52Y107_SLICE_X78Y107_AO6;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_D = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_D = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X53Y107_SLICE_X81Y107_DX = CLBLM_R_X53Y107_SLICE_X80Y107_CO6;
  assign CLBLM_R_X53Y107_SLICE_X80Y107_A1 = 1'b1;
  assign CLBLM_R_X53Y107_SLICE_X80Y107_A2 = 1'b1;
  assign CLBLM_R_X53Y107_SLICE_X80Y107_A3 = CLBLL_R_X57Y100_SLICE_X87Y100_AQ;
  assign CLBLM_R_X53Y107_SLICE_X80Y107_A4 = CLBLM_L_X56Y101_SLICE_X85Y101_BQ;
  assign CLBLM_R_X53Y107_SLICE_X80Y107_A5 = CLBLL_R_X57Y101_SLICE_X87Y101_CQ;
  assign CLBLM_R_X53Y107_SLICE_X80Y107_A6 = 1'b1;
  assign CLBLM_R_X53Y107_SLICE_X80Y107_B1 = CLBLL_R_X57Y100_SLICE_X87Y100_AQ;
  assign CLBLM_R_X53Y107_SLICE_X80Y107_B2 = CLBLM_R_X53Y107_SLICE_X81Y107_D_XOR;
  assign CLBLM_R_X53Y107_SLICE_X80Y107_B3 = CLBLL_R_X57Y99_SLICE_X86Y99_BQ;
  assign CLBLM_R_X53Y107_SLICE_X80Y107_B4 = 1'b1;
  assign CLBLM_R_X53Y107_SLICE_X80Y107_B5 = CLBLM_R_X53Y105_SLICE_X81Y105_C_CY;
  assign CLBLM_R_X53Y107_SLICE_X80Y107_B6 = 1'b1;
  assign CLBLM_R_X53Y107_SLICE_X80Y107_C1 = CLBLL_R_X57Y100_SLICE_X87Y100_BQ;
  assign CLBLM_R_X53Y107_SLICE_X80Y107_C2 = CLBLL_R_X57Y100_SLICE_X87Y100_CQ;
  assign CLBLM_R_X53Y107_SLICE_X80Y107_C3 = CLBLL_R_X57Y101_SLICE_X87Y101_AQ;
  assign CLBLM_R_X53Y107_SLICE_X80Y107_C4 = CLBLM_L_X56Y101_SLICE_X85Y101_BQ;
  assign CLBLM_R_X53Y107_SLICE_X80Y107_C5 = CLBLM_L_X56Y101_SLICE_X85Y101_DQ;
  assign CLBLM_R_X53Y107_SLICE_X80Y107_C6 = CLBLL_R_X57Y101_SLICE_X87Y101_CQ;
  assign CLBLM_L_X56Y111_SLICE_X84Y111_D1 = 1'b1;
  assign CLBLM_R_X53Y107_SLICE_X80Y107_D1 = CLBLL_R_X57Y100_SLICE_X87Y100_AQ;
  assign CLBLM_R_X53Y107_SLICE_X80Y107_D2 = CLBLL_R_X57Y100_SLICE_X87Y100_CQ;
  assign CLBLM_R_X53Y107_SLICE_X80Y107_D3 = CLBLL_R_X57Y101_SLICE_X87Y101_AQ;
  assign CLBLM_R_X53Y107_SLICE_X80Y107_D4 = CLBLL_R_X57Y101_SLICE_X87Y101_CQ;
  assign CLBLM_R_X53Y107_SLICE_X80Y107_D5 = CLBLM_L_X56Y101_SLICE_X85Y101_DQ;
  assign CLBLM_R_X53Y107_SLICE_X80Y107_D6 = CLBLM_L_X56Y101_SLICE_X85Y101_BQ;
  assign RIOI3_X105Y123_OLOGIC_X1Y123_T1 = 1'b1;
  assign CLBLM_L_X56Y111_SLICE_X84Y111_D3 = 1'b1;
  assign CLBLM_L_X56Y111_SLICE_X84Y111_D4 = 1'b1;
  assign CLBLL_L_X52Y107_SLICE_X78Y107_A1 = CLBLM_L_X56Y101_SLICE_X85Y101_DQ;
  assign CLBLL_L_X52Y107_SLICE_X78Y107_A2 = CLBLL_L_X54Y100_SLICE_X82Y100_BQ;
  assign CLBLL_L_X52Y107_SLICE_X78Y107_A3 = CLBLM_R_X53Y101_SLICE_X80Y101_BQ;
  assign CLBLL_L_X52Y107_SLICE_X78Y107_A4 = CLBLM_L_X56Y101_SLICE_X85Y101_BQ;
  assign CLBLL_L_X52Y107_SLICE_X78Y107_A5 = CLBLL_R_X57Y100_SLICE_X86Y100_CQ;
  assign CLBLL_L_X52Y107_SLICE_X78Y107_A6 = 1'b1;
  assign CLBLL_L_X52Y107_SLICE_X78Y107_B1 = CLBLM_L_X56Y101_SLICE_X85Y101_CQ;
  assign CLBLL_L_X52Y107_SLICE_X78Y107_B2 = CLBLL_R_X57Y100_SLICE_X87Y100_BQ;
  assign CLBLL_L_X52Y107_SLICE_X78Y107_B3 = CLBLM_R_X53Y101_SLICE_X80Y101_BQ;
  assign CLBLL_L_X52Y107_SLICE_X78Y107_B4 = CLBLL_L_X54Y100_SLICE_X82Y100_BQ;
  assign CLBLL_L_X52Y107_SLICE_X78Y107_B5 = CLBLL_R_X57Y101_SLICE_X87Y101_DQ;
  assign CLBLL_L_X52Y107_SLICE_X78Y107_B6 = 1'b1;
  assign CLBLL_L_X52Y107_SLICE_X78Y107_C1 = 1'b1;
  assign CLBLL_L_X52Y107_SLICE_X78Y107_C2 = 1'b1;
  assign CLBLL_L_X52Y107_SLICE_X78Y107_C3 = 1'b1;
  assign CLBLL_L_X52Y107_SLICE_X78Y107_C4 = 1'b1;
  assign CLBLL_L_X52Y107_SLICE_X78Y107_C5 = 1'b1;
  assign CLBLL_L_X52Y107_SLICE_X78Y107_C6 = 1'b1;
  assign CLBLL_L_X52Y107_SLICE_X78Y107_D1 = 1'b1;
  assign CLBLL_L_X52Y107_SLICE_X78Y107_D2 = 1'b1;
  assign CLBLL_L_X52Y107_SLICE_X78Y107_D3 = 1'b1;
  assign CLBLL_L_X52Y107_SLICE_X78Y107_D4 = 1'b1;
  assign CLBLL_L_X52Y107_SLICE_X78Y107_D5 = 1'b1;
  assign CLBLL_L_X52Y107_SLICE_X78Y107_D6 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_A1 = CLBLM_L_X56Y98_SLICE_X85Y98_DQ;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_A2 = CLBLM_L_X64Y96_SLICE_X96Y96_BO6;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_A3 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_A4 = CLBLM_R_X63Y98_SLICE_X95Y98_A5Q;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_A5 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_A6 = CLBLM_L_X50Y105_SLICE_X77Y105_AQ;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_B1 = CLBLM_L_X56Y98_SLICE_X85Y98_DQ;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_B2 = CLBLM_L_X64Y97_SLICE_X96Y97_AQ;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_B3 = CLBLM_L_X64Y96_SLICE_X96Y96_CO5;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_B4 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_B5 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_B6 = CLBLM_R_X49Y105_SLICE_X75Y105_CQ;
  assign CLBLL_L_X52Y107_SLICE_X79Y107_A1 = 1'b1;
  assign CLBLL_L_X52Y107_SLICE_X79Y107_A2 = 1'b1;
  assign CLBLL_L_X52Y107_SLICE_X79Y107_A3 = 1'b1;
  assign CLBLL_L_X52Y107_SLICE_X79Y107_A4 = 1'b1;
  assign CLBLL_L_X52Y107_SLICE_X79Y107_A5 = 1'b1;
  assign CLBLL_L_X52Y107_SLICE_X79Y107_A6 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_C1 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_C2 = CLBLM_L_X64Y96_SLICE_X96Y96_CO6;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLL_L_X52Y107_SLICE_X79Y107_B1 = 1'b1;
  assign CLBLL_L_X52Y107_SLICE_X79Y107_B2 = 1'b1;
  assign CLBLL_L_X52Y107_SLICE_X79Y107_B3 = 1'b1;
  assign CLBLL_L_X52Y107_SLICE_X79Y107_B4 = 1'b1;
  assign CLBLL_L_X52Y107_SLICE_X79Y107_B5 = 1'b1;
  assign CLBLL_L_X52Y107_SLICE_X79Y107_B6 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_D3 = CLBLM_L_X64Y96_SLICE_X96Y96_BO5;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_D4 = CLBLM_L_X50Y104_SLICE_X76Y104_AQ;
  assign CLBLL_L_X52Y107_SLICE_X79Y107_C1 = 1'b1;
  assign CLBLL_L_X52Y107_SLICE_X79Y107_C2 = 1'b1;
  assign CLBLL_L_X52Y107_SLICE_X79Y107_C3 = 1'b1;
  assign CLBLL_L_X52Y107_SLICE_X79Y107_C4 = 1'b1;
  assign CLBLL_L_X52Y107_SLICE_X79Y107_C5 = 1'b1;
  assign CLBLL_L_X52Y107_SLICE_X79Y107_C6 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_D5 = CLBLM_L_X56Y98_SLICE_X85Y98_DQ;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_D6 = CLBLM_R_X63Y98_SLICE_X95Y98_AQ;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_A1 = CLBLM_L_X62Y95_SLICE_X92Y95_AQ;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_A2 = CLBLM_L_X62Y98_SLICE_X92Y98_CQ;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_A3 = CLBLM_L_X62Y98_SLICE_X92Y98_DQ;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_A4 = CLBLM_L_X62Y98_SLICE_X92Y98_AQ;
  assign CLBLL_L_X52Y107_SLICE_X79Y107_D1 = 1'b1;
  assign CLBLL_L_X52Y107_SLICE_X79Y107_D2 = 1'b1;
  assign CLBLL_L_X52Y107_SLICE_X79Y107_D3 = 1'b1;
  assign CLBLL_L_X52Y107_SLICE_X79Y107_D4 = 1'b1;
  assign CLBLL_L_X52Y107_SLICE_X79Y107_D5 = 1'b1;
  assign CLBLL_L_X52Y107_SLICE_X79Y107_D6 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_AX = CLBLM_R_X63Y95_SLICE_X95Y95_D5Q;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_B1 = CLBLM_L_X62Y95_SLICE_X92Y95_AQ;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_B2 = CLBLM_L_X62Y98_SLICE_X92Y98_CQ;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_B3 = CLBLM_L_X62Y98_SLICE_X92Y98_DQ;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_B5 = CLBLM_L_X62Y95_SLICE_X92Y95_A5Q;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_B6 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_BX = CLBLM_L_X64Y96_SLICE_X97Y96_AQ;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_B4 = CLBLM_L_X62Y98_SLICE_X92Y98_AQ;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_C1 = CLBLM_L_X62Y95_SLICE_X92Y95_AQ;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_C2 = CLBLM_L_X62Y98_SLICE_X92Y98_CQ;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_C3 = CLBLM_L_X62Y98_SLICE_X92Y98_DQ;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_C4 = CLBLM_L_X62Y98_SLICE_X92Y98_AQ;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_C5 = CLBLM_L_X62Y95_SLICE_X92Y95_A5Q;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_C6 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_CE = CLBLM_L_X60Y98_SLICE_X91Y98_BQ;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_CI = CLBLM_L_X64Y96_SLICE_X97Y96_BQ;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_CX = CLBLM_L_X64Y96_SLICE_X97Y96_CQ;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_D1 = CLBLM_L_X62Y95_SLICE_X93Y95_DQ;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_D2 = CLBLM_L_X62Y95_SLICE_X93Y95_D5Q;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_D3 = CLBLM_L_X62Y95_SLICE_X93Y95_AQ;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_D4 = CLBLM_L_X62Y95_SLICE_X93Y95_BQ;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_D5 = CLBLM_L_X62Y95_SLICE_X93Y95_CQ;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_D6 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_DI = 1'b1;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_C1 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_DX = 1'b1;
  assign CLBLM_R_X53Y108_SLICE_X81Y108_A1 = CLBLL_R_X57Y100_SLICE_X87Y100_CQ;
  assign CLBLM_R_X53Y108_SLICE_X81Y108_A2 = CLBLL_R_X57Y99_SLICE_X86Y99_AQ;
  assign CLBLM_R_X53Y108_SLICE_X81Y108_A3 = CLBLM_L_X56Y101_SLICE_X85Y101_DQ;
  assign CLBLM_R_X53Y108_SLICE_X81Y108_A4 = CLBLL_R_X57Y101_SLICE_X87Y101_CQ;
  assign CLBLM_R_X53Y108_SLICE_X81Y108_A5 = CLBLL_R_X57Y100_SLICE_X87Y100_BQ;
  assign CLBLM_R_X53Y108_SLICE_X81Y108_A6 = CLBLM_L_X56Y101_SLICE_X85Y101_BQ;
  assign CLBLM_R_X53Y108_SLICE_X81Y108_AX = CLBLM_R_X53Y108_SLICE_X80Y108_CO6;
  assign CLBLM_R_X53Y108_SLICE_X81Y108_B1 = CLBLL_R_X57Y101_SLICE_X87Y101_CQ;
  assign CLBLM_R_X53Y108_SLICE_X81Y108_B2 = CLBLL_R_X57Y99_SLICE_X86Y99_AQ;
  assign CLBLM_R_X53Y108_SLICE_X81Y108_B3 = CLBLM_L_X56Y101_SLICE_X85Y101_DQ;
  assign CLBLM_R_X53Y108_SLICE_X81Y108_B4 = 1'b1;
  assign CLBLM_R_X53Y108_SLICE_X81Y108_B5 = CLBLL_R_X57Y100_SLICE_X87Y100_BQ;
  assign CLBLM_R_X53Y108_SLICE_X81Y108_B6 = 1'b1;
  assign CLBLM_R_X53Y108_SLICE_X81Y108_C1 = 1'b1;
  assign CLBLM_R_X53Y108_SLICE_X81Y108_C2 = 1'b1;
  assign CLBLM_R_X53Y108_SLICE_X81Y108_C3 = 1'b1;
  assign CLBLM_R_X53Y108_SLICE_X81Y108_C4 = 1'b1;
  assign CLBLM_R_X53Y108_SLICE_X81Y108_C5 = 1'b1;
  assign CLBLM_R_X53Y108_SLICE_X81Y108_C6 = 1'b1;
  assign CLBLM_R_X53Y108_SLICE_X81Y108_CIN = CLBLM_R_X53Y107_SLICE_X81Y107_COUT;
  assign CLBLM_R_X53Y108_SLICE_X81Y108_CX = 1'b0;
  assign CLBLM_R_X53Y108_SLICE_X81Y108_D1 = 1'b1;
  assign CLBLM_R_X53Y108_SLICE_X81Y108_D2 = 1'b1;
  assign CLBLM_R_X53Y108_SLICE_X81Y108_D3 = 1'b1;
  assign CLBLM_R_X53Y108_SLICE_X81Y108_D4 = 1'b1;
  assign CLBLM_R_X53Y108_SLICE_X81Y108_D5 = 1'b1;
  assign CLBLM_R_X53Y108_SLICE_X81Y108_D6 = 1'b1;
  assign CLBLM_R_X53Y108_SLICE_X81Y108_DX = 1'b0;
  assign CLBLM_R_X53Y108_SLICE_X80Y108_A1 = CLBLM_L_X56Y101_SLICE_X85Y101_DQ;
  assign CLBLM_R_X53Y108_SLICE_X80Y108_A2 = CLBLL_R_X57Y101_SLICE_X87Y101_CQ;
  assign CLBLM_R_X53Y108_SLICE_X80Y108_A3 = CLBLM_L_X56Y101_SLICE_X85Y101_AQ;
  assign CLBLM_R_X53Y108_SLICE_X80Y108_A4 = CLBLL_R_X57Y101_SLICE_X87Y101_AQ;
  assign CLBLM_R_X53Y108_SLICE_X80Y108_A5 = CLBLL_R_X57Y100_SLICE_X87Y100_AQ;
  assign CLBLM_R_X53Y108_SLICE_X80Y108_A6 = CLBLL_R_X57Y100_SLICE_X87Y100_CQ;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_D1 = 1'b1;
  assign CLBLM_R_X53Y108_SLICE_X80Y108_B1 = CLBLL_R_X57Y100_SLICE_X87Y100_AQ;
  assign CLBLM_R_X53Y108_SLICE_X80Y108_B2 = CLBLL_R_X57Y100_SLICE_X86Y100_BQ;
  assign CLBLM_R_X53Y108_SLICE_X80Y108_B3 = CLBLM_L_X56Y101_SLICE_X85Y101_AQ;
  assign CLBLM_R_X53Y108_SLICE_X80Y108_B4 = CLBLL_R_X57Y100_SLICE_X87Y100_CQ;
  assign CLBLM_R_X53Y108_SLICE_X80Y108_B5 = CLBLM_L_X56Y101_SLICE_X85Y101_DQ;
  assign CLBLM_R_X53Y108_SLICE_X80Y108_B6 = CLBLL_R_X57Y101_SLICE_X87Y101_CQ;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_D4 = 1'b1;
  assign CLBLM_R_X53Y108_SLICE_X80Y108_C1 = CLBLM_L_X56Y101_SLICE_X85Y101_DQ;
  assign CLBLM_R_X53Y108_SLICE_X80Y108_C2 = CLBLL_R_X57Y100_SLICE_X87Y100_BQ;
  assign CLBLM_R_X53Y108_SLICE_X80Y108_C3 = CLBLL_R_X57Y101_SLICE_X87Y101_CQ;
  assign CLBLM_R_X53Y108_SLICE_X80Y108_C4 = CLBLM_L_X56Y101_SLICE_X85Y101_BQ;
  assign CLBLM_R_X53Y108_SLICE_X80Y108_C5 = CLBLL_R_X57Y100_SLICE_X87Y100_CQ;
  assign CLBLM_R_X53Y108_SLICE_X80Y108_C6 = CLBLL_R_X57Y99_SLICE_X86Y99_AQ;
  assign CLBLM_R_X53Y108_SLICE_X80Y108_D1 = 1'b1;
  assign CLBLM_R_X53Y108_SLICE_X80Y108_D2 = 1'b1;
  assign CLBLM_R_X53Y108_SLICE_X80Y108_D3 = 1'b1;
  assign CLBLM_R_X53Y108_SLICE_X80Y108_D4 = 1'b1;
  assign CLBLM_R_X53Y108_SLICE_X80Y108_D5 = 1'b1;
  assign CLBLM_R_X53Y108_SLICE_X80Y108_D6 = 1'b1;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_A1 = CLBLM_L_X50Y106_SLICE_X76Y106_AQ;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_A2 = CLBLM_L_X56Y98_SLICE_X85Y98_DQ;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_A3 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_A4 = CLBLM_R_X63Y98_SLICE_X95Y98_BQ;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_A5 = 1'b1;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_A6 = CLBLM_R_X63Y96_SLICE_X94Y96_AO5;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_B1 = CLBLM_R_X63Y99_SLICE_X95Y99_AQ;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_B2 = CLBLM_L_X50Y107_SLICE_X76Y107_BQ;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_B3 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_B4 = CLBLM_L_X56Y98_SLICE_X85Y98_DQ;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_B5 = CLBLM_R_X63Y96_SLICE_X94Y96_BO5;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_B6 = 1'b1;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_C1 = 1'b1;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_C2 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_C3 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_C4 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_C5 = CLBLM_L_X56Y97_SLICE_X85Y97_AQ;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_C6 = CLBLM_R_X63Y95_SLICE_X95Y95_AQ;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_CE = CLBLM_L_X62Y99_SLICE_X93Y99_AO6;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_D1 = 1'b1;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_D2 = 1'b1;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_D3 = 1'b1;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_D4 = 1'b1;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_D5 = 1'b1;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_D6 = 1'b1;
  assign CLBLM_L_X64Y97_SLICE_X97Y97_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_A1 = CLBLM_R_X63Y97_SLICE_X95Y97_D5Q;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_A2 = CLBLM_R_X63Y97_SLICE_X95Y97_DQ;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_A3 = CLBLM_L_X64Y99_SLICE_X96Y99_AQ;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_A4 = CLBLM_R_X63Y99_SLICE_X94Y99_DO5;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_A5 = CLBLM_R_X65Y102_SLICE_X99Y102_AQ;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_A6 = 1'b1;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_B1 = CLBLM_R_X63Y99_SLICE_X94Y99_DO5;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_B2 = CLBLM_L_X62Y97_SLICE_X92Y97_BQ;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_B3 = CLBLM_L_X62Y97_SLICE_X92Y97_AQ;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_B4 = CLBLM_R_X65Y104_SLICE_X99Y104_BQ;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_B5 = CLBLM_R_X65Y103_SLICE_X99Y103_BQ;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_B6 = 1'b1;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_C1 = CLBLM_L_X64Y96_SLICE_X97Y96_AQ;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_C2 = 1'b1;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_C3 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_C4 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_C5 = CLBLM_L_X56Y97_SLICE_X85Y97_AQ;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_C6 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_CE = CLBLM_L_X60Y98_SLICE_X91Y98_DQ;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_D1 = 1'b1;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_D2 = 1'b1;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_D3 = 1'b1;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_D4 = 1'b1;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_D5 = 1'b1;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_D6 = 1'b1;
  assign CLBLM_L_X64Y97_SLICE_X96Y97_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_D = LIOB33_X0Y103_IOB_X0Y104_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_D = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_A1 = CLBLM_L_X64Y101_SLICE_X96Y101_C_XOR;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_A2 = CLBLM_R_X65Y97_SLICE_X98Y97_AO5;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_A3 = CLBLM_R_X65Y97_SLICE_X98Y97_AO6;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_A4 = CLBLM_L_X64Y98_SLICE_X97Y98_BO6;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_A5 = CLBLM_L_X64Y98_SLICE_X97Y98_DO6;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_A6 = CLBLM_L_X64Y98_SLICE_X97Y98_CO6;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_B1 = CLBLM_L_X64Y96_SLICE_X97Y96_DQ;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_B2 = CLBLM_L_X56Y97_SLICE_X85Y97_AQ;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_B3 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_B4 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_B5 = 1'b1;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_B6 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_C1 = CLBLM_L_X60Y98_SLICE_X90Y98_AQ;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_C2 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_C3 = 1'b1;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_C4 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_C5 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_C6 = CLBLM_R_X65Y101_SLICE_X98Y101_D_XOR;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_CE = CLBLM_L_X60Y98_SLICE_X91Y98_BQ;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_D1 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_D2 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_D3 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_D4 = CLBLM_L_X64Y101_SLICE_X97Y101_D_XOR;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_D5 = CLBLM_L_X62Y101_SLICE_X93Y101_CQ;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_D6 = 1'b1;
  assign CLBLM_L_X64Y98_SLICE_X97Y98_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_A1 = CLBLM_R_X63Y101_SLICE_X95Y101_DO6;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_A2 = CLBLM_R_X65Y97_SLICE_X98Y97_AO6;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_A3 = CLBLM_L_X64Y97_SLICE_X96Y97_CO6;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_A4 = CLBLM_L_X64Y101_SLICE_X96Y101_D_XOR;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_A5 = CLBLM_R_X65Y98_SLICE_X98Y98_DO6;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_A6 = CLBLM_R_X65Y97_SLICE_X98Y97_AO5;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_B1 = CLBLM_R_X63Y95_SLICE_X95Y95_DQ;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_B2 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_B3 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_B4 = CLBLM_L_X56Y97_SLICE_X85Y97_AQ;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_B5 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_B6 = CLBLM_L_X64Y98_SLICE_X96Y98_CO6;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_C1 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_C2 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_C3 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_C4 = CLBLM_L_X64Y100_SLICE_X97Y100_A_XOR;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_C5 = CLBLM_L_X64Y98_SLICE_X96Y98_DO6;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_C6 = CLBLM_L_X62Y100_SLICE_X92Y100_AQ;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_CE = CLBLM_L_X60Y98_SLICE_X91Y98_BQ;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_D1 = CLBLM_L_X60Y98_SLICE_X90Y98_AQ;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_D2 = CLBLM_L_X62Y100_SLICE_X92Y100_AQ;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_D3 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_D4 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_D5 = CLBLM_R_X65Y100_SLICE_X99Y100_CQ;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_D6 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_L_X64Y98_SLICE_X96Y98_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_C3 = CLBLM_L_X64Y97_SLICE_X96Y97_A5Q;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_C4 = CLBLM_R_X49Y106_SLICE_X74Y106_AQ;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_C5 = CLBLM_L_X56Y98_SLICE_X85Y98_DQ;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_C6 = 1'b1;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_CE = CLBLM_L_X62Y99_SLICE_X93Y99_AO6;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_D1 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X64Y96_SLICE_X97Y96_D2 = 1'b1;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_A1 = CLBLM_R_X65Y97_SLICE_X98Y97_AO5;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_A2 = CLBLM_L_X64Y100_SLICE_X96Y100_C_XOR;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_A3 = CLBLM_R_X65Y97_SLICE_X98Y97_AO6;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_A4 = CLBLM_R_X63Y100_SLICE_X95Y100_BO6;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_A5 = CLBLM_L_X64Y97_SLICE_X97Y97_CO6;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_A6 = CLBLM_R_X65Y99_SLICE_X99Y99_DO6;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_B1 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_B2 = CLBLM_L_X60Y98_SLICE_X90Y98_AQ;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_B3 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_B4 = 1'b1;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_B5 = CLBLM_R_X65Y102_SLICE_X98Y102_C_XOR;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_B6 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_C1 = CLBLM_L_X64Y101_SLICE_X97Y101_C_XOR;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_C2 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_C3 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_C4 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_C5 = 1'b1;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_C6 = CLBLM_L_X62Y101_SLICE_X93Y101_BQ;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_CE = CLBLM_L_X60Y98_SLICE_X91Y98_BQ;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_D1 = 1'b1;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_D2 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_D3 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_D4 = CLBLM_L_X56Y97_SLICE_X85Y97_AQ;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_D5 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_D6 = CLBLM_L_X64Y96_SLICE_X97Y96_BQ;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_A5 = CLBLM_L_X62Y95_SLICE_X92Y95_A5Q;
  assign CLBLM_L_X64Y99_SLICE_X97Y99_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_A6 = 1'b1;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_A1 = CLBLM_R_X63Y101_SLICE_X95Y101_CO6;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_A2 = CLBLM_L_X64Y99_SLICE_X97Y99_BO6;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_A3 = CLBLM_R_X65Y97_SLICE_X98Y97_AO5;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_A4 = CLBLM_R_X65Y97_SLICE_X98Y97_AO6;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_AI = CLBLM_R_X63Y95_SLICE_X95Y95_C5Q;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_A5 = CLBLM_L_X64Y102_SLICE_X96Y102_B_XOR;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_A6 = CLBLM_L_X64Y99_SLICE_X96Y99_CO6;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_B1 = CLBLM_L_X64Y99_SLICE_X96Y99_DO6;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_B2 = CLBLM_L_X64Y101_SLICE_X96Y101_B_XOR;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_B3 = CLBLM_R_X65Y97_SLICE_X98Y97_AO5;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_B4 = CLBLM_L_X64Y99_SLICE_X97Y99_CO6;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_B5 = CLBLM_R_X65Y96_SLICE_X98Y96_BO6;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_B6 = CLBLM_R_X65Y97_SLICE_X98Y97_AO6;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_C1 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_C2 = CLBLM_L_X56Y97_SLICE_X85Y97_AQ;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_C3 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_C4 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_C5 = 1'b1;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_C6 = CLBLM_L_X64Y96_SLICE_X97Y96_CQ;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_CE = CLBLM_L_X60Y98_SLICE_X91Y98_BQ;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_D1 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_D2 = 1'b1;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_D3 = CLBLM_L_X60Y98_SLICE_X90Y98_AQ;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_D4 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_D5 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_D6 = CLBLM_R_X65Y101_SLICE_X98Y101_C_XOR;
  assign CLBLM_L_X64Y99_SLICE_X96Y99_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X64Y96_SLICE_X96Y96_BI = CLBLM_L_X64Y96_SLICE_X97Y96_DQ;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_A1 = CLBLM_R_X65Y100_SLICE_X99Y100_CQ;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_A2 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_A3 = CLBLM_L_X62Y100_SLICE_X92Y100_AQ;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_A4 = CLBLM_R_X49Y104_SLICE_X75Y104_DQ;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_A5 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_A6 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_AX = CLBLM_R_X65Y100_SLICE_X99Y100_CQ;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_B1 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_B2 = CLBLM_R_X65Y100_SLICE_X99Y100_AQ;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_B3 = CLBLM_R_X49Y106_SLICE_X75Y106_CQ;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_B4 = CLBLM_L_X62Y100_SLICE_X92Y100_BQ;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_B5 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_B6 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_BX = CLBLM_R_X65Y100_SLICE_X99Y100_AQ;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_C1 = CLBLM_L_X62Y101_SLICE_X93Y101_AQ;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_C2 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_C3 = CLBLM_R_X65Y106_SLICE_X98Y106_CQ;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_C4 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_C5 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_C6 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_CE = CLBLM_L_X62Y101_SLICE_X93Y101_AO6;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_CX = CLBLM_R_X65Y106_SLICE_X98Y106_CQ;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_D1 = CLBLM_L_X64Y106_SLICE_X97Y106_DQ;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_D2 = CLBLM_L_X62Y100_SLICE_X92Y100_CQ;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_D3 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_D4 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_D5 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_D6 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_DX = CLBLM_L_X64Y106_SLICE_X97Y106_DQ;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_A1 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_A2 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_A3 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_A4 = CLBLM_R_X65Y100_SLICE_X99Y100_AQ;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_A5 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_A6 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_AX = CLBLM_R_X65Y100_SLICE_X99Y100_CQ;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_B1 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_B2 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_B3 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_B4 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_B5 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_B6 = CLBLM_R_X65Y106_SLICE_X98Y106_CQ;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_D = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_D = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_BX = 1'b0;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_C1 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_C2 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_C3 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_C4 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_C5 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_C6 = CLBLM_L_X64Y106_SLICE_X97Y106_DQ;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_CX = 1'b0;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_D1 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_D2 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_D3 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_D4 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_D5 = 1'b1;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_D6 = CLBLM_R_X65Y100_SLICE_X99Y100_BQ;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_DX = 1'b0;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_A1 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_A2 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_A3 = CLBLM_L_X64Y100_SLICE_X97Y100_AQ;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_A4 = CLBLM_R_X65Y100_SLICE_X99Y100_BQ;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_A5 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_A6 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_AX = CLBLM_R_X65Y100_SLICE_X99Y100_BQ;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_B1 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_B2 = CLBLM_R_X65Y106_SLICE_X98Y106_DQ;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_B3 = CLBLM_L_X64Y100_SLICE_X97Y100_BQ;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_B4 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_B5 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_B6 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_BX = CLBLM_R_X65Y106_SLICE_X98Y106_DQ;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_C1 = CLBLM_R_X63Y103_SLICE_X95Y103_BQ;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_C2 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_C3 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_C4 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_C5 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_C6 = CLBLM_L_X62Y101_SLICE_X93Y101_BQ;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_CIN = CLBLM_L_X64Y100_SLICE_X97Y100_COUT;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_CX = CLBLM_R_X63Y103_SLICE_X95Y103_BQ;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_D1 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_D2 = CLBLM_L_X62Y101_SLICE_X93Y101_CQ;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_D3 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_D4 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_D5 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_D6 = CLBLM_R_X63Y101_SLICE_X95Y101_AQ;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_DX = CLBLM_R_X63Y101_SLICE_X95Y101_AQ;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_A1 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_A2 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_A3 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_A4 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_A5 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_A6 = CLBLM_R_X65Y106_SLICE_X98Y106_DQ;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_B3 = CLBLM_L_X64Y96_SLICE_X97Y96_AQ;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_AX = 1'b0;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_B1 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_B2 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_B3 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_B4 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_B5 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_B6 = CLBLM_R_X63Y103_SLICE_X95Y103_BQ;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_B4 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_BX = 1'b0;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_C1 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_C2 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_C3 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_C4 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_C5 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_C6 = CLBLM_R_X63Y101_SLICE_X95Y101_AQ;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_B6 = CLBLM_L_X62Y98_SLICE_X92Y98_CQ;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_CIN = CLBLM_L_X64Y100_SLICE_X96Y100_COUT;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_CX = 1'b0;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_D1 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_D2 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_D3 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_D4 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_D5 = 1'b1;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_D6 = CLBLM_R_X63Y103_SLICE_X95Y103_CQ;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_DX = 1'b0;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_C4 = CLBLM_L_X50Y105_SLICE_X77Y105_AQ;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_C6 = 1'b1;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_CE = CLBLM_R_X63Y100_SLICE_X94Y100_BO6;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_D1 = CLBLM_L_X64Y97_SLICE_X96Y97_AQ;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_D4 = CLBLM_R_X49Y105_SLICE_X75Y105_CQ;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_D = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_A1 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_A2 = CLBLM_L_X64Y102_SLICE_X97Y102_BQ;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_A3 = CLBLM_R_X63Y103_SLICE_X95Y103_CQ;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_A4 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_A5 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_A6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1 = CLBLM_R_X49Y111_SLICE_X74Y111_CQ;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_AX = CLBLM_R_X63Y103_SLICE_X95Y103_CQ;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_B1 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_B2 = CLBLM_R_X65Y107_SLICE_X98Y107_DQ;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_B3 = CLBLM_L_X64Y102_SLICE_X97Y102_CQ;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_B4 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_D3 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_B5 = CLBLM_R_X49Y108_SLICE_X75Y108_DQ;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_D4 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_B6 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_BX = CLBLM_R_X65Y107_SLICE_X98Y107_DQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_C1 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_C2 = CLBLM_R_X65Y107_SLICE_X98Y107_AQ;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_C3 = CLBLM_R_X49Y107_SLICE_X75Y107_DQ;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_C4 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_C5 = CLBLM_L_X64Y102_SLICE_X97Y102_AQ;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_C6 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_CE = CLBLM_L_X62Y101_SLICE_X93Y101_AO6;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_CIN = CLBLM_L_X64Y101_SLICE_X97Y101_COUT;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_D1 = CLBLM_R_X49Y107_SLICE_X74Y107_AQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1 = CLBLM_R_X49Y109_SLICE_X74Y109_BQ;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_CX = CLBLM_L_X64Y102_SLICE_X97Y102_AQ;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_D1 = CLBLM_R_X65Y107_SLICE_X98Y107_BQ;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_D2 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_D3 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_D4 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_D5 = CLBLM_L_X64Y102_SLICE_X97Y102_AQ;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_D6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_A1 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_A2 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_A3 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_A4 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_A5 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_A6 = CLBLM_R_X65Y107_SLICE_X98Y107_DQ;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_AX = 1'b0;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_B1 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_B2 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_B3 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_B4 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_B5 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_B6 = CLBLM_R_X65Y107_SLICE_X98Y107_AQ;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_BX = 1'b0;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_C1 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_C2 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_C3 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_C4 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_C5 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_C6 = CLBLM_R_X65Y107_SLICE_X98Y107_BQ;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_CIN = CLBLM_L_X64Y101_SLICE_X96Y101_COUT;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_T1 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_CX = 1'b0;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_D1 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_D2 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_D3 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_D4 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_D5 = 1'b1;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_D6 = CLBLM_R_X65Y107_SLICE_X98Y107_CQ;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_DX = 1'b0;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_D = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_D = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_A1 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_A2 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_A3 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_A4 = CLBLM_R_X65Y107_SLICE_X98Y107_BQ;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_A5 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_A6 = CLBLM_R_X65Y107_SLICE_X98Y107_CQ;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_AX = CLBLM_R_X65Y107_SLICE_X98Y107_BQ;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_B1 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_B2 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_B3 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_B4 = CLBLM_R_X65Y106_SLICE_X98Y106_AQ;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_B5 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_B6 = CLBLM_R_X65Y107_SLICE_X98Y107_CQ;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_BX = CLBLM_R_X65Y107_SLICE_X98Y107_CQ;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_C1 = CLBLM_L_X64Y106_SLICE_X97Y106_AQ;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_C2 = CLBLM_R_X65Y106_SLICE_X98Y106_AQ;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_C3 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_C4 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_C5 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_C6 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_CIN = CLBLM_L_X64Y102_SLICE_X97Y102_COUT;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_CX = CLBLM_R_X65Y106_SLICE_X98Y106_AQ;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_D1 = CLBLM_L_X64Y106_SLICE_X97Y106_AQ;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_D2 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_D3 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_D4 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_D5 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_D6 = CLBLM_R_X63Y103_SLICE_X95Y103_AQ;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_DX = CLBLM_L_X64Y106_SLICE_X97Y106_AQ;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_A1 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_A2 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_A3 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_A4 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_A5 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_A6 = CLBLM_R_X65Y106_SLICE_X98Y106_AQ;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_AX = 1'b0;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_B1 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_B2 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_B3 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_B4 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_B5 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_B6 = CLBLM_L_X64Y106_SLICE_X97Y106_AQ;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_BX = 1'b0;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_C1 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_C2 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_C3 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_C4 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_C5 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_C6 = CLBLM_R_X63Y103_SLICE_X95Y103_AQ;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_CIN = CLBLM_L_X64Y102_SLICE_X96Y102_COUT;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_CX = 1'b0;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_D1 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_D2 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_D3 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_D4 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_D5 = 1'b1;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_D6 = CLBLM_R_X65Y106_SLICE_X98Y106_BQ;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_DX = 1'b0;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_A1 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_A2 = CLBLM_R_X65Y106_SLICE_X98Y106_BQ;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_A3 = CLBLM_R_X63Y103_SLICE_X95Y103_AQ;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_A4 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_A5 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_A6 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_AX = CLBLM_R_X63Y103_SLICE_X95Y103_AQ;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_B1 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_B2 = CLBLM_L_X64Y106_SLICE_X97Y106_BQ;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_B3 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_B4 = CLBLM_R_X65Y106_SLICE_X98Y106_BQ;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_B5 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_B6 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_BX = CLBLM_R_X65Y106_SLICE_X98Y106_BQ;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_C1 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_C2 = CLBLM_L_X64Y106_SLICE_X97Y106_BQ;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_C3 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_C4 = CLBLM_L_X64Y106_SLICE_X97Y106_CQ;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_C5 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_C6 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_CIN = CLBLM_L_X64Y103_SLICE_X97Y103_COUT;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_CX = 1'b0;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_D1 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_D2 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_D3 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_D4 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_D5 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_D6 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X97Y104_DX = 1'b0;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_A1 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_A2 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_A3 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_A4 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_A5 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_A6 = CLBLM_L_X64Y106_SLICE_X97Y106_BQ;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_AX = 1'b0;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_B1 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_B2 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_B3 = 1'b1;
  assign CLBLL_R_X57Y99_SLICE_X86Y99_A4 = CLBLL_L_X54Y99_SLICE_X82Y99_AQ;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_B4 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_B5 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_B6 = CLBLM_L_X64Y106_SLICE_X97Y106_CQ;
  assign CLBLL_R_X57Y99_SLICE_X86Y99_A5 = CLBLL_L_X54Y98_SLICE_X83Y98_BQ;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_BX = 1'b0;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_C1 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_C2 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_C3 = 1'b1;
  assign CLBLL_R_X57Y99_SLICE_X86Y99_A6 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_C4 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_C5 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_C6 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_CIN = CLBLM_L_X64Y103_SLICE_X96Y103_COUT;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_CX = 1'b0;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_D1 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_D2 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_D3 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_D4 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_D5 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_D6 = 1'b1;
  assign CLBLM_L_X64Y104_SLICE_X96Y104_DX = 1'b0;
  assign CLBLL_R_X57Y99_SLICE_X86Y99_B3 = CLBLM_L_X56Y99_SLICE_X85Y99_BQ;
  assign CLBLL_R_X57Y99_SLICE_X86Y99_C2 = 1'b1;
  assign CLBLL_R_X57Y99_SLICE_X86Y99_C3 = 1'b1;
  assign CLBLL_R_X57Y99_SLICE_X86Y99_C4 = 1'b1;
  assign CLBLL_R_X57Y99_SLICE_X86Y99_C5 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_D = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_D = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_A1 = CLBLM_R_X63Y105_SLICE_X95Y105_C_XOR;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_A2 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_A3 = CLBLM_L_X64Y105_SLICE_X97Y105_AQ;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_A4 = CLBLM_L_X64Y105_SLICE_X97Y105_BO6;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_A5 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_A6 = CLBLM_L_X62Y105_SLICE_X92Y105_BO5;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_B1 = CLBLM_R_X63Y105_SLICE_X95Y105_C_XOR;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_B2 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_B3 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_B4 = CLBLM_R_X49Y106_SLICE_X74Y106_AQ;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_B5 = CLBLM_L_X62Y105_SLICE_X93Y105_AO6;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_B6 = CLBLM_R_X63Y105_SLICE_X94Y105_D_XOR;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_C1 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_C2 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_C3 = CLBLM_R_X49Y104_SLICE_X75Y104_DQ;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_C4 = CLBLM_L_X64Y103_SLICE_X97Y103_A_XOR;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_C5 = 1'b1;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_C6 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_CE = CLBLM_L_X62Y100_SLICE_X92Y100_CO6;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_D1 = CLBLM_L_X64Y104_SLICE_X97Y104_C_XOR;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_D2 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_D3 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_D4 = 1'b1;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_D5 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_D6 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLM_L_X64Y105_SLICE_X97Y105_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_A1 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_A2 = CLBLM_L_X62Y105_SLICE_X92Y105_BO5;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_A3 = CLBLM_L_X64Y105_SLICE_X96Y105_AQ;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_A4 = CLBLM_L_X64Y105_SLICE_X96Y105_BO6;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_A5 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_A6 = CLBLM_R_X63Y105_SLICE_X95Y105_B_XOR;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_B1 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_B2 = CLBLM_R_X49Y105_SLICE_X75Y105_CQ;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_B3 = CLBLM_L_X62Y105_SLICE_X93Y105_AO6;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_B4 = CLBLM_R_X63Y105_SLICE_X95Y105_B_XOR;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_B5 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_B6 = CLBLM_R_X63Y105_SLICE_X94Y105_C_XOR;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_C1 = CLBLM_L_X64Y103_SLICE_X97Y103_C_XOR;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_C2 = 1'b1;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_C3 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_C4 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_C5 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_C6 = CLBLM_R_X49Y106_SLICE_X75Y106_DQ;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_CE = CLBLM_L_X62Y100_SLICE_X92Y100_CO6;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_D1 = CLBLM_R_X49Y111_SLICE_X74Y111_AQ;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_D2 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_D3 = CLBLM_L_X64Y105_SLICE_X96Y105_AQ;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_D4 = 1'b1;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_D5 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_D6 = CLBLM_L_X64Y107_SLICE_X96Y107_BQ;
  assign CLBLM_L_X64Y105_SLICE_X96Y105_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_A1 = CLBLL_R_X57Y103_SLICE_X86Y103_AQ;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_A2 = 1'b1;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_A3 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_A4 = CLBLM_L_X64Y108_SLICE_X96Y108_BQ;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_A5 = CLBLM_R_X65Y103_SLICE_X99Y103_AQ;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_A6 = CLBLL_R_X57Y103_SLICE_X86Y103_A5Q;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_B1 = CLBLL_R_X57Y103_SLICE_X86Y103_AQ;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_B2 = 1'b1;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_B3 = CLBLM_R_X63Y105_SLICE_X94Y105_AQ;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_B4 = CLBLM_R_X65Y105_SLICE_X98Y105_BQ;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_B5 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_B6 = CLBLL_R_X57Y103_SLICE_X86Y103_A5Q;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_A3 = CLBLM_L_X64Y98_SLICE_X97Y98_AQ;
  assign CLBLM_R_X47Y119_SLICE_X73Y119_C6 = 1'b1;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_C1 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_C2 = CLBLL_R_X57Y103_SLICE_X86Y103_A5Q;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_C3 = CLBLM_L_X64Y109_SLICE_X96Y109_A5Q;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_C4 = CLBLL_R_X57Y103_SLICE_X86Y103_AQ;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_C5 = CLBLM_R_X65Y105_SLICE_X99Y105_AQ;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_C6 = 1'b1;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_CE = CLBLM_L_X62Y105_SLICE_X93Y105_DO6;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_D1 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_D2 = CLBLL_R_X57Y103_SLICE_X86Y103_A5Q;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_D3 = CLBLM_L_X64Y99_SLICE_X97Y99_AQ;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_D4 = CLBLL_R_X57Y103_SLICE_X86Y103_AQ;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_D5 = 1'b1;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_D6 = CLBLM_R_X63Y104_SLICE_X94Y104_BQ;
  assign CLBLM_L_X64Y106_SLICE_X97Y106_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_A1 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_A2 = CLBLM_L_X62Y105_SLICE_X92Y105_BO5;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_A3 = CLBLM_L_X64Y106_SLICE_X96Y106_AQ;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_A4 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_A5 = CLBLM_L_X64Y106_SLICE_X96Y106_CO6;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_A6 = CLBLM_R_X63Y106_SLICE_X95Y106_B_XOR;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_B1 = CLBLM_R_X63Y106_SLICE_X95Y106_C_XOR;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_B2 = CLBLM_L_X64Y106_SLICE_X96Y106_BQ;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_B3 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_B4 = CLBLM_L_X64Y106_SLICE_X96Y106_DO6;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_B5 = CLBLM_L_X62Y105_SLICE_X92Y105_BO5;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_B6 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_B2 = CLBLM_R_X63Y98_SLICE_X94Y98_CQ;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_B3 = CLBLM_R_X63Y98_SLICE_X94Y98_C5Q;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_C1 = CLBLM_L_X50Y107_SLICE_X76Y107_BQ;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_C2 = CLBLM_L_X62Y105_SLICE_X93Y105_AO6;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_C3 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_C4 = CLBLM_R_X63Y106_SLICE_X95Y106_B_XOR;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_C5 = CLBLM_R_X63Y106_SLICE_X94Y106_C_XOR;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_C6 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_CE = CLBLM_L_X62Y100_SLICE_X92Y100_CO6;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_B4 = CLBLM_R_X65Y98_SLICE_X98Y98_AQ;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_B5 = CLBLM_R_X65Y104_SLICE_X99Y104_AQ;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_B6 = 1'b1;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_D1 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_D2 = CLBLM_L_X62Y105_SLICE_X93Y105_AO6;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_D3 = CLBLM_L_X50Y107_SLICE_X77Y107_AQ;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_D4 = CLBLM_R_X63Y106_SLICE_X94Y106_D_XOR;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_D5 = CLBLM_R_X63Y106_SLICE_X95Y106_C_XOR;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_D6 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X64Y106_SLICE_X96Y106_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_D3 = CLBLM_R_X65Y101_SLICE_X99Y101_AQ;
  assign CLBLM_L_X64Y107_SLICE_X97Y107_A1 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X64Y107_SLICE_X97Y107_A2 = CLBLM_R_X63Y107_SLICE_X95Y107_C_XOR;
  assign CLBLM_L_X64Y107_SLICE_X97Y107_A3 = CLBLM_L_X64Y107_SLICE_X97Y107_AQ;
  assign CLBLM_L_X64Y107_SLICE_X97Y107_A4 = CLBLM_L_X64Y107_SLICE_X97Y107_DO6;
  assign CLBLM_L_X64Y107_SLICE_X97Y107_A5 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X64Y107_SLICE_X97Y107_A6 = CLBLM_L_X62Y105_SLICE_X92Y105_BO5;
  assign CLBLM_L_X64Y107_SLICE_X97Y107_B1 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X64Y107_SLICE_X97Y107_B2 = CLBLM_L_X64Y107_SLICE_X97Y107_BQ;
  assign CLBLM_L_X64Y107_SLICE_X97Y107_B3 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X64Y107_SLICE_X97Y107_B4 = CLBLM_R_X63Y106_SLICE_X95Y106_D_XOR;
  assign CLBLM_L_X64Y107_SLICE_X97Y107_B5 = CLBLM_L_X62Y105_SLICE_X92Y105_BO5;
  assign CLBLM_L_X64Y107_SLICE_X97Y107_B6 = CLBLM_L_X64Y107_SLICE_X97Y107_CO6;
  assign CLBLM_L_X64Y107_SLICE_X97Y107_C1 = CLBLM_R_X63Y107_SLICE_X94Y107_A_XOR;
  assign CLBLM_L_X64Y107_SLICE_X97Y107_C2 = CLBLM_L_X50Y104_SLICE_X76Y104_AQ;
  assign CLBLM_L_X64Y107_SLICE_X97Y107_C3 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X64Y107_SLICE_X97Y107_C4 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X64Y107_SLICE_X97Y107_C5 = CLBLM_L_X62Y105_SLICE_X93Y105_AO6;
  assign CLBLM_L_X64Y107_SLICE_X97Y107_C6 = CLBLM_R_X63Y106_SLICE_X95Y106_D_XOR;
  assign CLBLM_L_X64Y107_SLICE_X97Y107_CE = CLBLM_R_X63Y100_SLICE_X94Y100_CO6;
  assign CLBLM_L_X64Y107_SLICE_X97Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X64Y107_SLICE_X97Y107_D1 = CLBLM_R_X49Y106_SLICE_X74Y106_AQ;
  assign CLBLM_L_X64Y107_SLICE_X97Y107_D2 = CLBLM_R_X63Y107_SLICE_X94Y107_D_XOR;
  assign CLBLM_L_X64Y107_SLICE_X97Y107_D3 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X64Y107_SLICE_X97Y107_D4 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X64Y107_SLICE_X97Y107_D5 = CLBLM_L_X62Y105_SLICE_X93Y105_AO6;
  assign CLBLM_L_X64Y107_SLICE_X97Y107_D6 = CLBLM_R_X63Y107_SLICE_X95Y107_C_XOR;
  assign CLBLM_L_X64Y107_SLICE_X97Y107_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X64Y107_SLICE_X96Y107_A1 = CLBLM_R_X63Y107_SLICE_X95Y107_A_XOR;
  assign CLBLM_L_X64Y107_SLICE_X96Y107_A2 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X64Y107_SLICE_X96Y107_A3 = CLBLM_L_X64Y107_SLICE_X96Y107_AQ;
  assign CLBLM_L_X64Y107_SLICE_X96Y107_A4 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X64Y107_SLICE_X96Y107_A5 = CLBLM_L_X62Y105_SLICE_X92Y105_BO5;
  assign CLBLM_L_X64Y107_SLICE_X96Y107_A6 = CLBLM_L_X64Y107_SLICE_X96Y107_CO6;
  assign CLBLM_L_X64Y107_SLICE_X96Y107_B1 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X64Y107_SLICE_X96Y107_B2 = CLBLM_L_X64Y107_SLICE_X96Y107_BQ;
  assign CLBLM_L_X64Y107_SLICE_X96Y107_B3 = CLBLM_L_X64Y107_SLICE_X96Y107_DO6;
  assign CLBLM_L_X64Y107_SLICE_X96Y107_B4 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X64Y107_SLICE_X96Y107_B5 = CLBLM_L_X62Y105_SLICE_X92Y105_BO5;
  assign CLBLM_L_X64Y107_SLICE_X96Y107_B6 = CLBLM_R_X63Y107_SLICE_X95Y107_B_XOR;
  assign CLBLM_L_X64Y107_SLICE_X96Y107_C1 = CLBLM_R_X63Y107_SLICE_X94Y107_B_XOR;
  assign CLBLM_L_X64Y107_SLICE_X96Y107_C2 = CLBLM_L_X50Y105_SLICE_X77Y105_AQ;
  assign CLBLM_L_X64Y107_SLICE_X96Y107_C3 = CLBLM_L_X62Y105_SLICE_X93Y105_AO6;
  assign CLBLM_L_X64Y107_SLICE_X96Y107_C4 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X64Y107_SLICE_X96Y107_C5 = CLBLM_R_X63Y107_SLICE_X95Y107_A_XOR;
  assign CLBLM_L_X64Y107_SLICE_X96Y107_C6 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X64Y107_SLICE_X96Y107_CE = CLBLM_R_X63Y100_SLICE_X94Y100_CO6;
  assign CLBLM_L_X64Y107_SLICE_X96Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X64Y107_SLICE_X96Y107_D1 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X64Y107_SLICE_X96Y107_D2 = CLBLM_R_X63Y107_SLICE_X94Y107_C_XOR;
  assign CLBLM_L_X64Y107_SLICE_X96Y107_D3 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X64Y107_SLICE_X96Y107_D4 = CLBLM_R_X63Y107_SLICE_X95Y107_B_XOR;
  assign CLBLM_L_X64Y107_SLICE_X96Y107_D5 = CLBLM_L_X62Y105_SLICE_X93Y105_AO6;
  assign CLBLM_L_X64Y107_SLICE_X96Y107_D6 = CLBLM_R_X49Y105_SLICE_X75Y105_CQ;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_D = LIOB33_X0Y115_IOB_X0Y116_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_D = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_L_X64Y107_SLICE_X96Y107_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X64Y108_SLICE_X97Y108_A1 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X64Y108_SLICE_X97Y108_A2 = CLBLM_R_X63Y108_SLICE_X95Y108_A_XOR;
  assign CLBLM_L_X64Y108_SLICE_X97Y108_A3 = CLBLM_L_X64Y108_SLICE_X97Y108_AQ;
  assign CLBLM_L_X64Y108_SLICE_X97Y108_A4 = CLBLM_L_X64Y108_SLICE_X97Y108_BO6;
  assign CLBLM_L_X64Y108_SLICE_X97Y108_A5 = CLBLM_L_X62Y105_SLICE_X92Y105_BO5;
  assign CLBLM_L_X64Y108_SLICE_X97Y108_A6 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X64Y108_SLICE_X97Y108_B1 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X64Y108_SLICE_X97Y108_B2 = CLBLM_L_X62Y105_SLICE_X93Y105_AO6;
  assign CLBLM_L_X64Y108_SLICE_X97Y108_B3 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X64Y108_SLICE_X97Y108_B4 = CLBLM_L_X50Y106_SLICE_X76Y106_CQ;
  assign CLBLM_L_X64Y108_SLICE_X97Y108_B5 = CLBLM_R_X63Y108_SLICE_X95Y108_A_XOR;
  assign CLBLM_L_X64Y108_SLICE_X97Y108_B6 = CLBLM_R_X63Y108_SLICE_X94Y108_B_XOR;
  assign CLBLM_L_X64Y108_SLICE_X97Y108_C1 = 1'b1;
  assign CLBLM_L_X64Y108_SLICE_X97Y108_C2 = 1'b1;
  assign CLBLM_L_X64Y108_SLICE_X97Y108_C3 = 1'b1;
  assign CLBLM_L_X64Y108_SLICE_X97Y108_C4 = 1'b1;
  assign CLBLM_L_X60Y96_SLICE_X91Y96_A1 = 1'b1;
  assign CLBLM_L_X60Y96_SLICE_X91Y96_A2 = 1'b1;
  assign CLBLM_L_X60Y96_SLICE_X91Y96_A3 = 1'b1;
  assign CLBLM_L_X60Y96_SLICE_X91Y96_A4 = 1'b1;
  assign CLBLM_L_X60Y96_SLICE_X91Y96_A5 = 1'b1;
  assign CLBLM_L_X60Y96_SLICE_X91Y96_A6 = 1'b1;
  assign CLBLM_L_X64Y108_SLICE_X97Y108_C5 = 1'b1;
  assign CLBLM_L_X64Y108_SLICE_X97Y108_C6 = 1'b1;
  assign CLBLM_L_X64Y108_SLICE_X97Y108_CE = CLBLM_R_X63Y100_SLICE_X94Y100_CO6;
  assign CLBLM_L_X60Y96_SLICE_X91Y96_B1 = 1'b1;
  assign CLBLM_L_X60Y96_SLICE_X91Y96_B2 = 1'b1;
  assign CLBLM_L_X60Y96_SLICE_X91Y96_B3 = 1'b1;
  assign CLBLM_L_X60Y96_SLICE_X91Y96_B4 = 1'b1;
  assign CLBLM_L_X60Y96_SLICE_X91Y96_B5 = 1'b1;
  assign CLBLM_L_X60Y96_SLICE_X91Y96_B6 = 1'b1;
  assign CLBLM_L_X64Y108_SLICE_X97Y108_D1 = 1'b1;
  assign CLBLM_L_X64Y108_SLICE_X97Y108_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X60Y96_SLICE_X91Y96_C1 = 1'b1;
  assign CLBLM_L_X60Y96_SLICE_X91Y96_C2 = 1'b1;
  assign CLBLM_L_X60Y96_SLICE_X91Y96_C3 = 1'b1;
  assign CLBLM_L_X64Y108_SLICE_X96Y108_A1 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X64Y108_SLICE_X96Y108_A2 = CLBLM_L_X62Y105_SLICE_X92Y105_BO5;
  assign CLBLM_L_X64Y108_SLICE_X96Y108_A3 = CLBLM_L_X64Y108_SLICE_X96Y108_AQ;
  assign CLBLM_L_X64Y108_SLICE_X96Y108_A4 = CLBLM_R_X63Y107_SLICE_X95Y107_D_XOR;
  assign CLBLM_L_X64Y108_SLICE_X96Y108_A5 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X64Y108_SLICE_X96Y108_A6 = CLBLM_L_X64Y108_SLICE_X96Y108_CO6;
  assign CLBLM_L_X60Y96_SLICE_X91Y96_C6 = 1'b1;
  assign CLBLM_L_X60Y96_SLICE_X91Y96_C4 = 1'b1;
  assign CLBLM_L_X60Y96_SLICE_X91Y96_C5 = 1'b1;
  assign CLBLM_L_X64Y108_SLICE_X96Y108_B1 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X60Y96_SLICE_X91Y96_D2 = 1'b1;
  assign CLBLM_L_X64Y108_SLICE_X96Y108_B2 = CLBLM_L_X64Y108_SLICE_X96Y108_DO6;
  assign CLBLM_L_X64Y108_SLICE_X96Y108_B3 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X64Y108_SLICE_X96Y108_B4 = CLBLM_L_X62Y105_SLICE_X93Y105_AO6;
  assign CLBLM_L_X64Y108_SLICE_X96Y108_B5 = CLBLM_R_X63Y108_SLICE_X94Y108_D_XOR;
  assign CLBLM_L_X64Y108_SLICE_X96Y108_B6 = CLBLM_R_X63Y108_SLICE_X95Y108_C_XOR;
  assign CLBLM_L_X60Y96_SLICE_X91Y96_D1 = 1'b1;
  assign CLBLM_L_X60Y96_SLICE_X91Y96_D3 = 1'b1;
  assign CLBLM_L_X60Y96_SLICE_X91Y96_D4 = 1'b1;
  assign CLBLM_L_X64Y108_SLICE_X96Y108_C1 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X64Y108_SLICE_X96Y108_C2 = CLBLM_L_X50Y106_SLICE_X76Y106_AQ;
  assign CLBLM_L_X64Y108_SLICE_X96Y108_C3 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X64Y108_SLICE_X96Y108_C4 = CLBLM_R_X63Y107_SLICE_X95Y107_D_XOR;
  assign CLBLM_L_X64Y108_SLICE_X96Y108_C5 = CLBLM_R_X63Y108_SLICE_X94Y108_A_XOR;
  assign CLBLM_L_X60Y96_SLICE_X90Y96_A4 = 1'b1;
  assign CLBLM_L_X60Y96_SLICE_X90Y96_A5 = 1'b1;
  assign CLBLM_L_X60Y96_SLICE_X90Y96_A6 = 1'b1;
  assign CLBLM_L_X64Y108_SLICE_X96Y108_C6 = CLBLM_L_X62Y105_SLICE_X93Y105_AO6;
  assign CLBLM_L_X64Y108_SLICE_X96Y108_CE = CLBLM_R_X63Y100_SLICE_X94Y100_CO6;
  assign CLBLM_L_X64Y108_SLICE_X96Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X60Y96_SLICE_X90Y96_AX = CLBLM_R_X59Y96_SLICE_X89Y96_AQ;
  assign CLBLM_L_X60Y96_SLICE_X90Y96_A2 = 1'b1;
  assign CLBLM_L_X60Y96_SLICE_X90Y96_A3 = 1'b1;
  assign CLBLM_L_X60Y96_SLICE_X90Y96_B1 = 1'b1;
  assign CLBLM_L_X64Y108_SLICE_X96Y108_D1 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X60Y96_SLICE_X90Y96_B5 = 1'b1;
  assign CLBLM_L_X64Y108_SLICE_X96Y108_D2 = CLBLM_L_X50Y107_SLICE_X77Y107_AQ;
  assign CLBLM_L_X60Y96_SLICE_X90Y96_B6 = 1'b1;
  assign CLBLM_L_X60Y96_SLICE_X90Y96_B2 = 1'b1;
  assign CLBLM_L_X60Y96_SLICE_X90Y96_B3 = 1'b1;
  assign CLBLM_L_X60Y96_SLICE_X90Y96_BX = CLBLM_R_X59Y96_SLICE_X89Y96_A5Q;
  assign CLBLM_L_X60Y96_SLICE_X90Y96_B4 = 1'b1;
  assign CLBLM_L_X60Y96_SLICE_X90Y96_C1 = 1'b1;
  assign CLBLM_L_X64Y108_SLICE_X96Y108_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X60Y96_SLICE_X90Y96_C2 = 1'b1;
  assign CLBLM_L_X60Y96_SLICE_X90Y96_C3 = 1'b1;
  assign CLBLM_L_X60Y96_SLICE_X90Y96_C4 = 1'b1;
  assign CLBLM_L_X60Y96_SLICE_X90Y96_C5 = 1'b1;
  assign CLBLM_L_X60Y96_SLICE_X90Y96_C6 = 1'b1;
  assign CLBLM_L_X60Y96_SLICE_X90Y96_CE = CLBLL_R_X57Y97_SLICE_X87Y97_AO6;
  assign CLBLM_L_X60Y96_SLICE_X90Y96_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X60Y96_SLICE_X90Y96_D1 = 1'b1;
  assign CLBLM_L_X60Y96_SLICE_X90Y96_D2 = 1'b1;
  assign CLBLM_L_X60Y96_SLICE_X90Y96_D3 = 1'b1;
  assign CLBLM_L_X60Y96_SLICE_X90Y96_D4 = 1'b1;
  assign CLBLM_L_X60Y96_SLICE_X90Y96_D5 = 1'b1;
  assign CLBLM_L_X60Y96_SLICE_X90Y96_D6 = 1'b1;
  assign CLBLM_L_X60Y96_SLICE_X90Y96_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X64Y109_SLICE_X97Y109_A1 = 1'b1;
  assign CLBLM_L_X64Y109_SLICE_X97Y109_A2 = 1'b1;
  assign CLBLM_L_X64Y109_SLICE_X97Y109_A3 = 1'b1;
  assign CLBLM_L_X64Y109_SLICE_X97Y109_A4 = 1'b1;
  assign CLBLM_L_X64Y109_SLICE_X97Y109_A5 = 1'b1;
  assign CLBLM_L_X64Y109_SLICE_X97Y109_A6 = 1'b1;
  assign CLBLM_L_X64Y109_SLICE_X97Y109_B1 = 1'b1;
  assign CLBLM_L_X64Y109_SLICE_X97Y109_B2 = 1'b1;
  assign CLBLM_L_X64Y109_SLICE_X97Y109_B3 = 1'b1;
  assign CLBLM_L_X64Y109_SLICE_X97Y109_B4 = 1'b1;
  assign CLBLM_L_X64Y109_SLICE_X97Y109_B5 = 1'b1;
  assign CLBLM_L_X64Y109_SLICE_X97Y109_B6 = 1'b1;
  assign CLBLM_L_X64Y109_SLICE_X97Y109_C1 = 1'b1;
  assign CLBLM_L_X64Y109_SLICE_X97Y109_C2 = 1'b1;
  assign CLBLM_L_X64Y109_SLICE_X97Y109_C3 = 1'b1;
  assign CLBLM_L_X64Y109_SLICE_X97Y109_C4 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_A1 = CLBLM_L_X50Y106_SLICE_X76Y106_AQ;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_A2 = CLBLM_L_X50Y104_SLICE_X76Y104_AQ;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_A3 = CLBLM_L_X50Y105_SLICE_X77Y105_AQ;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_A4 = CLBLM_L_X50Y107_SLICE_X77Y107_AQ;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_A5 = CLBLM_L_X62Y100_SLICE_X92Y100_AO6;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_A6 = 1'b1;
  assign CLBLM_L_X64Y109_SLICE_X97Y109_C5 = 1'b1;
  assign CLBLM_L_X64Y109_SLICE_X97Y109_C6 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_AX = CLBLM_R_X49Y108_SLICE_X75Y108_DQ;
  assign CLBLL_R_X57Y100_SLICE_X86Y100_A1 = CLBLL_L_X54Y99_SLICE_X82Y99_AQ;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_B1 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_B2 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_B3 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_B4 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_B5 = CLBLM_R_X63Y99_SLICE_X94Y99_DO5;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_B6 = CLBLM_L_X62Y97_SLICE_X92Y97_CQ;
  assign CLBLM_L_X64Y109_SLICE_X97Y109_D1 = 1'b1;
  assign CLBLM_L_X64Y109_SLICE_X97Y109_D2 = 1'b1;
  assign CLBLM_L_X64Y109_SLICE_X97Y109_D3 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_C1 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_C2 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_C3 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_C4 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_C5 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_C6 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_CE = CLBLM_L_X60Y98_SLICE_X91Y98_DQ;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X64Y109_SLICE_X96Y109_A1 = CLBLM_L_X64Y109_SLICE_X96Y109_DO6;
  assign CLBLM_L_X64Y109_SLICE_X96Y109_A2 = CLBLM_R_X49Y106_SLICE_X74Y106_AQ;
  assign CLBLM_L_X64Y109_SLICE_X96Y109_A3 = CLBLM_L_X50Y104_SLICE_X76Y104_AQ;
  assign CLBLM_L_X64Y109_SLICE_X96Y109_A4 = CLBLM_L_X64Y109_SLICE_X96Y109_BO6;
  assign CLBLM_L_X64Y109_SLICE_X96Y109_A5 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_D1 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_D2 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_D3 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_D4 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_D5 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_D6 = 1'b1;
  assign CLBLM_L_X64Y109_SLICE_X96Y109_B1 = CLBLM_R_X63Y109_SLICE_X94Y109_A_XOR;
  assign CLBLM_L_X60Y97_SLICE_X91Y97_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X64Y109_SLICE_X96Y109_B2 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X64Y109_SLICE_X96Y109_B3 = CLBLM_L_X64Y109_SLICE_X96Y109_AQ;
  assign CLBLM_L_X64Y109_SLICE_X96Y109_B4 = CLBLM_L_X62Y105_SLICE_X93Y105_AO6;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_A1 = CLBLM_L_X56Y97_SLICE_X85Y97_DO6;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_A2 = CLBLM_R_X63Y99_SLICE_X94Y99_DO5;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_A3 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_A4 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_A5 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_A6 = 1'b1;
  assign CLBLM_L_X64Y109_SLICE_X96Y109_C1 = CLBLM_L_X62Y105_SLICE_X92Y105_BO5;
  assign CLBLM_L_X64Y109_SLICE_X96Y109_C2 = CLBLM_L_X62Y105_SLICE_X93Y105_AO6;
  assign CLBLM_L_X64Y109_SLICE_X96Y109_C3 = CLBLM_R_X63Y105_SLICE_X94Y105_AQ;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_AX = CLBLM_R_X49Y107_SLICE_X75Y107_DQ;
  assign CLBLM_L_X64Y109_SLICE_X96Y109_C4 = CLBLM_R_X63Y109_SLICE_X95Y109_B_XOR;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_B1 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_B2 = CLBLM_L_X50Y107_SLICE_X76Y107_BQ;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_B4 = CLBLM_R_X49Y105_SLICE_X75Y105_CQ;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_B5 = CLBLM_R_X49Y106_SLICE_X74Y106_AQ;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_B6 = CLBLM_L_X50Y106_SLICE_X76Y106_CQ;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_B3 = CLBLM_L_X60Y97_SLICE_X91Y97_AO6;
  assign CLBLM_L_X64Y109_SLICE_X96Y109_D1 = CLBLM_L_X62Y105_SLICE_X92Y105_BO5;
  assign CLBLM_L_X64Y109_SLICE_X96Y109_D2 = CLBLM_R_X63Y109_SLICE_X94Y109_D_XOR;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_BX = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLM_L_X64Y109_SLICE_X96Y109_D3 = CLBLM_L_X62Y105_SLICE_X93Y105_AO6;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_C1 = CLBLM_L_X60Y97_SLICE_X91Y97_AQ;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_C2 = CLBLM_R_X59Y96_SLICE_X88Y96_AQ;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_C3 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_C4 = CLBLM_L_X60Y97_SLICE_X90Y97_A5Q;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_C5 = CLBLM_R_X59Y96_SLICE_X88Y96_BQ;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_C6 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_CE = CLBLM_L_X60Y98_SLICE_X91Y98_DQ;
  assign CLBLM_L_X64Y109_SLICE_X96Y109_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLL_R_X57Y100_SLICE_X86Y100_B4 = CLBLM_R_X59Y98_SLICE_X89Y98_A5Q;
  assign CLBLL_R_X57Y100_SLICE_X86Y100_B5 = CLBLM_L_X60Y100_SLICE_X90Y100_AO5;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_CX = CLBLM_L_X56Y97_SLICE_X84Y97_CO6;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_D1 = CLBLM_R_X59Y97_SLICE_X88Y97_BQ;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_D2 = CLBLM_L_X60Y97_SLICE_X91Y97_AQ;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_D3 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_D4 = CLBLM_L_X60Y97_SLICE_X90Y97_A5Q;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_D5 = 1'b1;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_D6 = CLBLL_R_X57Y97_SLICE_X86Y97_AQ;
  assign CLBLM_L_X60Y97_SLICE_X90Y97_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLL_R_X57Y100_SLICE_X86Y100_C5 = CLBLL_L_X54Y99_SLICE_X82Y99_CQ;
  assign CLBLL_R_X57Y100_SLICE_X86Y100_C6 = CLBLM_L_X56Y100_SLICE_X85Y100_AQ;
  assign CLBLL_R_X57Y100_SLICE_X86Y100_CE = CLBLL_R_X57Y100_SLICE_X87Y100_DO6;
  assign CLBLL_R_X57Y100_SLICE_X86Y100_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_X0Y117_ILOGIC_X0Y118_D = LIOB33_X0Y117_IOB_X0Y118_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_D = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_C5 = 1'b1;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_C6 = 1'b1;
  assign CLBLM_L_X60Y98_SLICE_X91Y98_A1 = 1'b1;
  assign CLBLM_L_X60Y98_SLICE_X91Y98_A2 = 1'b1;
  assign CLBLM_L_X60Y98_SLICE_X91Y98_A3 = 1'b1;
  assign CLBLM_L_X60Y98_SLICE_X91Y98_A4 = 1'b1;
  assign CLBLM_L_X60Y98_SLICE_X91Y98_A5 = 1'b1;
  assign CLBLM_L_X60Y98_SLICE_X91Y98_A6 = CLBLM_L_X60Y98_SLICE_X91Y98_DQ;
  assign CLBLM_L_X60Y98_SLICE_X91Y98_AX = CLBLM_L_X60Y98_SLICE_X90Y98_CO6;
  assign CLBLM_L_X60Y98_SLICE_X91Y98_B1 = 1'b1;
  assign CLBLM_L_X60Y98_SLICE_X91Y98_B2 = 1'b1;
  assign CLBLM_L_X60Y98_SLICE_X91Y98_B3 = 1'b1;
  assign CLBLM_L_X60Y98_SLICE_X91Y98_B4 = 1'b1;
  assign CLBLM_L_X60Y98_SLICE_X91Y98_B5 = 1'b1;
  assign CLBLM_L_X60Y98_SLICE_X91Y98_B6 = 1'b1;
  assign CLBLM_L_X60Y98_SLICE_X91Y98_BX = CLBLM_L_X60Y98_SLICE_X91Y98_AQ;
  assign CLBLM_L_X60Y98_SLICE_X91Y98_C1 = 1'b1;
  assign CLBLM_L_X60Y98_SLICE_X91Y98_C2 = 1'b1;
  assign CLBLM_L_X60Y98_SLICE_X91Y98_C3 = 1'b1;
  assign CLBLM_L_X60Y98_SLICE_X91Y98_C4 = 1'b1;
  assign CLBLM_L_X60Y98_SLICE_X91Y98_C5 = 1'b1;
  assign CLBLM_L_X60Y98_SLICE_X91Y98_C6 = 1'b1;
  assign CLBLM_L_X60Y98_SLICE_X91Y98_CE = CLBLM_L_X62Y110_SLICE_X93Y110_BO6;
  assign CLBLM_L_X60Y98_SLICE_X91Y98_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X60Y98_SLICE_X91Y98_CX = CLBLM_L_X60Y98_SLICE_X91Y98_BQ;
  assign CLBLM_L_X60Y98_SLICE_X91Y98_D1 = 1'b1;
  assign CLBLM_L_X60Y98_SLICE_X91Y98_D2 = 1'b1;
  assign CLBLM_L_X60Y98_SLICE_X91Y98_D3 = 1'b1;
  assign CLBLM_L_X60Y98_SLICE_X91Y98_D4 = 1'b1;
  assign CLBLM_L_X60Y98_SLICE_X91Y98_D5 = 1'b1;
  assign CLBLM_L_X60Y98_SLICE_X91Y98_D6 = 1'b1;
  assign CLBLM_L_X60Y98_SLICE_X91Y98_DX = CLBLM_L_X60Y98_SLICE_X91Y98_CQ;
  assign CLBLM_L_X60Y98_SLICE_X91Y98_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X60Y98_SLICE_X90Y98_A1 = 1'b1;
  assign CLBLM_L_X60Y98_SLICE_X90Y98_A2 = CLBLM_L_X60Y97_SLICE_X90Y97_CO6;
  assign CLBLM_L_X60Y98_SLICE_X90Y98_A3 = CLBLM_L_X60Y98_SLICE_X90Y98_AQ;
  assign CLBLM_L_X60Y98_SLICE_X90Y98_A4 = CLBLM_L_X60Y97_SLICE_X90Y97_BQ;
  assign CLBLM_L_X60Y98_SLICE_X90Y98_A5 = CLBLM_L_X60Y98_SLICE_X91Y98_AQ;
  assign CLBLM_L_X60Y98_SLICE_X90Y98_A6 = CLBLM_L_X60Y97_SLICE_X90Y97_DO6;
  assign CLBLM_L_X60Y98_SLICE_X90Y98_B1 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X60Y98_SLICE_X90Y98_B2 = CLBLM_L_X60Y98_SLICE_X90Y98_BQ;
  assign CLBLM_L_X60Y98_SLICE_X90Y98_B3 = CLBLM_L_X62Y99_SLICE_X92Y99_AO6;
  assign CLBLM_L_X60Y98_SLICE_X90Y98_B4 = CLBLM_R_X53Y100_SLICE_X80Y100_A5Q;
  assign CLBLM_L_X60Y98_SLICE_X90Y98_B5 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X60Y98_SLICE_X90Y98_B6 = CLBLM_R_X53Y100_SLICE_X80Y100_AQ;
  assign CLBLM_L_X60Y98_SLICE_X90Y98_C1 = CLBLM_R_X53Y100_SLICE_X80Y100_A5Q;
  assign CLBLM_L_X60Y98_SLICE_X90Y98_C2 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X60Y98_SLICE_X90Y98_C3 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X60Y98_SLICE_X90Y98_C4 = CLBLM_R_X53Y100_SLICE_X80Y100_AQ;
  assign CLBLM_L_X60Y98_SLICE_X90Y98_C5 = 1'b1;
  assign CLBLM_L_X60Y98_SLICE_X90Y98_C6 = 1'b1;
  assign CLBLM_L_X60Y98_SLICE_X90Y98_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X60Y98_SLICE_X90Y98_D1 = CLBLM_L_X60Y100_SLICE_X91Y100_CO5;
  assign CLBLM_L_X60Y98_SLICE_X90Y98_D2 = CLBLM_R_X53Y100_SLICE_X80Y100_AQ;
  assign CLBLM_L_X60Y98_SLICE_X90Y98_D3 = CLBLM_L_X62Y104_SLICE_X93Y104_AQ;
  assign CLBLM_L_X60Y98_SLICE_X90Y98_D4 = CLBLM_L_X60Y99_SLICE_X90Y99_AO6;
  assign CLBLM_L_X60Y98_SLICE_X90Y98_D5 = CLBLM_R_X59Y102_SLICE_X89Y102_AQ;
  assign CLBLM_L_X60Y98_SLICE_X90Y98_D6 = CLBLM_R_X53Y100_SLICE_X80Y100_A5Q;
  assign CLBLM_L_X60Y98_SLICE_X90Y98_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_A1 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_A2 = CLBLM_L_X60Y98_SLICE_X90Y98_BQ;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_A3 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_A4 = CLBLM_R_X59Y102_SLICE_X88Y102_AQ;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_A5 = CLBLM_L_X60Y99_SLICE_X91Y99_CO6;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_A6 = 1'b1;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_A4 = CLBLM_R_X65Y103_SLICE_X99Y103_AQ;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_D5 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_B1 = CLBLM_L_X62Y103_SLICE_X92Y103_AQ;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_B2 = CLBLM_L_X60Y110_SLICE_X91Y110_AQ;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_B3 = CLBLM_L_X62Y110_SLICE_X92Y110_DO6;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_B4 = CLBLM_L_X62Y106_SLICE_X93Y106_AQ;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_B5 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_B6 = 1'b1;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_A5 = CLBLM_R_X63Y99_SLICE_X94Y99_CQ;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_A6 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_C1 = CLBLM_L_X62Y106_SLICE_X93Y106_AQ;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_C2 = CLBLM_L_X62Y111_SLICE_X92Y111_BO6;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_C3 = CLBLM_R_X59Y102_SLICE_X89Y102_AQ;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_C4 = CLBLM_L_X62Y103_SLICE_X92Y103_AQ;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_C5 = CLBLM_L_X60Y110_SLICE_X91Y110_AQ;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_C6 = CLBLM_L_X62Y104_SLICE_X93Y104_AQ;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_D6 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_D1 = CLBLM_R_X59Y102_SLICE_X88Y102_AQ;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_D2 = CLBLM_L_X62Y111_SLICE_X92Y111_BO6;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_D3 = CLBLM_R_X59Y102_SLICE_X89Y102_AQ;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_D4 = CLBLM_L_X60Y98_SLICE_X90Y98_BQ;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_D5 = CLBLM_L_X60Y99_SLICE_X91Y99_BO5;
  assign CLBLM_L_X60Y99_SLICE_X91Y99_D6 = CLBLM_L_X62Y104_SLICE_X93Y104_AQ;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_A1 = CLBLM_R_X59Y102_SLICE_X89Y102_AQ;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_A2 = CLBLM_L_X60Y99_SLICE_X91Y99_BO6;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_A3 = CLBLM_R_X59Y102_SLICE_X88Y102_AQ;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_A4 = CLBLM_L_X62Y104_SLICE_X93Y104_AQ;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_A5 = CLBLM_L_X60Y98_SLICE_X90Y98_BQ;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_A6 = 1'b1;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_B3 = CLBLM_L_X50Y104_SLICE_X76Y104_AQ;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_AX = CLBLM_L_X60Y99_SLICE_X90Y99_BO6;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_B1 = CLBLM_L_X60Y110_SLICE_X91Y110_AQ;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_B2 = CLBLM_L_X62Y106_SLICE_X93Y106_AQ;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_B3 = CLBLM_R_X63Y98_SLICE_X94Y98_F7AMUX_O;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_B4 = CLBLM_R_X59Y103_SLICE_X88Y103_CO6;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_B5 = CLBLM_R_X59Y102_SLICE_X89Y102_AQ;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_B6 = 1'b1;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_B5 = CLBLM_R_X65Y98_SLICE_X98Y98_BQ;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_B6 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_C1 = CLBLM_L_X62Y106_SLICE_X93Y106_AQ;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_C2 = CLBLM_R_X63Y97_SLICE_X95Y97_F7AMUX_O;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_C3 = 1'b1;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_C4 = CLBLM_R_X59Y102_SLICE_X88Y102_DO6;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_C5 = CLBLM_R_X59Y102_SLICE_X89Y102_AQ;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_C6 = CLBLM_L_X60Y110_SLICE_X91Y110_AQ;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_CE = CLBLM_L_X62Y99_SLICE_X92Y99_DO6;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_D1 = CLBLM_L_X60Y100_SLICE_X91Y100_CO5;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_D2 = CLBLM_L_X60Y100_SLICE_X91Y100_AO6;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_D3 = CLBLM_R_X59Y100_SLICE_X88Y100_DO6;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_D4 = CLBLM_L_X62Y99_SLICE_X92Y99_AO6;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_D5 = CLBLM_R_X59Y102_SLICE_X89Y102_AQ;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_D6 = CLBLM_L_X62Y104_SLICE_X93Y104_AQ;
  assign CLBLM_L_X60Y99_SLICE_X90Y99_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign LIOI3_X0Y121_ILOGIC_X0Y122_D = LIOB33_X0Y121_IOB_X0Y122_I;
  assign LIOI3_X0Y121_ILOGIC_X0Y121_D = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLM_L_X60Y100_SLICE_X91Y100_A1 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X60Y100_SLICE_X91Y100_A2 = CLBLM_R_X59Y102_SLICE_X88Y102_AQ;
  assign CLBLM_L_X60Y100_SLICE_X91Y100_A3 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X60Y100_SLICE_X91Y100_A4 = CLBLM_L_X60Y98_SLICE_X90Y98_BQ;
  assign CLBLM_L_X60Y100_SLICE_X91Y100_A5 = CLBLM_L_X62Y104_SLICE_X93Y104_AQ;
  assign CLBLM_L_X60Y100_SLICE_X91Y100_A6 = 1'b1;
  assign CLBLM_L_X60Y100_SLICE_X91Y100_B1 = CLBLM_L_X60Y101_SLICE_X91Y101_DO6;
  assign CLBLM_L_X60Y100_SLICE_X91Y100_B2 = CLBLM_R_X63Y99_SLICE_X94Y99_F7AMUX_O;
  assign CLBLM_L_X60Y100_SLICE_X91Y100_B3 = CLBLM_R_X59Y102_SLICE_X89Y102_AQ;
  assign CLBLM_L_X60Y100_SLICE_X91Y100_B4 = CLBLM_L_X60Y110_SLICE_X91Y110_AQ;
  assign CLBLM_L_X60Y100_SLICE_X91Y100_B5 = 1'b1;
  assign CLBLM_L_X60Y100_SLICE_X91Y100_B6 = CLBLM_L_X62Y106_SLICE_X93Y106_AQ;
  assign CLBLM_L_X60Y100_SLICE_X91Y100_C1 = CLBLM_L_X62Y103_SLICE_X92Y103_AQ;
  assign CLBLM_L_X60Y100_SLICE_X91Y100_C2 = CLBLM_L_X62Y106_SLICE_X93Y106_AQ;
  assign CLBLM_L_X60Y100_SLICE_X91Y100_C3 = CLBLM_L_X62Y110_SLICE_X92Y110_DO6;
  assign CLBLM_L_X60Y100_SLICE_X91Y100_C4 = CLBLM_L_X60Y110_SLICE_X91Y110_AQ;
  assign CLBLM_L_X60Y100_SLICE_X91Y100_C5 = 1'b1;
  assign CLBLM_L_X60Y100_SLICE_X91Y100_C6 = 1'b1;
  assign CLBLM_L_X60Y100_SLICE_X91Y100_CE = CLBLM_L_X62Y99_SLICE_X92Y99_DO6;
  assign CLBLM_L_X60Y100_SLICE_X91Y100_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X60Y100_SLICE_X91Y100_D1 = CLBLM_R_X59Y97_SLICE_X88Y97_BQ;
  assign CLBLM_L_X60Y100_SLICE_X91Y100_D2 = CLBLM_L_X62Y107_SLICE_X92Y107_AQ;
  assign CLBLM_L_X60Y100_SLICE_X91Y100_D3 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_L_X60Y100_SLICE_X91Y100_D4 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_L_X60Y100_SLICE_X91Y100_D5 = 1'b1;
  assign CLBLM_L_X60Y100_SLICE_X91Y100_D6 = CLBLM_L_X62Y104_SLICE_X92Y104_AQ;
  assign CLBLM_L_X60Y100_SLICE_X91Y100_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X60Y100_SLICE_X90Y100_A1 = CLBLM_L_X60Y99_SLICE_X90Y99_CQ;
  assign CLBLM_L_X60Y100_SLICE_X90Y100_A2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X60Y100_SLICE_X90Y100_A3 = CLBLM_L_X60Y99_SLICE_X90Y99_AQ;
  assign CLBLM_L_X60Y100_SLICE_X90Y100_A4 = CLBLM_L_X62Y99_SLICE_X92Y99_BQ;
  assign CLBLM_L_X60Y100_SLICE_X90Y100_A5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X60Y100_SLICE_X90Y100_A6 = 1'b1;
  assign CLBLM_L_X60Y100_SLICE_X90Y100_AX = CLBLM_R_X59Y100_SLICE_X88Y100_AO5;
  assign CLBLM_L_X60Y100_SLICE_X90Y100_B1 = CLBLM_R_X59Y101_SLICE_X88Y101_AO6;
  assign CLBLM_L_X60Y100_SLICE_X90Y100_B2 = CLBLM_L_X62Y99_SLICE_X92Y99_AO6;
  assign CLBLM_L_X60Y100_SLICE_X90Y100_B3 = CLBLM_L_X60Y100_SLICE_X91Y100_AO6;
  assign CLBLM_L_X60Y100_SLICE_X90Y100_B4 = CLBLM_L_X60Y100_SLICE_X91Y100_CO5;
  assign CLBLM_L_X60Y100_SLICE_X90Y100_B5 = CLBLM_R_X59Y102_SLICE_X89Y102_AQ;
  assign CLBLM_L_X60Y100_SLICE_X90Y100_B6 = CLBLM_L_X62Y104_SLICE_X93Y104_AQ;
  assign CLBLM_L_X60Y100_SLICE_X90Y100_C1 = CLBLM_R_X59Y102_SLICE_X89Y102_AQ;
  assign CLBLM_L_X60Y100_SLICE_X90Y100_C2 = CLBLM_L_X60Y100_SLICE_X91Y100_AO5;
  assign CLBLM_L_X60Y100_SLICE_X90Y100_C3 = CLBLM_R_X59Y101_SLICE_X88Y101_AO6;
  assign CLBLM_L_X60Y100_SLICE_X90Y100_C4 = CLBLM_L_X62Y99_SLICE_X92Y99_AO6;
  assign CLBLM_L_X60Y100_SLICE_X90Y100_C5 = 1'b1;
  assign CLBLM_L_X60Y100_SLICE_X90Y100_C6 = CLBLM_L_X60Y100_SLICE_X91Y100_CO5;
  assign CLBLM_L_X60Y100_SLICE_X90Y100_CE = CLBLM_L_X60Y99_SLICE_X90Y99_DO6;
  assign CLBLM_L_X60Y100_SLICE_X90Y100_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X60Y100_SLICE_X90Y100_D1 = CLBLM_R_X59Y102_SLICE_X89Y102_AQ;
  assign CLBLM_L_X60Y100_SLICE_X90Y100_D2 = CLBLM_L_X60Y100_SLICE_X91Y100_AO5;
  assign CLBLM_L_X60Y100_SLICE_X90Y100_D3 = CLBLM_L_X60Y100_SLICE_X91Y100_CO5;
  assign CLBLM_L_X60Y100_SLICE_X90Y100_D4 = CLBLM_L_X62Y99_SLICE_X92Y99_AO6;
  assign CLBLM_L_X60Y100_SLICE_X90Y100_D5 = 1'b1;
  assign CLBLM_L_X60Y100_SLICE_X90Y100_D6 = CLBLM_R_X59Y100_SLICE_X88Y100_DO6;
  assign CLBLM_L_X60Y100_SLICE_X90Y100_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_A1 = CLBLM_L_X60Y99_SLICE_X90Y99_BO5;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_A2 = CLBLM_R_X63Y96_SLICE_X95Y96_CO6;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_A3 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_A4 = CLBLM_R_X59Y102_SLICE_X89Y102_BO6;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_A5 = CLBLM_R_X63Y101_SLICE_X95Y101_BO6;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_A6 = CLBLM_L_X62Y106_SLICE_X93Y106_CO6;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_B1 = CLBLM_L_X60Y99_SLICE_X90Y99_BO5;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_B2 = CLBLM_L_X62Y103_SLICE_X93Y103_BO6;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_B3 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_B4 = CLBLM_L_X62Y105_SLICE_X92Y105_DO6;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_B5 = CLBLM_R_X59Y105_SLICE_X89Y105_F7AMUX_O;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_B6 = CLBLM_L_X62Y97_SLICE_X93Y97_F7AMUX_O;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_C1 = CLBLM_L_X62Y99_SLICE_X92Y99_BQ;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_C2 = CLBLM_L_X60Y100_SLICE_X91Y100_BQ;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_C3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_C4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_C5 = CLBLM_L_X60Y101_SLICE_X91Y101_AQ;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_C6 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_CE = CLBLM_L_X62Y99_SLICE_X92Y99_DO6;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_D1 = CLBLL_R_X57Y104_SLICE_X87Y104_DO6;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_D2 = CLBLM_L_X62Y103_SLICE_X93Y103_BO6;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_D3 = CLBLM_L_X64Y105_SLICE_X96Y105_DO6;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_D4 = CLBLM_L_X62Y106_SLICE_X93Y106_CO6;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_D5 = CLBLM_L_X60Y100_SLICE_X91Y100_DO6;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_D6 = CLBLM_R_X59Y101_SLICE_X89Y101_CO6;
  assign CLBLM_L_X60Y101_SLICE_X91Y101_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_A1 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_A2 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_A3 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_A4 = CLBLM_L_X60Y106_SLICE_X91Y106_D_XOR;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_A5 = CLBLM_L_X62Y97_SLICE_X92Y97_AO6;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_A6 = CLBLM_L_X60Y103_SLICE_X91Y103_D_XOR;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_B1 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_B2 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_B3 = CLBLL_L_X54Y101_SLICE_X83Y101_AO6;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_B4 = CLBLM_R_X59Y101_SLICE_X89Y101_BO6;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_B5 = CLBLM_L_X64Y100_SLICE_X97Y100_BQ;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_B6 = CLBLM_L_X64Y100_SLICE_X97Y100_AQ;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_C1 = CLBLM_L_X60Y105_SLICE_X90Y105_C_XOR;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_C2 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_C3 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_C4 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_C5 = CLBLM_R_X59Y105_SLICE_X89Y105_CQ;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_C6 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_CE = CLBLM_L_X62Y102_SLICE_X92Y102_CO6;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_D1 = CLBLM_R_X59Y104_SLICE_X89Y104_CQ;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_D2 = CLBLM_L_X60Y105_SLICE_X90Y105_D_XOR;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_D3 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_D4 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_D5 = 1'b1;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_D6 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X60Y101_SLICE_X90Y101_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_D1 = CLBLM_R_X49Y109_SLICE_X74Y109_DQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_T1 = 1'b1;
  assign CLBLL_R_X57Y101_SLICE_X86Y101_A1 = CLBLM_L_X50Y104_SLICE_X76Y104_AQ;
  assign CLBLL_R_X57Y101_SLICE_X86Y101_A2 = CLBLM_R_X49Y104_SLICE_X74Y104_AQ;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_A1 = 1'b1;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_A2 = CLBLM_L_X60Y102_SLICE_X90Y102_CQ;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_A3 = 1'b1;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_A4 = 1'b1;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_A5 = 1'b1;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_A6 = 1'b1;
  assign CLBLL_R_X57Y101_SLICE_X86Y101_A3 = CLBLL_R_X57Y101_SLICE_X86Y101_AQ;
  assign CLBLL_R_X57Y101_SLICE_X86Y101_A4 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_AX = CLBLM_L_X62Y102_SLICE_X92Y102_BQ;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_B1 = 1'b1;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_B2 = CLBLM_L_X62Y104_SLICE_X92Y104_AQ;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_B3 = 1'b1;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_B4 = CLBLM_L_X62Y102_SLICE_X92Y102_AO6;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_B5 = 1'b1;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_B6 = 1'b1;
  assign CLBLL_R_X57Y101_SLICE_X86Y101_A5 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLL_R_X57Y101_SLICE_X86Y101_A6 = 1'b1;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_BX = CLBLM_L_X62Y104_SLICE_X92Y104_AQ;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_C1 = CLBLM_L_X60Y102_SLICE_X90Y102_AQ;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_C2 = 1'b1;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_C3 = 1'b1;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_C4 = 1'b1;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_C5 = 1'b1;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_C6 = 1'b1;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_CE = CLBLM_L_X62Y102_SLICE_X92Y102_CO6;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_CX = CLBLM_L_X60Y102_SLICE_X90Y102_AQ;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_D1 = 1'b1;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_D2 = 1'b1;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_D3 = 1'b1;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_D4 = 1'b1;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_D5 = 1'b1;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_D6 = CLBLM_L_X60Y102_SLICE_X90Y102_BQ;
  assign CLBLL_R_X57Y101_SLICE_X86Y101_B1 = CLBLL_L_X54Y101_SLICE_X83Y101_CO6;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_DX = CLBLM_L_X60Y102_SLICE_X90Y102_BQ;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLL_R_X57Y101_SLICE_X86Y101_B2 = CLBLM_L_X62Y99_SLICE_X92Y99_AO6;
  assign CLBLM_L_X60Y102_SLICE_X90Y102_A1 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X60Y102_SLICE_X90Y102_A2 = CLBLM_L_X60Y105_SLICE_X91Y105_C_XOR;
  assign CLBLM_L_X60Y102_SLICE_X90Y102_A3 = CLBLM_L_X60Y102_SLICE_X91Y102_C_XOR;
  assign CLBLM_L_X60Y102_SLICE_X90Y102_A4 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X60Y102_SLICE_X90Y102_A5 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X60Y102_SLICE_X90Y102_A6 = CLBLM_L_X62Y98_SLICE_X92Y98_AO6;
  assign CLBLL_R_X57Y101_SLICE_X86Y101_B4 = CLBLL_R_X57Y97_SLICE_X86Y97_CO6;
  assign CLBLM_L_X60Y102_SLICE_X90Y102_B1 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X60Y102_SLICE_X90Y102_B2 = CLBLM_L_X60Y102_SLICE_X91Y102_D_XOR;
  assign CLBLM_L_X60Y102_SLICE_X90Y102_B3 = CLBLM_L_X62Y102_SLICE_X92Y102_AO5;
  assign CLBLM_L_X60Y102_SLICE_X90Y102_B4 = CLBLM_L_X60Y105_SLICE_X91Y105_D_XOR;
  assign CLBLM_L_X60Y102_SLICE_X90Y102_B5 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X60Y102_SLICE_X90Y102_B6 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLL_R_X57Y101_SLICE_X86Y101_B5 = CLBLL_L_X52Y105_SLICE_X78Y105_AO5;
  assign CLBLL_R_X57Y101_SLICE_X86Y101_B6 = CLBLL_R_X57Y101_SLICE_X86Y101_AO5;
  assign CLBLM_L_X60Y102_SLICE_X90Y102_C1 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X60Y102_SLICE_X90Y102_C2 = CLBLM_L_X60Y102_SLICE_X91Y102_A_XOR;
  assign CLBLM_L_X60Y102_SLICE_X90Y102_C3 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X60Y102_SLICE_X90Y102_C4 = CLBLM_L_X60Y105_SLICE_X91Y105_A_XOR;
  assign CLBLM_L_X60Y102_SLICE_X90Y102_C5 = CLBLM_L_X62Y103_SLICE_X93Y103_AO6;
  assign CLBLM_L_X60Y102_SLICE_X90Y102_C6 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X60Y102_SLICE_X90Y102_CE = CLBLM_L_X62Y102_SLICE_X92Y102_DO6;
  assign CLBLM_L_X60Y102_SLICE_X90Y102_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X60Y102_SLICE_X90Y102_D1 = CLBLM_L_X60Y105_SLICE_X91Y105_C_XOR;
  assign CLBLM_L_X60Y102_SLICE_X90Y102_D2 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X60Y102_SLICE_X90Y102_D3 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_L_X60Y102_SLICE_X90Y102_D4 = CLBLM_L_X60Y102_SLICE_X90Y102_AQ;
  assign CLBLM_L_X60Y102_SLICE_X90Y102_D5 = CLBLM_R_X59Y103_SLICE_X89Y103_CQ;
  assign CLBLM_L_X60Y102_SLICE_X90Y102_D6 = CLBLM_L_X60Y101_SLICE_X90Y101_DO6;
  assign CLBLL_R_X57Y101_SLICE_X86Y101_C1 = 1'b1;
  assign LIOI3_X0Y123_ILOGIC_X0Y123_D = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLM_L_X60Y102_SLICE_X90Y102_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLL_R_X57Y101_SLICE_X86Y101_C3 = 1'b1;
  assign CLBLL_R_X57Y101_SLICE_X86Y101_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X57Y101_SLICE_X86Y101_D4 = 1'b1;
  assign CLBLL_R_X57Y101_SLICE_X86Y101_D5 = 1'b1;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_A1 = 1'b1;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_A2 = CLBLM_L_X62Y104_SLICE_X92Y104_BQ;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_A3 = CLBLM_L_X62Y102_SLICE_X92Y102_AO6;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_A4 = 1'b1;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_A5 = 1'b1;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_A6 = 1'b1;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_AX = CLBLM_L_X62Y104_SLICE_X92Y104_BQ;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_B1 = 1'b1;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_B2 = 1'b1;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_B3 = 1'b1;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_B4 = 1'b1;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_B5 = 1'b1;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_B6 = CLBLM_L_X62Y106_SLICE_X92Y106_BQ;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_BX = CLBLM_L_X62Y106_SLICE_X92Y106_BQ;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_C1 = 1'b1;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_C2 = 1'b1;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_C3 = CLBLM_L_X62Y106_SLICE_X92Y106_CQ;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_C4 = 1'b1;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_C5 = 1'b1;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_C6 = 1'b1;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_CE = CLBLM_L_X60Y100_SLICE_X90Y100_DO6;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_CIN = CLBLM_L_X60Y102_SLICE_X91Y102_COUT;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_CX = CLBLM_L_X62Y106_SLICE_X92Y106_CQ;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_D1 = 1'b1;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_D2 = 1'b1;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_D3 = 1'b1;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_D4 = 1'b1;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_D5 = CLBLM_L_X60Y101_SLICE_X90Y101_AQ;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_D6 = 1'b1;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_DX = CLBLM_L_X60Y101_SLICE_X90Y101_AQ;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X60Y103_SLICE_X90Y103_A1 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_L_X60Y103_SLICE_X90Y103_A2 = CLBLM_L_X56Y103_SLICE_X85Y103_BQ;
  assign CLBLM_L_X60Y103_SLICE_X90Y103_A3 = CLBLM_L_X60Y104_SLICE_X91Y104_AQ;
  assign CLBLM_L_X60Y103_SLICE_X90Y103_A4 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_L_X60Y103_SLICE_X90Y103_A5 = CLBLM_L_X56Y103_SLICE_X85Y103_AQ;
  assign CLBLM_L_X60Y103_SLICE_X90Y103_A6 = CLBLL_R_X57Y103_SLICE_X87Y103_AQ;
  assign CLBLM_L_X60Y103_SLICE_X90Y103_AX = CLBLM_L_X62Y106_SLICE_X93Y106_CO6;
  assign CLBLM_L_X60Y103_SLICE_X90Y103_B1 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_L_X60Y103_SLICE_X90Y103_B2 = CLBLM_L_X64Y108_SLICE_X96Y108_AQ;
  assign CLBLM_L_X60Y103_SLICE_X90Y103_B3 = CLBLM_R_X49Y109_SLICE_X74Y109_AQ;
  assign CLBLM_L_X60Y103_SLICE_X90Y103_B4 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_L_X60Y103_SLICE_X90Y103_B5 = 1'b1;
  assign CLBLM_L_X60Y103_SLICE_X90Y103_B6 = CLBLM_R_X63Y104_SLICE_X94Y104_BQ;
  assign CLBLM_L_X60Y103_SLICE_X90Y103_BX = CLBLM_L_X62Y103_SLICE_X93Y103_BO6;
  assign CLBLM_L_X60Y103_SLICE_X90Y103_C1 = CLBLM_R_X59Y96_SLICE_X88Y96_AQ;
  assign CLBLM_L_X60Y103_SLICE_X90Y103_C2 = 1'b1;
  assign CLBLM_L_X60Y103_SLICE_X90Y103_C3 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_L_X60Y103_SLICE_X90Y103_C4 = CLBLM_L_X60Y102_SLICE_X91Y102_BQ;
  assign CLBLM_L_X60Y103_SLICE_X90Y103_C5 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_L_X60Y103_SLICE_X90Y103_C6 = CLBLM_L_X60Y102_SLICE_X90Y102_BQ;
  assign CLBLM_L_X60Y103_SLICE_X90Y103_CX = CLBLM_L_X62Y106_SLICE_X93Y106_CO6;
  assign CLBLM_L_X60Y103_SLICE_X90Y103_D1 = CLBLM_L_X60Y103_SLICE_X91Y103_AQ;
  assign CLBLM_L_X60Y103_SLICE_X90Y103_D2 = CLBLM_R_X59Y98_SLICE_X88Y98_CQ;
  assign CLBLM_L_X60Y103_SLICE_X90Y103_D3 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_L_X60Y103_SLICE_X90Y103_D4 = CLBLM_L_X60Y104_SLICE_X90Y104_AQ;
  assign CLBLM_L_X60Y103_SLICE_X90Y103_D5 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_L_X60Y103_SLICE_X90Y103_D6 = CLBLM_R_X59Y98_SLICE_X89Y98_CQ;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_A1 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_A2 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_A3 = CLBLM_L_X62Y102_SLICE_X92Y102_AO6;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_A4 = CLBLM_L_X60Y109_SLICE_X91Y109_AQ;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_A5 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_A6 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_D1 = CLBLM_R_X49Y111_SLICE_X74Y111_AQ;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_AX = CLBLM_L_X60Y109_SLICE_X91Y109_AQ;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_B1 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_B2 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_B3 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_B4 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_B5 = CLBLM_L_X62Y107_SLICE_X92Y107_AQ;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_B6 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_T1 = 1'b1;
  assign CLBLM_R_X63Y100_SLICE_X95Y100_A4 = CLBLM_R_X65Y105_SLICE_X98Y105_BQ;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_BX = CLBLM_L_X62Y107_SLICE_X92Y107_AQ;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_C1 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_C2 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_C3 = 1'b1;
  assign CLBLM_R_X63Y100_SLICE_X95Y100_A5 = CLBLM_R_X65Y105_SLICE_X99Y105_AQ;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_C4 = CLBLM_L_X60Y109_SLICE_X91Y109_BQ;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_C5 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_C6 = 1'b1;
  assign CLBLM_R_X63Y100_SLICE_X95Y100_A6 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_CE = CLBLM_L_X60Y100_SLICE_X90Y100_CO6;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_CIN = CLBLM_L_X60Y103_SLICE_X91Y103_COUT;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_D1 = CLBLM_R_X49Y107_SLICE_X74Y107_AQ;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_CX = 1'b0;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_D1 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_D2 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_D3 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_D4 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_D5 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_D6 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_T1 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_DX = 1'b0;
  assign CLBLM_L_X60Y104_SLICE_X91Y104_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_A1 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_A2 = CLBLM_R_X59Y107_SLICE_X89Y107_D_XOR;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_A3 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_A4 = CLBLM_L_X62Y102_SLICE_X92Y102_AO5;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_A5 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_A6 = CLBLM_L_X60Y108_SLICE_X90Y108_D_XOR;
  assign CLBLM_R_X63Y100_SLICE_X95Y100_B2 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_B1 = CLBLM_L_X60Y104_SLICE_X90Y104_DO6;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_B2 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_B3 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_R_X63Y100_SLICE_X95Y100_B3 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_B4 = CLBLM_L_X60Y102_SLICE_X90Y102_CQ;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_B5 = CLBLM_R_X59Y103_SLICE_X89Y103_CQ;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_B6 = CLBLM_L_X60Y105_SLICE_X91Y105_A_XOR;
  assign CLBLM_R_X63Y100_SLICE_X95Y100_B4 = CLBLM_L_X62Y100_SLICE_X92Y100_CQ;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_C1 = CLBLM_L_X60Y106_SLICE_X90Y106_AQ;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_C2 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_R_X63Y100_SLICE_X95Y100_B5 = CLBLM_L_X64Y100_SLICE_X97Y100_D_XOR;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_C3 = CLBLM_R_X59Y98_SLICE_X89Y98_C5Q;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_C4 = CLBLM_R_X59Y100_SLICE_X89Y100_BQ;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_C5 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_C6 = CLBLM_R_X59Y112_SLICE_X89Y112_AQ;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_CE = CLBLM_L_X60Y99_SLICE_X90Y99_DO6;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_D1 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_D2 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_D3 = CLBLM_L_X60Y105_SLICE_X90Y105_B_XOR;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_D4 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_D5 = CLBLM_R_X59Y106_SLICE_X89Y106_CQ;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_D6 = 1'b1;
  assign CLBLM_L_X60Y104_SLICE_X90Y104_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X60Y110_SLICE_X90Y110_B5 = 1'b1;
  assign CLBLM_L_X60Y110_SLICE_X90Y110_B6 = CLBLM_R_X59Y111_SLICE_X89Y111_BQ;
  assign CLBLM_L_X60Y110_SLICE_X90Y110_BX = 1'b0;
  assign CLBLM_L_X60Y110_SLICE_X90Y110_C1 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X91Y105_A1 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X91Y105_A2 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X91Y105_A3 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X91Y105_A4 = CLBLM_L_X60Y102_SLICE_X90Y102_CQ;
  assign CLBLM_L_X60Y105_SLICE_X91Y105_A5 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X91Y105_A6 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X91Y105_AX = CLBLM_L_X62Y102_SLICE_X92Y102_BQ;
  assign CLBLM_L_X60Y105_SLICE_X91Y105_B1 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X91Y105_B2 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X91Y105_B3 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X91Y105_B4 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X91Y105_B5 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X91Y105_B6 = CLBLM_L_X62Y104_SLICE_X92Y104_AQ;
  assign CLBLM_L_X60Y105_SLICE_X91Y105_BX = 1'b0;
  assign CLBLM_L_X60Y105_SLICE_X91Y105_C1 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X91Y105_C2 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X91Y105_C3 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X91Y105_C4 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X91Y105_C5 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X91Y105_C6 = CLBLM_L_X60Y102_SLICE_X90Y102_AQ;
  assign CLBLM_L_X60Y110_SLICE_X90Y110_D4 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X91Y105_CX = 1'b0;
  assign CLBLM_L_X60Y105_SLICE_X91Y105_D1 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X91Y105_D2 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X91Y105_D3 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X91Y105_D4 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X91Y105_D5 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X91Y105_D6 = CLBLM_L_X60Y102_SLICE_X90Y102_BQ;
  assign CLBLM_L_X60Y105_SLICE_X91Y105_DX = 1'b0;
  assign CLBLM_L_X60Y105_SLICE_X90Y105_A1 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X90Y105_A2 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X90Y105_A3 = CLBLM_L_X62Y102_SLICE_X92Y102_BQ;
  assign CLBLM_L_X60Y105_SLICE_X90Y105_A4 = CLBLM_R_X59Y98_SLICE_X89Y98_AQ;
  assign CLBLM_L_X60Y105_SLICE_X90Y105_A5 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X90Y105_A6 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X90Y105_AX = CLBLM_L_X62Y102_SLICE_X92Y102_BQ;
  assign CLBLM_L_X60Y105_SLICE_X90Y105_B1 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X90Y105_B2 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X90Y105_B3 = CLBLM_L_X60Y102_SLICE_X90Y102_CQ;
  assign CLBLM_L_X60Y105_SLICE_X90Y105_B4 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X90Y105_B5 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X90Y105_B6 = CLBLM_R_X59Y98_SLICE_X89Y98_A5Q;
  assign CLBLM_L_X60Y105_SLICE_X90Y105_BX = CLBLM_L_X60Y102_SLICE_X90Y102_CQ;
  assign CLBLM_L_X60Y105_SLICE_X90Y105_C1 = CLBLM_R_X59Y98_SLICE_X89Y98_BQ;
  assign CLBLM_L_X60Y105_SLICE_X90Y105_C2 = CLBLM_L_X62Y104_SLICE_X92Y104_AQ;
  assign CLBLM_L_X60Y105_SLICE_X90Y105_C3 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X90Y105_C4 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X90Y105_C5 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X90Y105_C6 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X47Y119_A1 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X47Y119_A6 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X47Y119_A2 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X47Y119_A3 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X47Y119_A4 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X47Y119_A5 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X47Y119_B1 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X90Y105_CX = CLBLM_L_X62Y104_SLICE_X92Y104_AQ;
  assign CLBLM_L_X32Y119_SLICE_X47Y119_B2 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X90Y105_D1 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X90Y105_D2 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X90Y105_D3 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X90Y105_D4 = CLBLM_R_X59Y98_SLICE_X89Y98_B5Q;
  assign CLBLM_L_X60Y105_SLICE_X90Y105_D5 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X90Y105_D6 = CLBLM_L_X60Y102_SLICE_X90Y102_AQ;
  assign CLBLM_L_X32Y119_SLICE_X47Y119_B3 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X47Y119_B4 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X47Y119_B5 = 1'b1;
  assign CLBLM_L_X60Y105_SLICE_X90Y105_DX = CLBLM_L_X60Y102_SLICE_X90Y102_AQ;
  assign CLBLM_L_X32Y119_SLICE_X47Y119_B6 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X47Y119_C1 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X47Y119_C2 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X47Y119_C3 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X47Y119_C4 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X47Y119_C5 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X47Y119_C6 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X47Y119_D1 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X47Y119_D2 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X47Y119_D3 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X47Y119_D4 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X47Y119_D5 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X47Y119_D6 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X46Y119_A1 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X46Y119_A2 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X46Y119_A3 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X46Y119_A4 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X46Y119_A5 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X46Y119_A6 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X46Y119_AX = LIOB33_X0Y119_IOB_X0Y119_I;
  assign CLBLM_L_X32Y119_SLICE_X46Y119_B1 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X46Y119_B2 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X46Y119_B3 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X46Y119_B4 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X46Y119_B5 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X46Y119_B6 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X46Y119_BX = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_L_X32Y119_SLICE_X46Y119_C1 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X46Y119_C2 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X46Y119_C3 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X46Y119_C4 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X46Y119_C5 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X46Y119_C6 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X46Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X32Y119_SLICE_X46Y119_D1 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X46Y119_D2 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X46Y119_D3 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X46Y119_D4 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X46Y119_D5 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X46Y119_D6 = 1'b1;
  assign CLBLM_L_X32Y119_SLICE_X46Y119_SR = CLBLM_R_X15Y122_SLICE_X20Y122_AO6;
  assign CLBLM_L_X60Y106_SLICE_X91Y106_A1 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X91Y106_A2 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X91Y106_A3 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X91Y106_A4 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X91Y106_A5 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X91Y106_A6 = CLBLM_L_X62Y104_SLICE_X92Y104_BQ;
  assign CLBLM_L_X60Y106_SLICE_X91Y106_AX = 1'b0;
  assign CLBLM_L_X60Y106_SLICE_X91Y106_B1 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X91Y106_B2 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X91Y106_B3 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X91Y106_B4 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X91Y106_B5 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X91Y106_B6 = CLBLM_L_X62Y106_SLICE_X92Y106_BQ;
  assign CLBLM_L_X60Y106_SLICE_X91Y106_BX = 1'b0;
  assign CLBLM_L_X60Y106_SLICE_X91Y106_C1 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X91Y106_C2 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X91Y106_C3 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X91Y106_C4 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X91Y106_C5 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X91Y106_C6 = CLBLM_L_X62Y106_SLICE_X92Y106_CQ;
  assign CLBLM_L_X60Y106_SLICE_X91Y106_CIN = CLBLM_L_X60Y105_SLICE_X91Y105_COUT;
  assign CLBLM_L_X60Y106_SLICE_X91Y106_CX = 1'b0;
  assign CLBLM_L_X60Y106_SLICE_X91Y106_D1 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X91Y106_D2 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X91Y106_D3 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X91Y106_D4 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X91Y106_D5 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X91Y106_D6 = CLBLM_L_X60Y101_SLICE_X90Y101_AQ;
  assign CLBLM_L_X60Y106_SLICE_X91Y106_DX = 1'b0;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_A1 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_A2 = CLBLM_R_X59Y98_SLICE_X89Y98_CQ;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_A3 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_A4 = CLBLM_L_X62Y106_SLICE_X93Y106_BO6;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_A5 = CLBLM_L_X60Y102_SLICE_X90Y102_BQ;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_A6 = 1'b1;
  assign CLBLM_R_X65Y96_SLICE_X99Y96_A1 = 1'b1;
  assign CLBLM_R_X65Y96_SLICE_X99Y96_A2 = 1'b1;
  assign CLBLM_R_X65Y96_SLICE_X99Y96_A3 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_AX = CLBLM_L_X60Y102_SLICE_X90Y102_BQ;
  assign CLBLM_R_X65Y96_SLICE_X99Y96_A4 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_B1 = CLBLM_L_X62Y104_SLICE_X92Y104_BQ;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_B2 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_B3 = CLBLM_R_X59Y98_SLICE_X89Y98_C5Q;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_B4 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_B5 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_B6 = 1'b1;
  assign CLBLM_R_X65Y96_SLICE_X99Y96_A5 = 1'b1;
  assign CLBLM_R_X65Y96_SLICE_X99Y96_A6 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_BX = CLBLM_L_X62Y104_SLICE_X92Y104_BQ;
  assign CLBLM_R_X65Y96_SLICE_X99Y96_B1 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_C1 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_C2 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_C3 = CLBLM_R_X59Y96_SLICE_X89Y96_AQ;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_C4 = CLBLM_L_X62Y106_SLICE_X92Y106_BQ;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_C5 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_C6 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_CE = CLBLM_L_X60Y100_SLICE_X90Y100_DO6;
  assign CLBLM_R_X65Y96_SLICE_X99Y96_B5 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_CIN = CLBLM_L_X60Y105_SLICE_X90Y105_COUT;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X65Y96_SLICE_X99Y96_C1 = 1'b1;
  assign CLBLM_R_X65Y96_SLICE_X99Y96_C2 = 1'b1;
  assign CLBLM_R_X65Y96_SLICE_X99Y96_C3 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_CX = CLBLM_L_X62Y106_SLICE_X92Y106_BQ;
  assign CLBLM_R_X65Y96_SLICE_X99Y96_C4 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_D1 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_D2 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_D3 = CLBLM_L_X62Y106_SLICE_X92Y106_CQ;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_D4 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_D5 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_D6 = CLBLM_R_X59Y96_SLICE_X89Y96_A5Q;
  assign CLBLM_R_X65Y96_SLICE_X99Y96_D1 = 1'b1;
  assign CLBLM_R_X65Y96_SLICE_X99Y96_D2 = 1'b1;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_DX = CLBLM_L_X62Y106_SLICE_X92Y106_CQ;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X65Y96_SLICE_X99Y96_D3 = 1'b1;
  assign CLBLM_R_X65Y96_SLICE_X99Y96_D4 = 1'b1;
  assign CLBLM_R_X65Y96_SLICE_X99Y96_D5 = 1'b1;
  assign CLBLM_R_X65Y96_SLICE_X99Y96_D6 = 1'b1;
  assign CLBLM_R_X65Y96_SLICE_X98Y96_A1 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X65Y96_SLICE_X98Y96_A2 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_R_X65Y96_SLICE_X98Y96_A3 = CLBLM_L_X56Y97_SLICE_X85Y97_AQ;
  assign CLBLM_R_X65Y96_SLICE_X98Y96_A4 = CLBLM_R_X63Y95_SLICE_X95Y95_CQ;
  assign CLBLM_R_X65Y96_SLICE_X98Y96_A5 = 1'b1;
  assign CLBLM_R_X65Y96_SLICE_X98Y96_A6 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_R_X65Y96_SLICE_X98Y96_B1 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X65Y96_SLICE_X98Y96_B2 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_R_X65Y96_SLICE_X98Y96_B3 = CLBLM_L_X56Y97_SLICE_X85Y97_AQ;
  assign CLBLM_R_X65Y96_SLICE_X98Y96_B4 = 1'b1;
  assign CLBLM_R_X65Y96_SLICE_X98Y96_B5 = CLBLM_R_X63Y95_SLICE_X95Y95_D5Q;
  assign CLBLM_R_X65Y96_SLICE_X98Y96_B6 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_D1 = CLBLM_R_X49Y109_SLICE_X74Y109_AQ;
  assign CLBLM_R_X65Y96_SLICE_X98Y96_C1 = 1'b1;
  assign CLBLM_R_X65Y96_SLICE_X98Y96_C2 = 1'b1;
  assign CLBLM_R_X65Y96_SLICE_X98Y96_C3 = 1'b1;
  assign CLBLM_R_X65Y96_SLICE_X98Y96_C4 = 1'b1;
  assign CLBLM_R_X65Y96_SLICE_X98Y96_C5 = 1'b1;
  assign CLBLM_R_X65Y96_SLICE_X98Y96_C6 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_T1 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_D1 = CLBLM_R_X49Y111_SLICE_X74Y111_BQ;
  assign CLBLM_R_X65Y96_SLICE_X98Y96_D1 = 1'b1;
  assign CLBLM_R_X65Y96_SLICE_X98Y96_D2 = 1'b1;
  assign CLBLM_R_X65Y96_SLICE_X98Y96_D3 = 1'b1;
  assign CLBLM_R_X65Y96_SLICE_X98Y96_D4 = 1'b1;
  assign CLBLM_R_X65Y96_SLICE_X98Y96_D5 = 1'b1;
  assign CLBLM_R_X65Y96_SLICE_X98Y96_D6 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_T1 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_A1 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_A2 = CLBLM_L_X62Y107_SLICE_X92Y107_BO6;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_A3 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_A4 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_A5 = CLBLM_L_X60Y109_SLICE_X91Y109_AQ;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_A6 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_AX = 1'b0;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_B1 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_B2 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_B3 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_B4 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_B5 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_B6 = CLBLM_L_X62Y107_SLICE_X92Y107_AQ;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_BX = 1'b0;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_C1 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_C2 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_C3 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_C4 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_C5 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_C6 = CLBLM_L_X60Y109_SLICE_X91Y109_BQ;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_CE = CLBLM_L_X60Y100_SLICE_X90Y100_DO6;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_CIN = CLBLM_L_X60Y106_SLICE_X91Y106_COUT;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_CX = 1'b0;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_D1 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_D2 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_D3 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_D4 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_D5 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_D6 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_DX = 1'b0;
  assign CLBLM_L_X60Y107_SLICE_X91Y107_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_A1 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_A2 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_A3 = CLBLM_L_X60Y101_SLICE_X90Y101_AQ;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_A4 = CLBLM_L_X62Y107_SLICE_X92Y107_BO6;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_A5 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_A6 = 1'b1;
  assign CLBLM_R_X65Y97_SLICE_X99Y97_A1 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X65Y97_SLICE_X99Y97_A2 = 1'b1;
  assign CLBLM_R_X65Y97_SLICE_X99Y97_A3 = CLBLM_L_X56Y97_SLICE_X85Y97_AQ;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_AX = 1'b0;
  assign CLBLM_R_X65Y97_SLICE_X99Y97_A4 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_B1 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_B2 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_B3 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_B4 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_B5 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_B6 = CLBLM_L_X60Y109_SLICE_X91Y109_AQ;
  assign CLBLM_R_X65Y97_SLICE_X99Y97_A5 = CLBLM_L_X62Y96_SLICE_X93Y96_DQ;
  assign CLBLM_R_X65Y97_SLICE_X99Y97_A6 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_BX = 1'b0;
  assign CLBLM_R_X65Y97_SLICE_X99Y97_B1 = CLBLM_L_X62Y96_SLICE_X93Y96_CQ;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_C1 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_C2 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_C3 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_C4 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_C5 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_C6 = CLBLM_L_X62Y107_SLICE_X92Y107_AQ;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_CE = CLBLM_L_X60Y100_SLICE_X90Y100_CO6;
  assign CLBLM_R_X65Y97_SLICE_X99Y97_B5 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_CIN = CLBLM_L_X60Y106_SLICE_X90Y106_COUT;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X65Y97_SLICE_X99Y97_C1 = CLBLM_L_X56Y97_SLICE_X85Y97_AQ;
  assign CLBLM_R_X65Y97_SLICE_X99Y97_C2 = 1'b1;
  assign CLBLM_R_X65Y97_SLICE_X99Y97_C3 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_CX = 1'b0;
  assign CLBLM_R_X65Y97_SLICE_X99Y97_C4 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_D1 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_D2 = 1'b1;
  assign CLBLM_R_X65Y97_SLICE_X99Y97_D1 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_D5 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_D6 = CLBLM_L_X60Y109_SLICE_X91Y109_BQ;
  assign CLBLM_R_X65Y97_SLICE_X99Y97_D4 = 1'b1;
  assign CLBLM_R_X65Y97_SLICE_X99Y97_D5 = 1'b1;
  assign CLBLM_R_X65Y97_SLICE_X99Y97_D6 = 1'b1;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_DX = 1'b0;
  assign CLBLM_L_X60Y107_SLICE_X90Y107_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X65Y97_SLICE_X99Y97_D2 = 1'b1;
  assign CLBLM_R_X65Y97_SLICE_X99Y97_D3 = 1'b1;
  assign CLBLM_R_X65Y97_SLICE_X98Y97_A1 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X65Y97_SLICE_X98Y97_A2 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_R_X65Y97_SLICE_X98Y97_A3 = CLBLM_L_X60Y98_SLICE_X90Y98_AQ;
  assign CLBLM_R_X65Y97_SLICE_X98Y97_A4 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_R_X65Y97_SLICE_X98Y97_A5 = CLBLM_L_X56Y97_SLICE_X85Y97_AQ;
  assign CLBLM_R_X65Y97_SLICE_X98Y97_A6 = 1'b1;
  assign CLBLM_R_X47Y119_SLICE_X73Y119_A1 = CLBLM_R_X47Y119_SLICE_X73Y119_CQ;
  assign CLBLM_R_X47Y119_SLICE_X73Y119_A2 = 1'b1;
  assign CLBLM_R_X65Y97_SLICE_X98Y97_B1 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X47Y119_SLICE_X73Y119_A3 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLM_R_X47Y119_SLICE_X73Y119_A4 = CLBLM_R_X47Y119_SLICE_X73Y119_DQ;
  assign CLBLM_R_X47Y119_SLICE_X73Y119_A5 = CLBLM_L_X32Y119_SLICE_X46Y119_BQ;
  assign CLBLM_R_X47Y119_SLICE_X73Y119_A6 = 1'b1;
  assign CLBLM_R_X65Y97_SLICE_X98Y97_B4 = CLBLM_L_X64Y97_SLICE_X97Y97_AQ;
  assign CLBLM_R_X65Y97_SLICE_X98Y97_B2 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_R_X65Y97_SLICE_X98Y97_B3 = CLBLM_L_X56Y97_SLICE_X85Y97_AQ;
  assign CLBLM_R_X47Y119_SLICE_X73Y119_AX = CLBLM_L_X32Y119_SLICE_X46Y119_AQ;
  assign CLBLM_R_X47Y119_SLICE_X73Y119_B1 = 1'b1;
  assign CLBLM_R_X47Y119_SLICE_X73Y119_B2 = CLBLM_R_X47Y119_SLICE_X73Y119_BQ;
  assign CLBLM_R_X47Y119_SLICE_X73Y119_B3 = CLBLM_R_X47Y119_SLICE_X73Y119_AQ;
  assign CLBLM_R_X47Y119_SLICE_X73Y119_B4 = CLBLM_L_X32Y119_SLICE_X46Y119_AQ;
  assign CLBLM_R_X47Y119_SLICE_X73Y119_B5 = 1'b1;
  assign CLBLM_R_X47Y119_SLICE_X73Y119_B6 = 1'b1;
  assign CLBLM_R_X47Y119_SLICE_X73Y119_BX = CLBLM_R_X47Y119_SLICE_X73Y119_AQ;
  assign CLBLM_R_X47Y119_SLICE_X73Y119_C1 = 1'b1;
  assign CLBLM_R_X47Y119_SLICE_X73Y119_C2 = 1'b1;
  assign CLBLM_R_X47Y119_SLICE_X73Y119_C3 = 1'b1;
  assign CLBLM_R_X47Y119_SLICE_X73Y119_C4 = 1'b1;
  assign CLBLM_R_X47Y119_SLICE_X73Y119_C5 = 1'b1;
  assign CLBLM_R_X65Y97_SLICE_X98Y97_C3 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X65Y97_SLICE_X98Y97_C4 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_R_X65Y97_SLICE_X98Y97_C5 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_R_X47Y119_SLICE_X73Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X65Y97_SLICE_X98Y97_D1 = CLBLM_L_X56Y97_SLICE_X85Y97_AQ;
  assign CLBLM_R_X65Y97_SLICE_X98Y97_D2 = 1'b1;
  assign CLBLM_R_X65Y97_SLICE_X98Y97_D3 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_R_X47Y119_SLICE_X73Y119_CX = CLBLM_L_X32Y119_SLICE_X46Y119_BQ;
  assign CLBLM_R_X65Y97_SLICE_X98Y97_D4 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_R_X47Y119_SLICE_X73Y119_D1 = 1'b1;
  assign CLBLM_R_X47Y119_SLICE_X73Y119_D2 = 1'b1;
  assign CLBLM_R_X47Y119_SLICE_X73Y119_D3 = 1'b1;
  assign CLBLM_R_X47Y119_SLICE_X73Y119_D4 = 1'b1;
  assign CLBLM_R_X47Y119_SLICE_X73Y119_D5 = 1'b1;
  assign CLBLM_R_X47Y119_SLICE_X73Y119_D6 = 1'b1;
  assign CLBLM_R_X65Y97_SLICE_X98Y97_D5 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X47Y119_SLICE_X73Y119_DX = CLBLM_R_X47Y119_SLICE_X73Y119_CQ;
  assign CLBLM_R_X47Y119_SLICE_X73Y119_SR = CLBLM_R_X15Y122_SLICE_X20Y122_AO6;
  assign CLBLM_R_X47Y119_SLICE_X72Y119_A1 = 1'b1;
  assign CLBLM_R_X47Y119_SLICE_X72Y119_A2 = 1'b1;
  assign CLBLM_R_X47Y119_SLICE_X72Y119_A3 = 1'b1;
  assign CLBLM_R_X47Y119_SLICE_X72Y119_A4 = 1'b1;
  assign CLBLM_R_X47Y119_SLICE_X72Y119_A5 = 1'b1;
  assign CLBLM_R_X47Y119_SLICE_X72Y119_A6 = 1'b1;
  assign CLBLM_R_X47Y119_SLICE_X72Y119_B1 = 1'b1;
  assign CLBLM_R_X47Y119_SLICE_X72Y119_B2 = 1'b1;
  assign CLBLM_R_X47Y119_SLICE_X72Y119_B3 = 1'b1;
  assign CLBLM_R_X47Y119_SLICE_X72Y119_B4 = 1'b1;
  assign CLBLM_R_X47Y119_SLICE_X72Y119_B5 = 1'b1;
  assign CLBLM_R_X47Y119_SLICE_X72Y119_B6 = 1'b1;
  assign CLBLM_R_X47Y119_SLICE_X72Y119_C1 = 1'b1;
  assign CLBLM_R_X47Y119_SLICE_X72Y119_C2 = 1'b1;
  assign CLBLM_R_X47Y119_SLICE_X72Y119_C3 = 1'b1;
  assign CLBLM_R_X47Y119_SLICE_X72Y119_C4 = 1'b1;
  assign CLBLM_R_X47Y119_SLICE_X72Y119_C5 = 1'b1;
  assign CLBLM_R_X47Y119_SLICE_X72Y119_C6 = 1'b1;
  assign CLBLM_R_X47Y119_SLICE_X72Y119_D1 = 1'b1;
  assign CLBLM_R_X47Y119_SLICE_X72Y119_D2 = 1'b1;
  assign CLBLM_R_X47Y119_SLICE_X72Y119_D3 = 1'b1;
  assign CLBLM_R_X47Y119_SLICE_X72Y119_D4 = 1'b1;
  assign CLBLM_R_X47Y119_SLICE_X72Y119_D5 = 1'b1;
  assign CLBLM_R_X47Y119_SLICE_X72Y119_D6 = 1'b1;
  assign CLBLM_L_X60Y108_SLICE_X91Y108_A1 = CLBLL_R_X57Y106_SLICE_X87Y106_D_XOR;
  assign CLBLM_L_X60Y108_SLICE_X91Y108_A2 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X60Y108_SLICE_X91Y108_A3 = CLBLM_L_X62Y97_SLICE_X92Y97_AO6;
  assign CLBLM_L_X60Y108_SLICE_X91Y108_A4 = CLBLL_R_X57Y107_SLICE_X86Y107_D_XOR;
  assign CLBLM_L_X60Y108_SLICE_X91Y108_A5 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X60Y108_SLICE_X91Y108_A6 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X60Y108_SLICE_X91Y108_B1 = CLBLM_L_X62Y106_SLICE_X92Y106_AO5;
  assign CLBLM_L_X60Y108_SLICE_X91Y108_B2 = CLBLL_R_X57Y108_SLICE_X87Y108_CO6;
  assign CLBLM_L_X60Y108_SLICE_X91Y108_B3 = CLBLL_R_X57Y105_SLICE_X86Y105_AQ;
  assign CLBLM_L_X60Y108_SLICE_X91Y108_B4 = CLBLM_R_X59Y108_SLICE_X88Y108_C_XOR;
  assign CLBLM_L_X60Y108_SLICE_X91Y108_B5 = CLBLM_L_X60Y108_SLICE_X90Y108_B_XOR;
  assign CLBLM_L_X60Y108_SLICE_X91Y108_B6 = CLBLM_R_X59Y106_SLICE_X89Y106_AO6;
  assign CLBLM_L_X60Y108_SLICE_X91Y108_C1 = CLBLM_L_X60Y105_SLICE_X91Y105_D_XOR;
  assign CLBLM_L_X60Y108_SLICE_X91Y108_C2 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X60Y108_SLICE_X91Y108_C3 = CLBLM_R_X59Y103_SLICE_X89Y103_CQ;
  assign CLBLM_L_X60Y108_SLICE_X91Y108_C4 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_L_X60Y108_SLICE_X91Y108_C5 = CLBLM_L_X60Y102_SLICE_X90Y102_BQ;
  assign CLBLM_L_X60Y108_SLICE_X91Y108_C6 = CLBLM_R_X59Y106_SLICE_X89Y106_AO5;
  assign CLBLM_L_X60Y108_SLICE_X91Y108_CE = CLBLM_L_X60Y100_SLICE_X90Y100_CO6;
  assign CLBLM_L_X60Y108_SLICE_X91Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X60Y108_SLICE_X91Y108_D1 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_L_X60Y108_SLICE_X91Y108_D2 = CLBLL_R_X57Y106_SLICE_X86Y106_D_XOR;
  assign CLBLM_L_X60Y108_SLICE_X91Y108_D3 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X60Y108_SLICE_X91Y108_D4 = CLBLL_R_X57Y103_SLICE_X87Y103_AQ;
  assign CLBLM_L_X60Y108_SLICE_X91Y108_D5 = CLBLL_R_X57Y110_SLICE_X87Y110_A_XOR;
  assign CLBLM_L_X60Y108_SLICE_X91Y108_D6 = CLBLM_R_X59Y107_SLICE_X89Y107_BQ;
  assign CLBLM_L_X60Y108_SLICE_X91Y108_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_A1 = 1'b1;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_A2 = 1'b1;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_A3 = CLBLM_R_X59Y106_SLICE_X89Y106_CQ;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_A4 = 1'b1;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_A5 = 1'b1;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_A6 = 1'b1;
  assign CLBLM_R_X65Y98_SLICE_X99Y98_A1 = CLBLM_R_X65Y98_SLICE_X99Y98_DO6;
  assign CLBLM_R_X65Y98_SLICE_X99Y98_A2 = 1'b1;
  assign CLBLM_R_X65Y98_SLICE_X99Y98_A3 = CLBLM_R_X65Y98_SLICE_X98Y98_CO6;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_AX = CLBLM_L_X60Y100_SLICE_X90Y100_AQ;
  assign CLBLM_R_X65Y98_SLICE_X99Y98_A4 = CLBLM_R_X65Y98_SLICE_X99Y98_BO6;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_B1 = 1'b1;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_B2 = CLBLM_R_X59Y105_SLICE_X89Y105_CQ;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_B3 = 1'b1;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_B4 = CLBLM_L_X62Y108_SLICE_X92Y108_BO6;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_B5 = 1'b1;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_B6 = 1'b1;
  assign CLBLM_R_X65Y98_SLICE_X99Y98_B2 = CLBLM_L_X60Y98_SLICE_X90Y98_AQ;
  assign CLBLM_R_X65Y98_SLICE_X99Y98_B3 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_R_X65Y98_SLICE_X99Y98_B4 = CLBLM_L_X64Y100_SLICE_X96Y100_D_XOR;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_BX = 1'b0;
  assign CLBLM_R_X65Y98_SLICE_X99Y98_B5 = CLBLM_L_X56Y97_SLICE_X85Y97_AQ;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_C1 = 1'b1;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_C2 = 1'b1;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_C3 = 1'b1;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_C4 = 1'b1;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_C5 = 1'b1;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_C6 = CLBLM_R_X59Y104_SLICE_X89Y104_CQ;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_CE = CLBLM_L_X62Y102_SLICE_X92Y102_CO6;
  assign CLBLM_R_X65Y98_SLICE_X99Y98_B6 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X65Y98_SLICE_X99Y98_C1 = CLBLM_L_X64Y102_SLICE_X97Y102_D_XOR;
  assign CLBLM_R_X65Y98_SLICE_X99Y98_C2 = CLBLM_R_X49Y104_SLICE_X75Y104_CQ;
  assign CLBLM_R_X65Y98_SLICE_X99Y98_C3 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_R_X65Y98_SLICE_X99Y98_C4 = 1'b1;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_CX = 1'b0;
  assign CLBLM_R_X65Y98_SLICE_X99Y98_C5 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_D1 = 1'b1;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_D2 = 1'b1;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_D3 = 1'b1;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_D4 = 1'b1;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_D5 = 1'b1;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_D6 = CLBLM_L_X60Y104_SLICE_X90Y104_AQ;
  assign CLBLM_R_X65Y98_SLICE_X99Y98_D1 = 1'b1;
  assign CLBLM_R_X65Y98_SLICE_X99Y98_D6 = CLBLM_L_X64Y100_SLICE_X96Y100_D_XOR;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_DX = 1'b0;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X65Y98_SLICE_X99Y98_D2 = CLBLM_R_X63Y95_SLICE_X95Y95_B5Q;
  assign CLBLM_R_X65Y98_SLICE_X99Y98_D3 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_R_X65Y98_SLICE_X99Y98_D4 = 1'b1;
  assign CLBLM_R_X65Y98_SLICE_X99Y98_D5 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X65Y98_SLICE_X98Y98_A1 = CLBLM_R_X65Y98_SLICE_X99Y98_CO6;
  assign CLBLM_R_X65Y98_SLICE_X98Y98_A2 = CLBLM_R_X65Y97_SLICE_X98Y97_BO6;
  assign CLBLM_R_X65Y98_SLICE_X98Y98_A3 = CLBLM_R_X65Y97_SLICE_X98Y97_AO6;
  assign CLBLM_R_X65Y98_SLICE_X98Y98_A4 = CLBLM_R_X65Y97_SLICE_X98Y97_AO5;
  assign CLBLM_R_X65Y98_SLICE_X98Y98_A5 = CLBLM_L_X64Y102_SLICE_X96Y102_C_XOR;
  assign CLBLM_R_X65Y98_SLICE_X98Y98_A6 = CLBLM_R_X65Y102_SLICE_X99Y102_BO6;
  assign CLBLM_R_X65Y98_SLICE_X98Y98_B1 = 1'b1;
  assign CLBLM_R_X65Y98_SLICE_X98Y98_B2 = CLBLM_R_X65Y97_SLICE_X98Y97_AO5;
  assign CLBLM_R_X65Y98_SLICE_X98Y98_B3 = 1'b1;
  assign CLBLM_R_X65Y98_SLICE_X98Y98_B4 = 1'b1;
  assign CLBLM_R_X65Y98_SLICE_X98Y98_B5 = CLBLM_L_X64Y98_SLICE_X96Y98_BO6;
  assign CLBLM_R_X65Y98_SLICE_X98Y98_B6 = CLBLM_R_X65Y100_SLICE_X99Y100_CQ;
  assign CLBLM_R_X65Y98_SLICE_X98Y98_C1 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_R_X65Y98_SLICE_X98Y98_C2 = CLBLM_R_X65Y101_SLICE_X99Y101_BO6;
  assign CLBLM_R_X65Y98_SLICE_X98Y98_C3 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X65Y98_SLICE_X98Y98_C4 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_R_X65Y98_SLICE_X98Y98_C5 = CLBLM_L_X64Y100_SLICE_X97Y100_AQ;
  assign CLBLM_R_X65Y98_SLICE_X98Y98_C6 = CLBLM_L_X64Y100_SLICE_X96Y100_D_XOR;
  assign CLBLM_R_X65Y98_SLICE_X98Y98_CE = CLBLM_L_X60Y98_SLICE_X91Y98_BQ;
  assign CLBLM_R_X65Y98_SLICE_X98Y98_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X65Y98_SLICE_X98Y98_D1 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_R_X65Y98_SLICE_X98Y98_D2 = 1'b1;
  assign CLBLM_R_X65Y98_SLICE_X98Y98_D3 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_R_X65Y98_SLICE_X98Y98_D4 = CLBLM_R_X65Y102_SLICE_X98Y102_A_XOR;
  assign CLBLM_R_X65Y98_SLICE_X98Y98_D5 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X65Y98_SLICE_X98Y98_D6 = CLBLM_L_X60Y98_SLICE_X90Y98_AQ;
  assign CLBLM_R_X65Y98_SLICE_X98Y98_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_D1 = CLBLM_R_X49Y111_SLICE_X74Y111_CQ;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_D1 = CLBLM_R_X49Y109_SLICE_X74Y109_BQ;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_T1 = 1'b1;
  assign CLBLM_L_X60Y109_SLICE_X91Y109_A1 = CLBLM_L_X62Y97_SLICE_X92Y97_BO6;
  assign CLBLM_L_X60Y109_SLICE_X91Y109_A2 = CLBLM_L_X60Y107_SLICE_X91Y107_A_XOR;
  assign CLBLM_L_X60Y109_SLICE_X91Y109_A3 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X60Y109_SLICE_X91Y109_A4 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X60Y109_SLICE_X91Y109_A5 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X60Y109_SLICE_X91Y109_A6 = CLBLM_L_X60Y104_SLICE_X91Y104_A_XOR;
  assign CLBLM_L_X60Y109_SLICE_X91Y109_B1 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X60Y109_SLICE_X91Y109_B2 = CLBLM_L_X62Y100_SLICE_X93Y100_BO6;
  assign CLBLM_L_X60Y109_SLICE_X91Y109_B3 = CLBLM_L_X60Y107_SLICE_X91Y107_C_XOR;
  assign CLBLM_L_X60Y109_SLICE_X91Y109_B4 = CLBLM_L_X60Y104_SLICE_X91Y104_C_XOR;
  assign CLBLM_L_X60Y109_SLICE_X91Y109_B5 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X60Y109_SLICE_X91Y109_B6 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X60Y109_SLICE_X91Y109_C1 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_L_X60Y109_SLICE_X91Y109_C2 = CLBLM_L_X60Y107_SLICE_X91Y107_C_XOR;
  assign CLBLM_L_X60Y109_SLICE_X91Y109_C3 = CLBLM_L_X60Y109_SLICE_X91Y109_BQ;
  assign CLBLM_L_X60Y109_SLICE_X91Y109_C4 = CLBLM_R_X59Y103_SLICE_X89Y103_CQ;
  assign CLBLM_L_X60Y109_SLICE_X91Y109_C5 = CLBLM_L_X60Y109_SLICE_X91Y109_DO6;
  assign CLBLM_L_X60Y109_SLICE_X91Y109_C6 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X60Y109_SLICE_X91Y109_CE = CLBLM_L_X62Y102_SLICE_X92Y102_CO6;
  assign CLBLM_L_X60Y109_SLICE_X91Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X60Y109_SLICE_X91Y109_D1 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X60Y109_SLICE_X91Y109_D2 = 1'b1;
  assign CLBLM_L_X60Y109_SLICE_X91Y109_D3 = 1'b1;
  assign CLBLM_L_X60Y109_SLICE_X91Y109_D4 = CLBLM_R_X59Y110_SLICE_X89Y110_AQ;
  assign CLBLM_L_X60Y109_SLICE_X91Y109_D5 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_L_X60Y109_SLICE_X91Y109_D6 = CLBLM_L_X60Y107_SLICE_X90Y107_D_XOR;
  assign CLBLM_L_X60Y109_SLICE_X91Y109_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X60Y109_SLICE_X90Y109_A1 = 1'b1;
  assign CLBLM_L_X60Y109_SLICE_X90Y109_A2 = 1'b1;
  assign CLBLM_L_X60Y109_SLICE_X90Y109_A3 = 1'b1;
  assign CLBLM_L_X60Y109_SLICE_X90Y109_A4 = 1'b1;
  assign CLBLM_L_X60Y109_SLICE_X90Y109_A5 = 1'b1;
  assign CLBLM_L_X60Y109_SLICE_X90Y109_A6 = CLBLM_R_X59Y112_SLICE_X89Y112_AQ;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_A1 = CLBLM_L_X64Y100_SLICE_X96Y100_A_XOR;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_A2 = CLBLM_R_X65Y99_SLICE_X99Y99_CO6;
  assign CLBLM_L_X60Y109_SLICE_X90Y109_AX = 1'b0;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_A3 = CLBLM_R_X65Y100_SLICE_X99Y100_DO6;
  assign CLBLM_L_X60Y109_SLICE_X90Y109_B1 = 1'b1;
  assign CLBLM_L_X60Y109_SLICE_X90Y109_B2 = 1'b1;
  assign CLBLM_L_X60Y109_SLICE_X90Y109_B3 = 1'b1;
  assign CLBLM_L_X60Y109_SLICE_X90Y109_B4 = 1'b1;
  assign CLBLM_L_X60Y109_SLICE_X90Y109_B5 = 1'b1;
  assign CLBLM_L_X60Y109_SLICE_X90Y109_B6 = CLBLM_R_X59Y112_SLICE_X89Y112_BQ;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_A6 = CLBLM_R_X65Y97_SLICE_X98Y97_AO5;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_B1 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_L_X60Y109_SLICE_X90Y109_BX = 1'b0;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_B2 = CLBLM_R_X63Y95_SLICE_X95Y95_BQ;
  assign CLBLM_L_X60Y109_SLICE_X90Y109_C1 = 1'b1;
  assign CLBLM_L_X60Y109_SLICE_X90Y109_C2 = 1'b1;
  assign CLBLM_L_X60Y109_SLICE_X90Y109_C3 = 1'b1;
  assign CLBLM_L_X60Y109_SLICE_X90Y109_C4 = 1'b1;
  assign CLBLM_L_X60Y109_SLICE_X90Y109_C5 = 1'b1;
  assign CLBLM_L_X60Y109_SLICE_X90Y109_C6 = CLBLM_R_X59Y106_SLICE_X89Y106_BQ;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_C2 = 1'b1;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_B5 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_C5 = CLBLM_L_X60Y98_SLICE_X90Y98_AQ;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_C6 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_L_X60Y109_SLICE_X90Y109_CIN = CLBLM_L_X60Y108_SLICE_X90Y108_COUT;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_C3 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_C4 = CLBLM_R_X65Y100_SLICE_X98Y100_B_XOR;
  assign CLBLM_L_X60Y109_SLICE_X90Y109_CX = 1'b0;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_CE = CLBLM_L_X60Y98_SLICE_X91Y98_BQ;
  assign CLBLM_L_X60Y109_SLICE_X90Y109_D1 = 1'b1;
  assign CLBLM_L_X60Y109_SLICE_X90Y109_D2 = 1'b1;
  assign CLBLM_L_X60Y109_SLICE_X90Y109_D3 = 1'b1;
  assign CLBLM_L_X60Y109_SLICE_X90Y109_D4 = 1'b1;
  assign CLBLM_L_X60Y109_SLICE_X90Y109_D5 = 1'b1;
  assign CLBLM_L_X60Y109_SLICE_X90Y109_D6 = CLBLM_R_X59Y111_SLICE_X89Y111_CQ;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_D1 = CLBLM_R_X65Y100_SLICE_X98Y100_D_XOR;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_D2 = 1'b1;
  assign CLBLM_L_X60Y109_SLICE_X90Y109_DX = 1'b0;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_D3 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_D4 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_D5 = CLBLM_L_X60Y98_SLICE_X90Y98_AQ;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_D6 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_A1 = CLBLM_R_X65Y99_SLICE_X98Y99_DO6;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_A2 = CLBLM_R_X65Y97_SLICE_X98Y97_AO5;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_A3 = CLBLM_R_X65Y96_SLICE_X98Y96_AO6;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_A4 = CLBLM_L_X64Y100_SLICE_X96Y100_B_XOR;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_A5 = CLBLM_R_X65Y97_SLICE_X98Y97_AO6;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_A6 = CLBLM_R_X65Y99_SLICE_X98Y99_CO6;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_B1 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_B2 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_B3 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_B4 = CLBLM_L_X56Y97_SLICE_X85Y97_AQ;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_B5 = 1'b1;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_B6 = CLBLM_R_X63Y97_SLICE_X94Y97_DQ;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_C1 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_C2 = CLBLM_L_X60Y98_SLICE_X90Y98_AQ;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_C3 = 1'b1;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_C4 = CLBLM_R_X65Y100_SLICE_X98Y100_C_XOR;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_C5 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_C6 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_CE = CLBLM_L_X60Y98_SLICE_X91Y98_BQ;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_D1 = CLBLM_L_X64Y100_SLICE_X97Y100_C_XOR;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_D2 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_D3 = CLBLM_L_X62Y101_SLICE_X93Y101_AQ;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_D4 = 1'b1;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_D5 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_D6 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_R_X65Y99_SLICE_X98Y99_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X60Y111_SLICE_X90Y111_B4 = CLBLM_R_X59Y106_SLICE_X89Y106_AO6;
  assign CLBLM_L_X60Y111_SLICE_X90Y111_B5 = CLBLM_L_X60Y108_SLICE_X91Y108_AQ;
  assign CLBLM_L_X60Y111_SLICE_X90Y111_B6 = CLBLM_R_X59Y110_SLICE_X88Y110_A_XOR;
  assign CLBLM_L_X60Y111_SLICE_X90Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X60Y110_SLICE_X91Y110_A1 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X60Y110_SLICE_X91Y110_A2 = CLBLM_R_X49Y104_SLICE_X75Y104_DQ;
  assign CLBLM_L_X60Y110_SLICE_X91Y110_A3 = CLBLM_R_X59Y103_SLICE_X89Y103_DQ;
  assign CLBLM_L_X60Y110_SLICE_X91Y110_A4 = CLBLM_L_X60Y110_SLICE_X91Y110_BO6;
  assign CLBLM_L_X60Y110_SLICE_X91Y110_A5 = 1'b1;
  assign CLBLM_L_X60Y110_SLICE_X91Y110_A6 = CLBLM_L_X60Y108_SLICE_X91Y108_CO6;
  assign CLBLM_L_X60Y110_SLICE_X91Y110_B1 = CLBLM_L_X60Y108_SLICE_X91Y108_DO6;
  assign CLBLM_L_X60Y110_SLICE_X91Y110_B2 = CLBLM_R_X59Y106_SLICE_X89Y106_AO6;
  assign CLBLM_L_X60Y110_SLICE_X91Y110_B3 = CLBLM_L_X62Y106_SLICE_X92Y106_AO5;
  assign CLBLM_L_X60Y110_SLICE_X91Y110_B4 = CLBLM_L_X60Y108_SLICE_X90Y108_D_XOR;
  assign CLBLM_L_X60Y110_SLICE_X91Y110_B5 = CLBLL_R_X57Y103_SLICE_X87Y103_AQ;
  assign CLBLM_L_X60Y110_SLICE_X91Y110_B6 = CLBLM_R_X59Y109_SLICE_X88Y109_A_XOR;
  assign CLBLM_L_X60Y110_SLICE_X91Y110_C1 = CLBLM_L_X60Y107_SLICE_X90Y107_C_XOR;
  assign CLBLM_L_X60Y110_SLICE_X91Y110_C2 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_L_X60Y110_SLICE_X91Y110_C3 = 1'b1;
  assign CLBLM_L_X60Y110_SLICE_X91Y110_C4 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X60Y110_SLICE_X91Y110_C5 = 1'b1;
  assign CLBLM_L_X60Y110_SLICE_X91Y110_C6 = CLBLM_R_X59Y111_SLICE_X89Y111_BQ;
  assign CLBLM_L_X60Y110_SLICE_X91Y110_CE = CLBLM_R_X59Y99_SLICE_X89Y99_CO6;
  assign CLBLM_L_X60Y110_SLICE_X91Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X60Y110_SLICE_X91Y110_D1 = CLBLM_L_X60Y106_SLICE_X90Y106_C_XOR;
  assign CLBLM_L_X60Y110_SLICE_X91Y110_D2 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X60Y110_SLICE_X91Y110_D3 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_L_X60Y110_SLICE_X91Y110_D4 = CLBLM_R_X59Y112_SLICE_X89Y112_BQ;
  assign CLBLM_L_X60Y110_SLICE_X91Y110_D5 = 1'b1;
  assign CLBLM_L_X60Y110_SLICE_X91Y110_D6 = 1'b1;
  assign CLBLM_L_X60Y110_SLICE_X91Y110_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X60Y110_SLICE_X90Y110_A1 = 1'b1;
  assign CLBLM_L_X60Y110_SLICE_X90Y110_A2 = 1'b1;
  assign CLBLM_L_X60Y110_SLICE_X90Y110_A3 = 1'b1;
  assign CLBLM_L_X60Y110_SLICE_X90Y110_A4 = 1'b1;
  assign CLBLM_L_X60Y110_SLICE_X90Y110_A5 = 1'b1;
  assign CLBLM_L_X60Y110_SLICE_X90Y110_A6 = CLBLM_R_X59Y111_SLICE_X89Y111_AQ;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_A1 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_A2 = CLBLM_R_X65Y99_SLICE_X99Y99_AQ;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_A3 = 1'b1;
  assign CLBLM_L_X60Y110_SLICE_X90Y110_AX = 1'b0;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_A5 = CLBLL_R_X57Y103_SLICE_X86Y103_AQ;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_A6 = CLBLL_R_X57Y103_SLICE_X86Y103_A5Q;
  assign CLBLM_L_X60Y110_SLICE_X90Y110_B1 = 1'b1;
  assign CLBLM_L_X60Y110_SLICE_X90Y110_B2 = 1'b1;
  assign CLBLM_L_X60Y110_SLICE_X90Y110_B3 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_B1 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_B2 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_B3 = CLBLM_R_X65Y98_SLICE_X99Y98_AQ;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_B4 = CLBLM_L_X62Y105_SLICE_X93Y105_BQ;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_B5 = CLBLL_R_X57Y103_SLICE_X86Y103_AQ;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_B6 = CLBLL_R_X57Y103_SLICE_X86Y103_A5Q;
  assign CLBLM_L_X60Y110_SLICE_X90Y110_B4 = 1'b1;
  assign CLBLM_L_X60Y110_SLICE_X90Y110_C2 = 1'b1;
  assign CLBLM_L_X60Y110_SLICE_X90Y110_C3 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_C1 = CLBLL_R_X57Y103_SLICE_X86Y103_AQ;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_C2 = CLBLL_R_X57Y103_SLICE_X86Y103_A5Q;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_C3 = CLBLM_R_X63Y104_SLICE_X94Y104_AQ;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_C4 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_C5 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_C6 = CLBLM_R_X65Y98_SLICE_X98Y98_BQ;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_CE = CLBLM_L_X62Y105_SLICE_X93Y105_DO6;
  assign CLBLM_L_X60Y110_SLICE_X90Y110_C4 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X60Y110_SLICE_X90Y110_C5 = 1'b1;
  assign CLBLM_L_X60Y110_SLICE_X90Y110_C6 = CLBLM_R_X59Y110_SLICE_X89Y110_AQ;
  assign CLBLM_L_X60Y110_SLICE_X90Y110_CIN = CLBLM_L_X60Y109_SLICE_X90Y109_COUT;
  assign CLBLM_L_X60Y110_SLICE_X90Y110_CX = 1'b0;
  assign CLBLM_L_X60Y110_SLICE_X90Y110_D1 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_D1 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_D2 = CLBLM_L_X64Y100_SLICE_X97Y100_B_XOR;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_D3 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_D4 = CLBLM_L_X62Y100_SLICE_X92Y100_BQ;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_D5 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_D6 = 1'b1;
  assign CLBLM_L_X60Y110_SLICE_X90Y110_D2 = 1'b1;
  assign CLBLM_L_X60Y110_SLICE_X90Y110_D3 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X60Y110_SLICE_X90Y110_D5 = 1'b1;
  assign CLBLM_L_X60Y110_SLICE_X90Y110_D6 = 1'b1;
  assign CLBLM_L_X60Y110_SLICE_X90Y110_DX = 1'b0;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_A1 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_A2 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_A3 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_A4 = CLBLM_L_X62Y100_SLICE_X92Y100_AQ;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_A5 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_A6 = CLBLM_R_X65Y100_SLICE_X99Y100_CQ;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_AX = CLBLM_R_X65Y100_SLICE_X99Y100_CQ;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_B1 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_B2 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_B3 = CLBLM_L_X62Y100_SLICE_X92Y100_BQ;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_B4 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_B5 = CLBLM_R_X65Y100_SLICE_X99Y100_AQ;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_B6 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_BX = CLBLM_R_X65Y100_SLICE_X99Y100_AQ;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_C1 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_C2 = CLBLM_L_X62Y101_SLICE_X93Y101_AQ;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_C3 = CLBLM_R_X65Y106_SLICE_X98Y106_CQ;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_C4 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_C5 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_C6 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_CX = CLBLM_R_X65Y106_SLICE_X98Y106_CQ;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_D1 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_D2 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_D3 = CLBLM_L_X64Y106_SLICE_X97Y106_DQ;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_D4 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_D5 = 1'b1;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_D6 = CLBLM_L_X62Y100_SLICE_X92Y100_CQ;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_DX = CLBLM_L_X64Y106_SLICE_X97Y106_DQ;
  assign CLBLM_R_X65Y96_SLICE_X99Y96_B2 = 1'b1;
  assign CLBLM_R_X65Y96_SLICE_X99Y96_B3 = 1'b1;
  assign CLBLM_R_X65Y96_SLICE_X99Y96_B4 = 1'b1;
  assign CLBLM_R_X65Y96_SLICE_X99Y96_B6 = 1'b1;
  assign CLBLM_R_X65Y96_SLICE_X99Y96_C5 = 1'b1;
  assign CLBLM_R_X65Y96_SLICE_X99Y96_C6 = 1'b1;
  assign CLBLL_L_X54Y97_SLICE_X83Y97_B4 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLL_L_X54Y97_SLICE_X83Y97_B5 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign CLBLM_L_X60Y111_SLICE_X91Y111_A1 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLM_L_X60Y111_SLICE_X91Y111_A2 = CLBLM_L_X60Y109_SLICE_X91Y109_CO6;
  assign CLBLM_L_X60Y111_SLICE_X91Y111_A3 = 1'b1;
  assign CLBLM_L_X60Y111_SLICE_X91Y111_A4 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X60Y111_SLICE_X91Y111_A5 = CLBLM_R_X59Y103_SLICE_X89Y103_DQ;
  assign CLBLM_L_X60Y111_SLICE_X91Y111_A6 = CLBLM_R_X59Y111_SLICE_X89Y111_DO6;
  assign CLBLM_L_X60Y111_SLICE_X91Y111_B1 = CLBLM_R_X49Y108_SLICE_X75Y108_DQ;
  assign CLBLM_L_X60Y111_SLICE_X91Y111_B2 = CLBLM_L_X60Y111_SLICE_X90Y111_BO6;
  assign CLBLM_L_X60Y111_SLICE_X91Y111_B3 = 1'b1;
  assign CLBLM_L_X60Y111_SLICE_X91Y111_B4 = CLBLM_R_X59Y103_SLICE_X89Y103_DQ;
  assign CLBLM_L_X60Y111_SLICE_X91Y111_B5 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X60Y111_SLICE_X91Y111_B6 = CLBLM_L_X60Y111_SLICE_X91Y111_CO6;
  assign CLBLM_L_X60Y111_SLICE_X91Y111_C1 = CLBLM_R_X59Y103_SLICE_X89Y103_CQ;
  assign CLBLM_L_X60Y111_SLICE_X91Y111_C2 = CLBLM_L_X60Y106_SLICE_X91Y106_D_XOR;
  assign CLBLM_L_X60Y111_SLICE_X91Y111_C3 = CLBLM_L_X60Y101_SLICE_X90Y101_AQ;
  assign CLBLM_L_X60Y111_SLICE_X91Y111_C4 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_L_X60Y111_SLICE_X91Y111_C5 = CLBLM_L_X60Y111_SLICE_X91Y111_DO6;
  assign CLBLM_L_X60Y111_SLICE_X91Y111_C6 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X60Y111_SLICE_X91Y111_CE = CLBLM_R_X59Y99_SLICE_X89Y99_CO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_D1 = CLBLM_R_X49Y111_SLICE_X74Y111_AQ;
  assign CLBLM_L_X60Y111_SLICE_X91Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X60Y111_SLICE_X91Y111_D1 = CLBLM_R_X59Y111_SLICE_X89Y111_CQ;
  assign CLBLM_L_X60Y111_SLICE_X91Y111_D2 = CLBLM_L_X60Y107_SLICE_X90Y107_A_XOR;
  assign CLBLM_L_X60Y111_SLICE_X91Y111_D3 = 1'b1;
  assign CLBLM_L_X60Y111_SLICE_X91Y111_D4 = 1'b1;
  assign CLBLM_L_X60Y111_SLICE_X91Y111_D5 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_L_X60Y111_SLICE_X91Y111_D6 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_T1 = 1'b1;
  assign CLBLM_L_X60Y111_SLICE_X91Y111_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X60Y111_SLICE_X90Y111_A1 = CLBLM_R_X59Y111_SLICE_X88Y111_CO6;
  assign CLBLM_L_X60Y111_SLICE_X90Y111_A2 = CLBLM_R_X59Y103_SLICE_X89Y103_DQ;
  assign CLBLM_L_X60Y111_SLICE_X90Y111_A3 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X60Y111_SLICE_X90Y111_A4 = CLBLM_R_X49Y107_SLICE_X75Y107_DQ;
  assign CLBLM_L_X60Y111_SLICE_X90Y111_A5 = 1'b1;
  assign CLBLM_L_X60Y111_SLICE_X90Y111_A6 = CLBLM_L_X60Y111_SLICE_X90Y111_CO6;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_A1 = CLBLM_R_X65Y101_SLICE_X99Y101_DO6;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_A2 = CLBLM_R_X65Y97_SLICE_X99Y97_CO6;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_A3 = CLBLM_L_X64Y101_SLICE_X96Y101_A_XOR;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_A4 = CLBLM_R_X65Y97_SLICE_X98Y97_AO5;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_A5 = CLBLM_R_X65Y97_SLICE_X98Y97_AO6;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_A6 = CLBLM_R_X65Y101_SLICE_X99Y101_CO6;
  assign CLBLM_L_X60Y111_SLICE_X90Y111_B1 = CLBLM_L_X62Y106_SLICE_X92Y106_AO5;
  assign CLBLM_L_X60Y111_SLICE_X90Y111_B2 = CLBLM_L_X60Y109_SLICE_X90Y109_D_XOR;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_B1 = CLBLM_L_X60Y98_SLICE_X90Y98_AQ;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_B2 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_B3 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_B4 = CLBLM_R_X65Y101_SLICE_X98Y101_A_XOR;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_B5 = CLBLM_L_X64Y101_SLICE_X97Y101_A_XOR;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_B6 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_L_X60Y111_SLICE_X90Y111_B3 = CLBLM_R_X59Y111_SLICE_X88Y111_BO6;
  assign CLBLM_L_X60Y111_SLICE_X90Y111_C1 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_C1 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_C2 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_C3 = CLBLM_R_X65Y101_SLICE_X98Y101_B_XOR;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_C4 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_C5 = CLBLM_L_X60Y98_SLICE_X90Y98_AQ;
  assign CLBLM_L_X60Y111_SLICE_X90Y111_C2 = CLBLM_R_X59Y103_SLICE_X89Y103_CQ;
  assign CLBLM_L_X60Y111_SLICE_X90Y111_C3 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X60Y111_SLICE_X90Y111_C4 = CLBLM_L_X60Y109_SLICE_X91Y109_AQ;
  assign CLBLM_L_X60Y111_SLICE_X90Y111_C5 = CLBLM_L_X60Y111_SLICE_X90Y111_DO6;
  assign CLBLM_L_X60Y111_SLICE_X90Y111_C6 = CLBLM_L_X60Y107_SLICE_X91Y107_A_XOR;
  assign CLBLM_L_X60Y111_SLICE_X90Y111_CE = CLBLM_R_X59Y99_SLICE_X89Y99_CO6;
  assign CLBLM_L_X60Y111_SLICE_X90Y111_D1 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_L_X60Y111_SLICE_X90Y111_D2 = 1'b1;
  assign CLBLM_L_X60Y111_SLICE_X90Y111_D3 = CLBLM_L_X60Y107_SLICE_X90Y107_B_XOR;
  assign CLBLM_L_X60Y111_SLICE_X90Y111_D4 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X60Y111_SLICE_X90Y111_D5 = 1'b1;
  assign CLBLM_L_X60Y111_SLICE_X90Y111_D6 = CLBLM_R_X59Y111_SLICE_X89Y111_AQ;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_D5 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_D6 = CLBLM_L_X64Y100_SLICE_X97Y100_BQ;
  assign CLBLM_L_X60Y111_SLICE_X90Y111_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_D2 = CLBLM_L_X64Y101_SLICE_X97Y101_B_XOR;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_D3 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_D4 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_A1 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_A2 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_A3 = CLBLM_L_X64Y100_SLICE_X97Y100_AQ;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_A4 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_A5 = CLBLM_R_X65Y100_SLICE_X99Y100_BQ;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_A6 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_AX = CLBLM_R_X65Y100_SLICE_X99Y100_BQ;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_B1 = CLBLM_R_X65Y106_SLICE_X98Y106_DQ;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_B2 = CLBLM_L_X64Y100_SLICE_X97Y100_BQ;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_B3 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_B4 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_B5 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_B6 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_BX = CLBLM_R_X65Y106_SLICE_X98Y106_DQ;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_C1 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_C2 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_C3 = CLBLM_L_X62Y101_SLICE_X93Y101_BQ;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_C4 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_C5 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_C6 = CLBLM_R_X63Y103_SLICE_X95Y103_BQ;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_CIN = CLBLM_R_X65Y100_SLICE_X98Y100_COUT;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_CX = CLBLM_R_X63Y103_SLICE_X95Y103_BQ;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_D1 = CLBLM_R_X63Y101_SLICE_X95Y101_AQ;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_D2 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_D3 = CLBLM_L_X62Y101_SLICE_X93Y101_CQ;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_D4 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_D5 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_D6 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_DX = CLBLM_L_X62Y101_SLICE_X93Y101_CQ;
  assign CLBLM_L_X60Y112_SLICE_X91Y112_A1 = 1'b1;
  assign CLBLM_L_X60Y112_SLICE_X91Y112_A2 = 1'b1;
  assign CLBLM_L_X60Y112_SLICE_X91Y112_A3 = 1'b1;
  assign CLBLM_L_X60Y112_SLICE_X91Y112_A4 = 1'b1;
  assign CLBLM_L_X60Y112_SLICE_X91Y112_A5 = 1'b1;
  assign CLBLM_L_X60Y112_SLICE_X91Y112_A6 = 1'b1;
  assign CLBLM_L_X60Y112_SLICE_X91Y112_B1 = 1'b1;
  assign CLBLM_L_X60Y112_SLICE_X91Y112_B2 = 1'b1;
  assign CLBLM_L_X60Y112_SLICE_X91Y112_B3 = 1'b1;
  assign CLBLM_L_X60Y112_SLICE_X91Y112_B4 = 1'b1;
  assign CLBLM_L_X60Y112_SLICE_X91Y112_B5 = 1'b1;
  assign CLBLM_L_X60Y112_SLICE_X91Y112_B6 = 1'b1;
  assign CLBLM_L_X60Y112_SLICE_X91Y112_C1 = 1'b1;
  assign CLBLM_L_X60Y112_SLICE_X91Y112_C2 = 1'b1;
  assign CLBLM_L_X60Y112_SLICE_X91Y112_C3 = 1'b1;
  assign CLBLM_L_X60Y112_SLICE_X91Y112_C4 = 1'b1;
  assign CLBLM_L_X60Y112_SLICE_X91Y112_C5 = 1'b1;
  assign CLBLM_L_X60Y112_SLICE_X91Y112_C6 = 1'b1;
  assign CLBLM_L_X60Y112_SLICE_X91Y112_D1 = 1'b1;
  assign CLBLM_L_X60Y112_SLICE_X91Y112_D2 = 1'b1;
  assign CLBLM_L_X60Y112_SLICE_X91Y112_D3 = 1'b1;
  assign CLBLM_L_X60Y112_SLICE_X91Y112_D4 = 1'b1;
  assign CLBLM_L_X60Y112_SLICE_X91Y112_D5 = 1'b1;
  assign CLBLM_L_X60Y112_SLICE_X91Y112_D6 = 1'b1;
  assign CLBLM_L_X60Y112_SLICE_X90Y112_A1 = CLBLM_R_X59Y99_SLICE_X89Y99_AQ;
  assign CLBLM_L_X60Y112_SLICE_X90Y112_A2 = CLBLM_R_X59Y108_SLICE_X88Y108_AQ;
  assign CLBLM_L_X60Y112_SLICE_X90Y112_A3 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_L_X60Y112_SLICE_X90Y112_A4 = CLBLM_R_X59Y103_SLICE_X89Y103_DQ;
  assign CLBLM_L_X60Y112_SLICE_X90Y112_A5 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X60Y112_SLICE_X90Y112_A6 = CLBLM_R_X59Y103_SLICE_X89Y103_CQ;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_A1 = CLBLM_L_X64Y99_SLICE_X97Y99_DO6;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_A2 = CLBLM_L_X64Y102_SLICE_X96Y102_A_XOR;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_A3 = CLBLM_R_X65Y97_SLICE_X98Y97_AO6;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_A4 = CLBLM_R_X65Y97_SLICE_X98Y97_AO5;
  assign CLBLM_L_X60Y112_SLICE_X90Y112_B1 = CLBLM_R_X59Y99_SLICE_X89Y99_A5Q;
  assign CLBLM_L_X60Y112_SLICE_X90Y112_B2 = CLBLM_R_X59Y103_SLICE_X89Y103_DQ;
  assign CLBLM_L_X60Y112_SLICE_X90Y112_B3 = CLBLM_L_X60Y107_SLICE_X90Y107_AQ;
  assign CLBLM_L_X60Y112_SLICE_X90Y112_B4 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_L_X60Y112_SLICE_X90Y112_B5 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X60Y112_SLICE_X90Y112_B6 = CLBLM_R_X59Y103_SLICE_X89Y103_CQ;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_A5 = CLBLM_R_X63Y102_SLICE_X95Y102_AO6;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_A6 = CLBLM_R_X65Y102_SLICE_X99Y102_CO6;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_B1 = CLBLM_L_X60Y98_SLICE_X90Y98_AQ;
  assign CLBLM_L_X60Y112_SLICE_X90Y112_C1 = 1'b1;
  assign CLBLM_L_X60Y112_SLICE_X90Y112_C2 = 1'b1;
  assign CLBLM_L_X60Y112_SLICE_X90Y112_C3 = 1'b1;
  assign CLBLM_L_X60Y112_SLICE_X90Y112_C4 = 1'b1;
  assign CLBLM_L_X60Y112_SLICE_X90Y112_C5 = 1'b1;
  assign CLBLM_L_X60Y112_SLICE_X90Y112_C6 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_B4 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_B5 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_C5 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_C6 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_CE = CLBLM_L_X60Y98_SLICE_X91Y98_BQ;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_C1 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_C3 = CLBLM_R_X65Y102_SLICE_X98Y102_B_XOR;
  assign CLBLM_L_X60Y112_SLICE_X90Y112_D1 = 1'b1;
  assign CLBLM_L_X60Y112_SLICE_X90Y112_D2 = 1'b1;
  assign CLBLM_L_X60Y112_SLICE_X90Y112_D3 = 1'b1;
  assign CLBLM_L_X60Y112_SLICE_X90Y112_D4 = 1'b1;
  assign CLBLM_L_X60Y112_SLICE_X90Y112_D5 = 1'b1;
  assign CLBLM_L_X60Y112_SLICE_X90Y112_D6 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_D1 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_D2 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_D3 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_D4 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_D5 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_D6 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_A1 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_A2 = CLBLM_R_X63Y103_SLICE_X95Y103_CQ;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_A3 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_A4 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_A5 = CLBLM_L_X62Y101_SLICE_X93Y101_CQ;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_A6 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_B1 = CLBLM_R_X65Y107_SLICE_X98Y107_DQ;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_B2 = CLBLM_R_X63Y103_SLICE_X95Y103_CQ;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_B3 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_B4 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_B5 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_B6 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_BX = CLBLM_R_X63Y103_SLICE_X95Y103_CQ;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_C1 = CLBLM_R_X65Y107_SLICE_X98Y107_AQ;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_C2 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_C3 = CLBLM_R_X65Y107_SLICE_X98Y107_DQ;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_C4 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_C5 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_C6 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_CIN = CLBLM_R_X65Y101_SLICE_X98Y101_COUT;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_CX = CLBLM_R_X65Y107_SLICE_X98Y107_DQ;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_D1 = CLBLM_R_X65Y107_SLICE_X98Y107_AQ;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_D2 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_D3 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_D4 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_D5 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_D6 = CLBLM_R_X65Y107_SLICE_X98Y107_BQ;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_DX = CLBLM_R_X65Y107_SLICE_X98Y107_AQ;
  assign CLK_HROW_BOT_R_X139Y78_BUFHCE_X0Y20_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_A1 = CLBLM_L_X64Y105_SLICE_X96Y105_CO6;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_A2 = CLBLM_R_X63Y98_SLICE_X94Y98_DO6;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_A3 = CLBLM_R_X65Y97_SLICE_X98Y97_AO6;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_A4 = CLBLM_R_X65Y97_SLICE_X98Y97_AO5;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_A5 = CLBLM_R_X65Y103_SLICE_X99Y103_CO6;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_A6 = CLBLM_L_X64Y103_SLICE_X96Y103_B_XOR;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_B1 = CLBLM_R_X65Y103_SLICE_X99Y103_DO6;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_B2 = CLBLM_L_X64Y103_SLICE_X96Y103_C_XOR;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_B3 = CLBLM_R_X65Y97_SLICE_X98Y97_AO6;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_B4 = CLBLM_R_X65Y97_SLICE_X98Y97_AO5;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_B5 = CLBLM_R_X63Y103_SLICE_X95Y103_DO6;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_B6 = CLBLM_R_X65Y97_SLICE_X99Y97_AO6;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_C1 = CLBLM_L_X60Y98_SLICE_X90Y98_AQ;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_C2 = CLBLM_R_X65Y103_SLICE_X98Y103_C_XOR;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_C3 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_C4 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_C5 = 1'b1;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_C6 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_CE = CLBLM_L_X60Y98_SLICE_X91Y98_BQ;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_D1 = CLBLM_L_X60Y98_SLICE_X90Y98_AQ;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_D2 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_D3 = CLBLM_R_X65Y103_SLICE_X98Y103_D_XOR;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_D4 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_D5 = 1'b1;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_D6 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X65Y103_SLICE_X99Y103_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_A1 = CLBLM_R_X65Y107_SLICE_X98Y107_CQ;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_A2 = 1'b1;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_A3 = 1'b1;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_A4 = CLBLM_R_X65Y107_SLICE_X98Y107_BQ;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_A5 = 1'b1;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_A6 = 1'b1;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_AX = CLBLM_R_X65Y107_SLICE_X98Y107_BQ;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_B1 = CLBLM_R_X65Y107_SLICE_X98Y107_CQ;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_B2 = 1'b1;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_B3 = CLBLM_R_X65Y106_SLICE_X98Y106_AQ;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_B4 = 1'b1;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_B5 = 1'b1;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_B6 = 1'b1;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_BX = CLBLM_R_X65Y107_SLICE_X98Y107_CQ;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_C1 = 1'b1;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_C2 = 1'b1;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_C3 = CLBLM_R_X65Y106_SLICE_X98Y106_AQ;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_C4 = 1'b1;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_C5 = CLBLM_L_X64Y106_SLICE_X97Y106_AQ;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_C6 = 1'b1;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_CIN = CLBLM_R_X65Y102_SLICE_X98Y102_COUT;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_CX = CLBLM_R_X65Y106_SLICE_X98Y106_AQ;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_D1 = CLBLM_R_X63Y103_SLICE_X95Y103_AQ;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_D2 = 1'b1;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_D3 = CLBLM_L_X64Y106_SLICE_X97Y106_AQ;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_D4 = 1'b1;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_D5 = 1'b1;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_D6 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_D1 = CLBLM_R_X49Y109_SLICE_X74Y109_AQ;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_DX = CLBLM_L_X64Y106_SLICE_X97Y106_AQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_T1 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_D1 = CLBLM_R_X49Y111_SLICE_X74Y111_BQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_T1 = 1'b1;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_A1 = CLBLM_L_X64Y105_SLICE_X97Y105_CO6;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_A2 = CLBLM_R_X65Y104_SLICE_X99Y104_CO6;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_A3 = CLBLM_L_X64Y102_SLICE_X96Y102_D_XOR;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_A4 = CLBLM_L_X62Y97_SLICE_X93Y97_DO6;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_A5 = CLBLM_R_X65Y97_SLICE_X98Y97_AO6;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_A6 = CLBLM_R_X65Y97_SLICE_X98Y97_AO5;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_B1 = CLBLM_R_X65Y104_SLICE_X99Y104_DO6;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_B2 = CLBLM_R_X65Y97_SLICE_X98Y97_DO6;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_B3 = CLBLM_R_X65Y97_SLICE_X98Y97_AO6;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_B4 = CLBLM_L_X64Y103_SLICE_X96Y103_D_XOR;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_B5 = CLBLM_R_X63Y104_SLICE_X95Y104_AO6;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_B6 = CLBLM_R_X65Y97_SLICE_X98Y97_AO5;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_C1 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_C2 = 1'b1;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_C3 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_C4 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_C5 = CLBLM_L_X60Y98_SLICE_X90Y98_AQ;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_C6 = CLBLM_R_X65Y103_SLICE_X98Y103_A_XOR;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_CE = CLBLM_L_X60Y98_SLICE_X91Y98_BQ;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_D1 = 1'b1;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_D2 = CLBLM_R_X65Y104_SLICE_X98Y104_A_XOR;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_D3 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_D4 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_D5 = CLBLM_L_X60Y98_SLICE_X90Y98_AQ;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_D6 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_R_X65Y104_SLICE_X99Y104_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_A1 = 1'b1;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_A2 = 1'b1;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_A3 = CLBLM_R_X63Y103_SLICE_X95Y103_AQ;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_A4 = CLBLM_R_X65Y106_SLICE_X98Y106_BQ;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_A5 = 1'b1;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_A6 = 1'b1;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_AX = CLBLM_R_X63Y103_SLICE_X95Y103_AQ;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_B1 = 1'b1;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_B2 = 1'b1;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_B3 = 1'b1;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_B4 = CLBLM_R_X65Y106_SLICE_X98Y106_BQ;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_B5 = 1'b1;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_B6 = CLBLM_L_X64Y106_SLICE_X97Y106_BQ;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_BX = CLBLM_R_X65Y106_SLICE_X98Y106_BQ;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_C1 = 1'b1;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_C2 = 1'b1;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_C3 = CLBLM_L_X64Y106_SLICE_X97Y106_BQ;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_C4 = 1'b1;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_C5 = CLBLM_L_X64Y106_SLICE_X97Y106_CQ;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_C6 = 1'b1;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_CIN = CLBLM_R_X65Y103_SLICE_X98Y103_COUT;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_CX = 1'b0;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_D1 = 1'b1;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_D2 = 1'b1;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_D3 = 1'b1;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_D4 = 1'b1;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_D5 = 1'b1;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_D6 = 1'b1;
  assign CLBLM_R_X65Y104_SLICE_X98Y104_DX = 1'b0;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_A1 = CLBLM_R_X65Y105_SLICE_X99Y105_DO6;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_A2 = CLBLM_R_X65Y97_SLICE_X98Y97_AO5;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_A3 = CLBLM_R_X65Y97_SLICE_X98Y97_AO6;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_A4 = CLBLM_R_X65Y97_SLICE_X99Y97_BO6;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_A5 = CLBLM_L_X64Y104_SLICE_X96Y104_B_XOR;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_A6 = CLBLM_L_X64Y105_SLICE_X97Y105_DO6;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_B1 = CLBLM_R_X65Y103_SLICE_X98Y103_B_XOR;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_B2 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_B3 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_B4 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_B5 = CLBLM_L_X60Y98_SLICE_X90Y98_AQ;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_B6 = 1'b1;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_C1 = CLBLM_L_X60Y98_SLICE_X90Y98_AQ;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_C2 = CLBLM_R_X65Y104_SLICE_X98Y104_B_XOR;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_C3 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_C4 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_C5 = 1'b1;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_C6 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_CE = CLBLM_L_X60Y98_SLICE_X91Y98_BQ;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_D1 = CLBLM_L_X60Y98_SLICE_X90Y98_AQ;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_D2 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_D3 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_D4 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_D5 = 1'b1;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_D6 = CLBLM_R_X65Y104_SLICE_X98Y104_C_XOR;
  assign CLBLM_R_X65Y105_SLICE_X99Y105_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_A1 = CLBLM_R_X65Y97_SLICE_X98Y97_CO6;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_A2 = CLBLM_R_X65Y105_SLICE_X99Y105_BO6;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_A3 = CLBLM_R_X65Y97_SLICE_X98Y97_AO6;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_A4 = CLBLM_L_X64Y103_SLICE_X96Y103_A_XOR;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_A5 = CLBLM_R_X65Y97_SLICE_X98Y97_AO5;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_A6 = CLBLM_R_X65Y105_SLICE_X98Y105_CO6;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_B1 = CLBLM_R_X65Y105_SLICE_X98Y105_DO6;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_B2 = CLBLM_R_X65Y97_SLICE_X98Y97_AO5;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_B3 = CLBLM_R_X65Y99_SLICE_X98Y99_BO6;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_B4 = CLBLM_R_X65Y105_SLICE_X99Y105_CO6;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_B5 = CLBLM_R_X65Y97_SLICE_X98Y97_AO6;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_B6 = CLBLM_L_X64Y104_SLICE_X96Y104_A_XOR;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_C1 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_C2 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_C3 = CLBLM_R_X49Y106_SLICE_X75Y106_CQ;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_C4 = CLBLM_L_X64Y103_SLICE_X97Y103_B_XOR;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_C5 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_C6 = 1'b1;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_CE = CLBLM_L_X60Y98_SLICE_X91Y98_BQ;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_D1 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_D2 = 1'b1;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_D3 = CLBLM_L_X64Y104_SLICE_X97Y104_B_XOR;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_D4 = CLBLM_R_X49Y107_SLICE_X75Y107_DQ;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_D5 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_D6 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_R_X65Y105_SLICE_X98Y105_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign LIOB33_SING_X0Y149_IOB_X0Y149_O = CLBLM_R_X49Y111_SLICE_X75Y111_A5Q;
  assign CLBLM_R_X65Y97_SLICE_X99Y97_B2 = 1'b1;
  assign CLBLM_R_X65Y97_SLICE_X99Y97_B3 = CLBLM_L_X56Y97_SLICE_X85Y97_AQ;
  assign CLBLM_R_X65Y97_SLICE_X99Y97_B4 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X65Y97_SLICE_X99Y97_B6 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_R_X65Y97_SLICE_X99Y97_C5 = CLBLM_R_X63Y95_SLICE_X95Y95_C5Q;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_D1 = CLBLM_L_X50Y104_SLICE_X76Y104_AQ;
  assign CLBLM_R_X65Y97_SLICE_X99Y97_C6 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_T1 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_D1 = CLBLM_R_X49Y109_SLICE_X74Y109_CQ;
  assign CLBLL_L_X54Y98_SLICE_X83Y98_C5 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_T1 = 1'b1;
  assign CLBLL_L_X54Y98_SLICE_X83Y98_CE = CLBLM_L_X60Y98_SLICE_X91Y98_DQ;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_D1 = CLBLM_R_X65Y100_SLICE_X99Y100_CQ;
  assign CLBLM_L_X50Y104_SLICE_X77Y104_A1 = CLBLM_R_X53Y101_SLICE_X81Y101_AQ;
  assign CLBLM_L_X50Y104_SLICE_X77Y104_A2 = CLBLL_L_X54Y100_SLICE_X82Y100_BQ;
  assign CLBLM_L_X50Y104_SLICE_X77Y104_A3 = CLBLL_R_X57Y100_SLICE_X86Y100_BQ;
  assign CLBLM_L_X50Y104_SLICE_X77Y104_A4 = CLBLM_L_X56Y101_SLICE_X85Y101_DQ;
  assign CLBLM_L_X50Y104_SLICE_X77Y104_A5 = CLBLL_R_X57Y100_SLICE_X86Y100_CQ;
  assign CLBLM_L_X50Y104_SLICE_X77Y104_A6 = CLBLM_R_X53Y101_SLICE_X80Y101_BQ;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_T1 = 1'b1;
  assign CLBLM_L_X50Y104_SLICE_X77Y104_B1 = 1'b1;
  assign CLBLM_L_X50Y104_SLICE_X77Y104_B2 = 1'b1;
  assign CLBLM_L_X50Y104_SLICE_X77Y104_B3 = 1'b1;
  assign CLBLM_L_X50Y104_SLICE_X77Y104_B4 = 1'b1;
  assign CLBLM_L_X50Y104_SLICE_X77Y104_B5 = 1'b1;
  assign CLBLM_L_X50Y104_SLICE_X77Y104_B6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_D1 = 1'b0;
  assign CLBLM_L_X50Y104_SLICE_X77Y104_C1 = 1'b1;
  assign CLBLM_L_X50Y104_SLICE_X77Y104_C2 = 1'b1;
  assign CLBLM_L_X50Y104_SLICE_X77Y104_C3 = 1'b1;
  assign CLBLM_L_X50Y104_SLICE_X77Y104_C4 = 1'b1;
  assign CLBLM_L_X50Y104_SLICE_X77Y104_C5 = 1'b1;
  assign CLBLM_L_X50Y104_SLICE_X77Y104_C6 = 1'b1;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_A1 = 1'b1;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_A2 = 1'b1;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_A3 = 1'b1;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_A4 = 1'b1;
  assign CLBLM_L_X50Y104_SLICE_X77Y104_D1 = 1'b1;
  assign CLBLM_L_X50Y104_SLICE_X77Y104_D2 = 1'b1;
  assign CLBLM_L_X50Y104_SLICE_X77Y104_D3 = 1'b1;
  assign CLBLM_L_X50Y104_SLICE_X77Y104_D4 = 1'b1;
  assign CLBLM_L_X50Y104_SLICE_X77Y104_D5 = 1'b1;
  assign CLBLM_L_X50Y104_SLICE_X77Y104_D6 = 1'b1;
  assign CLBLM_L_X56Y97_SLICE_X85Y97_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_A5 = 1'b1;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_A6 = 1'b1;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_B1 = 1'b1;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_B2 = 1'b1;
  assign CLBLM_L_X50Y104_SLICE_X76Y104_A1 = CLBLM_L_X50Y107_SLICE_X76Y107_CO6;
  assign CLBLM_L_X50Y104_SLICE_X76Y104_A2 = CLBLM_R_X53Y100_SLICE_X81Y100_AQ;
  assign CLBLM_L_X50Y104_SLICE_X76Y104_A3 = CLBLM_R_X53Y101_SLICE_X81Y101_AQ;
  assign CLBLM_L_X50Y104_SLICE_X76Y104_A4 = CLBLM_L_X50Y104_SLICE_X76Y104_BO6;
  assign CLBLM_L_X50Y104_SLICE_X76Y104_A5 = 1'b1;
  assign CLBLM_L_X50Y104_SLICE_X76Y104_A6 = CLBLM_L_X50Y104_SLICE_X76Y104_CO6;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_B6 = 1'b1;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_C1 = 1'b1;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_C2 = 1'b1;
  assign CLBLM_L_X50Y104_SLICE_X76Y104_B1 = CLBLL_R_X57Y100_SLICE_X86Y100_AQ;
  assign CLBLM_L_X50Y104_SLICE_X76Y104_B2 = CLBLM_L_X50Y104_SLICE_X76Y104_DO6;
  assign CLBLM_L_X50Y104_SLICE_X76Y104_B3 = CLBLL_L_X54Y100_SLICE_X82Y100_BQ;
  assign CLBLM_L_X50Y104_SLICE_X76Y104_B4 = CLBLM_R_X53Y101_SLICE_X81Y101_AQ;
  assign CLBLM_L_X50Y104_SLICE_X76Y104_B5 = CLBLM_R_X53Y101_SLICE_X80Y101_BQ;
  assign CLBLM_L_X50Y104_SLICE_X76Y104_B6 = CLBLL_R_X57Y100_SLICE_X86Y100_DQ;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_D1 = 1'b1;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_D2 = 1'b1;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_D3 = 1'b1;
  assign CLBLM_L_X50Y104_SLICE_X76Y104_C1 = CLBLM_R_X53Y101_SLICE_X80Y101_BQ;
  assign CLBLM_L_X50Y104_SLICE_X76Y104_C2 = CLBLL_L_X54Y100_SLICE_X82Y100_BQ;
  assign CLBLM_L_X50Y104_SLICE_X76Y104_C3 = CLBLL_R_X57Y101_SLICE_X87Y101_CQ;
  assign CLBLM_L_X50Y104_SLICE_X76Y104_C4 = CLBLL_R_X57Y100_SLICE_X86Y100_DQ;
  assign CLBLM_L_X50Y104_SLICE_X76Y104_C5 = CLBLL_R_X57Y100_SLICE_X86Y100_AQ;
  assign CLBLM_L_X50Y104_SLICE_X76Y104_C6 = 1'b1;
  assign CLBLM_L_X50Y104_SLICE_X76Y104_CE = CLBLM_L_X56Y98_SLICE_X84Y98_DO6;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_D4 = 1'b1;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_A1 = 1'b1;
  assign CLBLM_L_X50Y104_SLICE_X76Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_A2 = CLBLL_R_X57Y103_SLICE_X86Y103_AQ;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_A3 = CLBLM_R_X63Y110_SLICE_X94Y110_AQ;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_A4 = CLBLL_R_X57Y103_SLICE_X86Y103_A5Q;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_A5 = CLBLM_R_X65Y105_SLICE_X98Y105_AQ;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_A6 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X50Y104_SLICE_X76Y104_D1 = CLBLL_R_X57Y100_SLICE_X86Y100_CQ;
  assign CLBLM_L_X50Y104_SLICE_X76Y104_D2 = CLBLL_R_X57Y97_SLICE_X86Y97_AQ;
  assign CLBLM_L_X50Y104_SLICE_X76Y104_D3 = 1'b1;
  assign CLBLM_L_X50Y104_SLICE_X76Y104_D4 = CLBLL_R_X57Y99_SLICE_X86Y99_BQ;
  assign CLBLM_L_X50Y104_SLICE_X76Y104_D5 = CLBLM_R_X53Y101_SLICE_X80Y101_BQ;
  assign CLBLM_L_X50Y104_SLICE_X76Y104_D6 = CLBLL_L_X54Y100_SLICE_X82Y100_BQ;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_B1 = CLBLM_L_X62Y103_SLICE_X93Y103_AQ;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_B2 = CLBLL_R_X57Y103_SLICE_X86Y103_A5Q;
  assign CLBLM_L_X50Y104_SLICE_X76Y104_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_B3 = CLBLL_R_X57Y103_SLICE_X86Y103_AQ;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_B4 = 1'b1;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_B5 = CLBLM_R_X65Y104_SLICE_X99Y104_BQ;
  assign CLBLM_L_X56Y97_SLICE_X85Y97_D6 = CLBLL_L_X54Y98_SLICE_X83Y98_AQ;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_B6 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_C1 = CLBLM_L_X64Y105_SLICE_X97Y105_AQ;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_C2 = CLBLL_R_X57Y103_SLICE_X86Y103_A5Q;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_C3 = CLBLL_R_X57Y103_SLICE_X86Y103_AQ;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_C4 = 1'b1;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_C5 = CLBLM_R_X65Y99_SLICE_X98Y99_AQ;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_C6 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_CE = CLBLM_L_X62Y105_SLICE_X93Y105_DO6;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X65Y97_SLICE_X98Y97_B5 = 1'b1;
  assign CLBLM_R_X65Y97_SLICE_X98Y97_B6 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_D1 = CLBLM_R_X65Y101_SLICE_X99Y101_AQ;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_D2 = CLBLL_R_X57Y103_SLICE_X86Y103_A5Q;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_D3 = CLBLM_L_X64Y106_SLICE_X96Y106_AQ;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_D4 = CLBLL_R_X57Y103_SLICE_X86Y103_AQ;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_D5 = 1'b1;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_D6 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X65Y106_SLICE_X98Y106_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X56Y97_SLICE_X84Y97_A1 = CLBLM_R_X49Y108_SLICE_X75Y108_DQ;
  assign CLBLM_L_X56Y97_SLICE_X84Y97_A2 = CLBLM_L_X56Y97_SLICE_X85Y97_BO5;
  assign CLBLM_R_X65Y97_SLICE_X98Y97_C1 = CLBLM_L_X56Y97_SLICE_X85Y97_AQ;
  assign CLBLM_L_X56Y97_SLICE_X84Y97_A3 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLM_R_X65Y97_SLICE_X98Y97_C2 = CLBLM_L_X64Y97_SLICE_X97Y97_BQ;
  assign CLBLM_L_X56Y97_SLICE_X84Y97_A4 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLM_R_X65Y97_SLICE_X98Y97_C6 = 1'b1;
  assign CLBLM_L_X56Y97_SLICE_X84Y97_B6 = CLBLM_R_X49Y107_SLICE_X75Y107_DQ;
  assign CLBLM_L_X56Y111_SLICE_X84Y111_B4 = 1'b1;
  assign CLBLM_R_X65Y97_SLICE_X98Y97_D6 = CLBLM_R_X63Y96_SLICE_X95Y96_BQ;
  assign CLBLM_L_X56Y97_SLICE_X84Y97_C2 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLM_L_X56Y111_SLICE_X84Y111_B5 = 1'b1;
  assign CLBLM_L_X56Y97_SLICE_X84Y97_C6 = 1'b1;
  assign CLBLM_L_X50Y105_SLICE_X77Y105_A1 = CLBLM_R_X49Y106_SLICE_X74Y106_CO6;
  assign CLBLM_L_X50Y105_SLICE_X77Y105_A2 = CLBLL_L_X52Y105_SLICE_X78Y105_BO5;
  assign CLBLM_L_X50Y105_SLICE_X77Y105_A3 = CLBLL_R_X57Y100_SLICE_X86Y100_CQ;
  assign CLBLM_L_X50Y105_SLICE_X77Y105_A4 = CLBLL_R_X57Y100_SLICE_X86Y100_DQ;
  assign CLBLM_L_X50Y105_SLICE_X77Y105_A5 = CLBLL_R_X57Y100_SLICE_X86Y100_BQ;
  assign CLBLM_L_X50Y105_SLICE_X77Y105_A6 = CLBLM_L_X50Y106_SLICE_X77Y106_AO5;
  assign CLBLM_L_X50Y105_SLICE_X77Y105_AX = CLBLM_R_X53Y100_SLICE_X81Y100_AQ;
  assign CLBLM_L_X50Y105_SLICE_X77Y105_B1 = CLBLM_R_X49Y108_SLICE_X75Y108_B_XOR;
  assign CLBLM_L_X50Y105_SLICE_X77Y105_B2 = CLBLM_L_X50Y106_SLICE_X77Y106_AO6;
  assign CLBLM_L_X50Y105_SLICE_X77Y105_B3 = CLBLM_L_X50Y104_SLICE_X77Y104_AO6;
  assign CLBLM_L_X50Y105_SLICE_X77Y105_B4 = 1'b1;
  assign CLBLM_L_X50Y105_SLICE_X77Y105_B5 = CLBLM_L_X50Y107_SLICE_X76Y107_AO6;
  assign CLBLM_L_X50Y105_SLICE_X77Y105_B6 = CLBLL_L_X54Y100_SLICE_X82Y100_BQ;
  assign CLBLM_L_X50Y105_SLICE_X77Y105_C1 = CLBLL_R_X57Y99_SLICE_X86Y99_BQ;
  assign CLBLM_L_X50Y105_SLICE_X77Y105_C2 = CLBLM_L_X50Y106_SLICE_X77Y106_AO5;
  assign CLBLM_L_X50Y105_SLICE_X77Y105_C3 = CLBLL_R_X57Y99_SLICE_X86Y99_AQ;
  assign CLBLM_L_X50Y105_SLICE_X77Y105_C4 = CLBLL_L_X52Y106_SLICE_X78Y106_AO5;
  assign CLBLM_L_X50Y105_SLICE_X77Y105_C5 = CLBLM_L_X50Y105_SLICE_X77Y105_DO6;
  assign CLBLM_L_X50Y105_SLICE_X77Y105_C6 = CLBLM_R_X49Y106_SLICE_X74Y106_CO6;
  assign CLBLM_L_X50Y105_SLICE_X77Y105_CE = CLBLM_L_X56Y98_SLICE_X84Y98_DO6;
  assign CLBLM_L_X50Y105_SLICE_X77Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X65Y107_SLICE_X99Y107_A1 = 1'b1;
  assign CLBLM_R_X65Y107_SLICE_X99Y107_A2 = 1'b1;
  assign CLBLM_R_X65Y107_SLICE_X99Y107_A3 = 1'b1;
  assign CLBLM_R_X65Y107_SLICE_X99Y107_A4 = 1'b1;
  assign CLBLM_L_X50Y105_SLICE_X77Y105_D1 = CLBLL_R_X57Y97_SLICE_X86Y97_AQ;
  assign CLBLM_L_X50Y105_SLICE_X77Y105_D2 = CLBLM_R_X53Y101_SLICE_X80Y101_BQ;
  assign CLBLM_L_X50Y105_SLICE_X77Y105_D3 = 1'b1;
  assign CLBLM_L_X50Y105_SLICE_X77Y105_D4 = CLBLL_R_X57Y101_SLICE_X87Y101_DQ;
  assign CLBLM_L_X50Y105_SLICE_X77Y105_D5 = CLBLL_L_X54Y100_SLICE_X82Y100_BQ;
  assign CLBLM_L_X50Y105_SLICE_X77Y105_D6 = CLBLL_R_X57Y100_SLICE_X86Y100_DQ;
  assign CLBLM_R_X65Y107_SLICE_X99Y107_A5 = 1'b1;
  assign CLBLM_R_X65Y107_SLICE_X99Y107_A6 = 1'b1;
  assign CLBLM_L_X50Y105_SLICE_X77Y105_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X65Y107_SLICE_X99Y107_B1 = 1'b1;
  assign CLBLM_R_X65Y107_SLICE_X99Y107_B2 = 1'b1;
  assign CLBLM_L_X50Y105_SLICE_X76Y105_A1 = CLBLM_L_X50Y105_SLICE_X76Y105_BO5;
  assign CLBLM_L_X50Y105_SLICE_X76Y105_A2 = CLBLL_L_X52Y105_SLICE_X78Y105_CO6;
  assign CLBLM_L_X50Y105_SLICE_X76Y105_A3 = CLBLM_L_X50Y111_SLICE_X76Y111_AO6;
  assign CLBLM_L_X50Y105_SLICE_X76Y105_A4 = CLBLM_L_X50Y111_SLICE_X76Y111_BO6;
  assign CLBLM_L_X50Y105_SLICE_X76Y105_A5 = CLBLM_L_X50Y105_SLICE_X76Y105_CO5;
  assign CLBLM_L_X50Y105_SLICE_X76Y105_A6 = 1'b1;
  assign CLBLM_R_X65Y107_SLICE_X99Y107_B6 = 1'b1;
  assign CLBLM_R_X65Y107_SLICE_X99Y107_C1 = 1'b1;
  assign CLBLM_R_X65Y107_SLICE_X99Y107_C2 = 1'b1;
  assign CLBLM_L_X50Y105_SLICE_X76Y105_B1 = CLBLL_R_X57Y99_SLICE_X86Y99_BQ;
  assign CLBLM_L_X50Y105_SLICE_X76Y105_B2 = CLBLM_R_X53Y100_SLICE_X81Y100_AQ;
  assign CLBLM_L_X50Y105_SLICE_X76Y105_B3 = CLBLM_L_X56Y101_SLICE_X85Y101_DQ;
  assign CLBLM_L_X50Y105_SLICE_X76Y105_B4 = CLBLL_R_X57Y97_SLICE_X86Y97_AQ;
  assign CLBLM_L_X50Y105_SLICE_X76Y105_B5 = CLBLL_L_X54Y100_SLICE_X82Y100_BQ;
  assign CLBLM_L_X50Y105_SLICE_X76Y105_B6 = 1'b1;
  assign CLBLM_R_X65Y107_SLICE_X99Y107_D1 = 1'b1;
  assign CLBLM_R_X65Y107_SLICE_X99Y107_D2 = 1'b1;
  assign CLBLM_R_X65Y107_SLICE_X99Y107_D3 = 1'b1;
  assign CLBLM_L_X50Y105_SLICE_X76Y105_C1 = CLBLM_R_X53Y100_SLICE_X81Y100_AQ;
  assign CLBLM_L_X50Y105_SLICE_X76Y105_C2 = CLBLL_R_X57Y97_SLICE_X86Y97_AQ;
  assign CLBLM_L_X50Y105_SLICE_X76Y105_C3 = CLBLL_L_X52Y105_SLICE_X78Y105_AO6;
  assign CLBLM_L_X50Y105_SLICE_X76Y105_C4 = CLBLM_R_X53Y101_SLICE_X80Y101_BQ;
  assign CLBLM_L_X50Y105_SLICE_X76Y105_C5 = CLBLM_R_X53Y101_SLICE_X81Y101_AQ;
  assign CLBLM_L_X50Y105_SLICE_X76Y105_C6 = 1'b1;
  assign CLBLM_L_X50Y105_SLICE_X76Y105_CE = CLBLM_L_X56Y98_SLICE_X84Y98_DO6;
  assign CLBLM_R_X65Y107_SLICE_X99Y107_D4 = 1'b1;
  assign CLBLM_R_X65Y107_SLICE_X98Y107_A1 = CLBLL_R_X57Y103_SLICE_X86Y103_AQ;
  assign CLBLM_L_X50Y105_SLICE_X76Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X65Y107_SLICE_X98Y107_A2 = CLBLL_R_X57Y103_SLICE_X86Y103_A5Q;
  assign CLBLM_R_X65Y107_SLICE_X98Y107_A3 = CLBLM_L_X64Y99_SLICE_X96Y99_AQ;
  assign CLBLM_R_X65Y107_SLICE_X98Y107_A4 = 1'b1;
  assign CLBLM_R_X65Y107_SLICE_X98Y107_A5 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X65Y107_SLICE_X98Y107_A6 = CLBLM_L_X64Y107_SLICE_X97Y107_AQ;
  assign CLBLM_L_X50Y105_SLICE_X76Y105_D1 = 1'b1;
  assign CLBLM_L_X50Y105_SLICE_X76Y105_D2 = 1'b1;
  assign CLBLM_L_X50Y105_SLICE_X76Y105_D3 = 1'b1;
  assign CLBLM_L_X50Y105_SLICE_X76Y105_D4 = 1'b1;
  assign CLBLM_L_X50Y105_SLICE_X76Y105_D5 = 1'b1;
  assign CLBLM_L_X50Y105_SLICE_X76Y105_D6 = 1'b1;
  assign CLBLM_R_X65Y107_SLICE_X98Y107_B1 = CLBLL_R_X57Y103_SLICE_X86Y103_AQ;
  assign CLBLM_R_X65Y107_SLICE_X98Y107_B2 = 1'b1;
  assign CLBLM_L_X50Y105_SLICE_X76Y105_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X65Y107_SLICE_X98Y107_B3 = CLBLM_L_X64Y108_SLICE_X96Y108_AQ;
  assign CLBLM_R_X65Y107_SLICE_X98Y107_B4 = CLBLL_R_X57Y103_SLICE_X86Y103_A5Q;
  assign CLBLM_R_X65Y107_SLICE_X98Y107_B5 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X65Y107_SLICE_X98Y107_B6 = CLBLM_R_X65Y98_SLICE_X98Y98_AQ;
  assign CLBLM_R_X65Y107_SLICE_X98Y107_C1 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X65Y107_SLICE_X98Y107_C2 = CLBLL_R_X57Y103_SLICE_X86Y103_AQ;
  assign CLBLM_R_X65Y107_SLICE_X98Y107_C3 = CLBLM_L_X64Y108_SLICE_X97Y108_AQ;
  assign CLBLM_R_X65Y107_SLICE_X98Y107_C4 = 1'b1;
  assign CLBLM_R_X65Y107_SLICE_X98Y107_C5 = CLBLM_R_X65Y104_SLICE_X99Y104_AQ;
  assign CLBLM_R_X65Y107_SLICE_X98Y107_C6 = CLBLL_R_X57Y103_SLICE_X86Y103_A5Q;
  assign CLBLM_R_X65Y107_SLICE_X98Y107_CE = CLBLM_L_X62Y105_SLICE_X93Y105_DO6;
  assign CLBLM_R_X65Y107_SLICE_X98Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X65Y107_SLICE_X98Y107_D1 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X65Y107_SLICE_X98Y107_D2 = CLBLL_R_X57Y103_SLICE_X86Y103_AQ;
  assign CLBLM_R_X65Y107_SLICE_X98Y107_D3 = CLBLM_R_X65Y102_SLICE_X99Y102_AQ;
  assign CLBLM_R_X65Y107_SLICE_X98Y107_D4 = CLBLM_L_X64Y107_SLICE_X96Y107_BQ;
  assign CLBLM_R_X65Y107_SLICE_X98Y107_D5 = 1'b1;
  assign CLBLM_R_X65Y107_SLICE_X98Y107_D6 = CLBLL_R_X57Y103_SLICE_X86Y103_A5Q;
  assign CLBLM_R_X65Y107_SLICE_X98Y107_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X50Y106_SLICE_X77Y106_A1 = CLBLM_R_X53Y101_SLICE_X80Y101_BQ;
  assign CLBLM_L_X50Y106_SLICE_X77Y106_A2 = CLBLM_L_X50Y108_SLICE_X76Y108_B_XOR;
  assign CLBLM_L_X50Y106_SLICE_X77Y106_A3 = CLBLM_R_X53Y101_SLICE_X81Y101_AQ;
  assign CLBLM_L_X50Y106_SLICE_X77Y106_A4 = CLBLL_L_X54Y100_SLICE_X82Y100_BQ;
  assign CLBLM_L_X50Y106_SLICE_X77Y106_A5 = CLBLM_L_X50Y108_SLICE_X77Y108_B_XOR;
  assign CLBLM_L_X50Y106_SLICE_X77Y106_A6 = 1'b1;
  assign CLBLM_L_X50Y106_SLICE_X77Y106_B1 = CLBLL_R_X57Y101_SLICE_X87Y101_CQ;
  assign CLBLM_L_X50Y106_SLICE_X77Y106_B2 = CLBLL_R_X57Y101_SLICE_X87Y101_DQ;
  assign CLBLM_L_X50Y106_SLICE_X77Y106_B3 = CLBLL_L_X54Y100_SLICE_X82Y100_BQ;
  assign CLBLM_L_X50Y106_SLICE_X77Y106_B4 = CLBLL_R_X57Y100_SLICE_X87Y100_CQ;
  assign CLBLM_L_X50Y106_SLICE_X77Y106_B5 = CLBLM_L_X56Y101_SLICE_X85Y101_DQ;
  assign CLBLM_L_X50Y106_SLICE_X77Y106_B6 = 1'b1;
  assign CLBLM_L_X50Y106_SLICE_X77Y106_C1 = CLBLM_L_X56Y101_SLICE_X85Y101_BQ;
  assign CLBLM_L_X50Y106_SLICE_X77Y106_C2 = CLBLM_R_X49Y106_SLICE_X74Y106_CO6;
  assign CLBLM_L_X50Y106_SLICE_X77Y106_C3 = CLBLM_L_X50Y106_SLICE_X76Y106_BO5;
  assign CLBLM_L_X50Y106_SLICE_X77Y106_C4 = CLBLM_L_X50Y106_SLICE_X77Y106_AO5;
  assign CLBLM_L_X50Y106_SLICE_X77Y106_C5 = CLBLM_L_X50Y106_SLICE_X77Y106_BO5;
  assign CLBLM_L_X50Y106_SLICE_X77Y106_C6 = CLBLM_L_X56Y101_SLICE_X85Y101_DQ;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_D1 = CLBLM_R_X49Y105_SLICE_X75Y105_CQ;
  assign CLBLM_L_X50Y106_SLICE_X77Y106_D1 = 1'b1;
  assign CLBLM_L_X50Y106_SLICE_X77Y106_D2 = 1'b1;
  assign CLBLM_L_X50Y106_SLICE_X77Y106_D3 = 1'b1;
  assign CLBLM_L_X50Y106_SLICE_X77Y106_D4 = 1'b1;
  assign CLBLM_L_X50Y106_SLICE_X77Y106_D5 = 1'b1;
  assign CLBLM_L_X50Y106_SLICE_X77Y106_D6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_T1 = 1'b1;
  assign CLBLM_L_X50Y106_SLICE_X76Y106_A1 = CLBLM_L_X50Y106_SLICE_X76Y106_DO6;
  assign CLBLM_L_X50Y106_SLICE_X76Y106_A2 = CLBLM_R_X49Y107_SLICE_X74Y107_BO6;
  assign CLBLM_L_X50Y106_SLICE_X76Y106_A3 = 1'b1;
  assign CLBLM_L_X50Y106_SLICE_X76Y106_A4 = CLBLL_L_X52Y106_SLICE_X79Y106_AO5;
  assign CLBLM_L_X50Y106_SLICE_X76Y106_A5 = CLBLM_R_X53Y100_SLICE_X81Y100_AQ;
  assign CLBLM_L_X50Y106_SLICE_X76Y106_A6 = CLBLM_R_X53Y101_SLICE_X81Y101_AQ;
  assign CLBLM_R_X59Y96_SLICE_X89Y96_A1 = CLBLM_L_X60Y98_SLICE_X90Y98_DO6;
  assign CLBLM_R_X59Y96_SLICE_X89Y96_A2 = CLBLM_L_X50Y107_SLICE_X76Y107_BQ;
  assign CLBLM_R_X59Y96_SLICE_X89Y96_A3 = CLBLM_L_X60Y96_SLICE_X90Y96_AQ;
  assign CLBLM_R_X59Y96_SLICE_X89Y96_A4 = CLBLM_L_X50Y107_SLICE_X77Y107_AQ;
  assign CLBLM_L_X50Y106_SLICE_X76Y106_B1 = CLBLL_R_X57Y101_SLICE_X87Y101_CQ;
  assign CLBLM_L_X50Y106_SLICE_X76Y106_B2 = CLBLL_R_X57Y100_SLICE_X86Y100_CQ;
  assign CLBLM_L_X50Y106_SLICE_X76Y106_B3 = CLBLL_R_X57Y100_SLICE_X86Y100_DQ;
  assign CLBLM_L_X50Y106_SLICE_X76Y106_B4 = CLBLL_R_X57Y100_SLICE_X87Y100_CQ;
  assign CLBLM_L_X50Y106_SLICE_X76Y106_B5 = CLBLM_L_X56Y101_SLICE_X85Y101_CQ;
  assign CLBLM_L_X50Y106_SLICE_X76Y106_B6 = 1'b1;
  assign CLBLM_R_X59Y96_SLICE_X89Y96_B2 = CLBLM_L_X56Y98_SLICE_X85Y98_CQ;
  assign CLBLM_R_X59Y96_SLICE_X89Y96_B3 = CLBLM_L_X56Y98_SLICE_X85Y98_BQ;
  assign CLBLM_R_X59Y96_SLICE_X89Y96_B4 = CLBLM_R_X59Y96_SLICE_X88Y96_BQ;
  assign CLBLM_R_X59Y96_SLICE_X89Y96_B5 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X59Y96_SLICE_X89Y96_B1 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X50Y106_SLICE_X76Y106_C1 = 1'b1;
  assign CLBLM_L_X50Y106_SLICE_X76Y106_C2 = CLBLM_L_X50Y106_SLICE_X77Y106_CO6;
  assign CLBLM_L_X50Y106_SLICE_X76Y106_C3 = CLBLM_R_X49Y108_SLICE_X74Y108_DO6;
  assign CLBLM_L_X50Y106_SLICE_X76Y106_C4 = CLBLM_R_X53Y101_SLICE_X81Y101_AQ;
  assign CLBLM_L_X50Y106_SLICE_X76Y106_C5 = CLBLM_R_X53Y100_SLICE_X81Y100_AQ;
  assign CLBLM_R_X59Y96_SLICE_X89Y96_C4 = 1'b1;
  assign CLBLM_R_X59Y96_SLICE_X89Y96_C5 = 1'b1;
  assign CLBLM_R_X59Y96_SLICE_X89Y96_C6 = 1'b1;
  assign CLBLM_R_X59Y96_SLICE_X89Y96_CE = CLBLM_R_X59Y98_SLICE_X89Y98_DO6;
  assign CLBLM_L_X50Y106_SLICE_X76Y106_C6 = CLBLL_L_X52Y107_SLICE_X78Y107_AO5;
  assign CLBLM_R_X59Y96_SLICE_X89Y96_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X50Y106_SLICE_X76Y106_CE = CLBLM_L_X56Y98_SLICE_X84Y98_DO6;
  assign CLBLM_L_X50Y106_SLICE_X76Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X50Y106_SLICE_X76Y106_D1 = CLBLM_L_X50Y106_SLICE_X77Y106_BO6;
  assign CLBLM_L_X50Y106_SLICE_X76Y106_D2 = CLBLM_L_X50Y106_SLICE_X77Y106_AO5;
  assign CLBLM_L_X50Y106_SLICE_X76Y106_D3 = CLBLL_R_X57Y101_SLICE_X87Y101_AQ;
  assign CLBLM_L_X50Y106_SLICE_X76Y106_D4 = CLBLL_R_X57Y101_SLICE_X87Y101_CQ;
  assign CLBLM_L_X50Y106_SLICE_X76Y106_D5 = CLBLM_R_X49Y106_SLICE_X74Y106_CO6;
  assign CLBLM_L_X50Y106_SLICE_X76Y106_D6 = CLBLM_L_X50Y106_SLICE_X76Y106_BO6;
  assign CLBLM_R_X59Y96_SLICE_X89Y96_D1 = 1'b1;
  assign CLBLM_R_X59Y96_SLICE_X89Y96_D2 = 1'b1;
  assign CLBLM_L_X50Y106_SLICE_X76Y106_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X59Y96_SLICE_X89Y96_D3 = 1'b1;
  assign CLBLM_R_X59Y96_SLICE_X89Y96_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X59Y96_SLICE_X89Y96_D4 = 1'b1;
  assign CLBLM_R_X59Y96_SLICE_X89Y96_D5 = 1'b1;
  assign CLBLM_R_X59Y96_SLICE_X89Y96_D6 = 1'b1;
  assign CLBLM_R_X59Y96_SLICE_X88Y96_A1 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X59Y96_SLICE_X88Y96_A2 = CLBLL_R_X57Y98_SLICE_X86Y98_CO6;
  assign CLBLM_R_X59Y96_SLICE_X88Y96_A3 = CLBLM_R_X59Y96_SLICE_X88Y96_AQ;
  assign CLBLM_R_X59Y96_SLICE_X88Y96_A4 = CLBLM_L_X50Y106_SLICE_X76Y106_AQ;
  assign CLBLM_R_X59Y96_SLICE_X88Y96_A5 = CLBLM_L_X60Y99_SLICE_X91Y99_DO6;
  assign CLBLM_R_X59Y96_SLICE_X88Y96_A6 = CLBLM_R_X59Y96_SLICE_X88Y96_CO6;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_D1 = CLBLM_R_X65Y107_SLICE_X98Y107_CQ;
  assign CLBLM_R_X59Y96_SLICE_X88Y96_B1 = CLBLM_L_X60Y99_SLICE_X91Y99_DO6;
  assign CLBLM_R_X59Y96_SLICE_X88Y96_B2 = CLBLM_R_X59Y96_SLICE_X88Y96_BQ;
  assign CLBLM_R_X59Y96_SLICE_X88Y96_B3 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X59Y96_SLICE_X88Y96_B4 = CLBLM_R_X59Y96_SLICE_X88Y96_DO6;
  assign CLBLM_R_X59Y96_SLICE_X88Y96_B5 = CLBLL_R_X57Y98_SLICE_X86Y98_BO6;
  assign CLBLM_R_X59Y96_SLICE_X88Y96_B6 = CLBLM_R_X49Y106_SLICE_X74Y106_AQ;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_T1 = 1'b1;
  assign CLBLM_R_X59Y96_SLICE_X88Y96_C1 = CLBLM_L_X50Y107_SLICE_X77Y107_AQ;
  assign CLBLM_R_X59Y96_SLICE_X88Y96_C2 = CLBLM_R_X59Y96_SLICE_X88Y96_AQ;
  assign CLBLM_R_X59Y96_SLICE_X88Y96_C3 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X59Y96_SLICE_X88Y96_C4 = CLBLL_R_X57Y97_SLICE_X86Y97_CO6;
  assign CLBLM_R_X59Y96_SLICE_X88Y96_C5 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X59Y96_SLICE_X88Y96_C6 = CLBLM_R_X59Y97_SLICE_X89Y97_B5Q;
  assign CLBLM_R_X59Y96_SLICE_X88Y96_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_D1 = CLBLM_R_X65Y107_SLICE_X98Y107_BQ;
  assign CLBLM_R_X59Y96_SLICE_X88Y96_D1 = CLBLM_L_X50Y107_SLICE_X77Y107_AQ;
  assign CLBLM_R_X59Y96_SLICE_X88Y96_D2 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X59Y96_SLICE_X88Y96_D3 = CLBLL_R_X57Y99_SLICE_X86Y99_AQ;
  assign CLBLM_R_X59Y96_SLICE_X88Y96_D4 = CLBLM_R_X59Y96_SLICE_X89Y96_BO6;
  assign CLBLM_R_X59Y96_SLICE_X88Y96_D5 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X59Y96_SLICE_X88Y96_D6 = CLBLL_R_X57Y99_SLICE_X86Y99_BQ;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_T1 = 1'b1;
  assign CLBLM_R_X59Y96_SLICE_X88Y96_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X50Y107_SLICE_X77Y107_A1 = 1'b1;
  assign CLBLM_L_X50Y107_SLICE_X77Y107_A2 = CLBLM_L_X50Y105_SLICE_X77Y105_CO6;
  assign CLBLM_L_X50Y107_SLICE_X77Y107_A3 = CLBLM_R_X53Y100_SLICE_X81Y100_AQ;
  assign CLBLM_L_X50Y107_SLICE_X77Y107_A4 = CLBLM_L_X50Y107_SLICE_X77Y107_BO6;
  assign CLBLM_L_X50Y107_SLICE_X77Y107_A5 = CLBLM_L_X50Y107_SLICE_X76Y107_DO6;
  assign CLBLM_L_X50Y107_SLICE_X77Y107_A6 = CLBLM_R_X53Y101_SLICE_X81Y101_AQ;
  assign CLBLM_L_X50Y107_SLICE_X77Y107_B1 = 1'b1;
  assign CLBLM_L_X50Y107_SLICE_X77Y107_B2 = CLBLL_R_X57Y99_SLICE_X86Y99_AQ;
  assign CLBLM_L_X50Y107_SLICE_X77Y107_B3 = CLBLL_L_X54Y100_SLICE_X82Y100_BQ;
  assign CLBLM_L_X50Y107_SLICE_X77Y107_B4 = CLBLL_R_X57Y100_SLICE_X87Y100_CQ;
  assign CLBLM_L_X50Y107_SLICE_X77Y107_B5 = CLBLM_R_X53Y101_SLICE_X80Y101_BQ;
  assign CLBLM_L_X50Y107_SLICE_X77Y107_B6 = CLBLL_R_X57Y99_SLICE_X86Y99_BQ;
  assign CLBLM_L_X50Y107_SLICE_X77Y107_C1 = 1'b1;
  assign CLBLM_L_X50Y107_SLICE_X77Y107_C2 = 1'b1;
  assign CLBLM_L_X50Y107_SLICE_X77Y107_C3 = 1'b1;
  assign CLBLM_L_X50Y107_SLICE_X77Y107_C4 = 1'b1;
  assign CLBLM_L_X50Y107_SLICE_X77Y107_C5 = 1'b1;
  assign CLBLM_L_X50Y107_SLICE_X77Y107_C6 = 1'b1;
  assign CLBLM_L_X50Y107_SLICE_X77Y107_CE = CLBLM_L_X56Y98_SLICE_X84Y98_DO6;
  assign CLBLM_L_X50Y107_SLICE_X77Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X50Y107_SLICE_X77Y107_D1 = 1'b1;
  assign CLBLM_L_X50Y107_SLICE_X77Y107_D2 = 1'b1;
  assign CLBLM_L_X50Y107_SLICE_X77Y107_D3 = 1'b1;
  assign CLBLM_L_X50Y107_SLICE_X77Y107_D4 = 1'b1;
  assign CLBLM_L_X50Y107_SLICE_X77Y107_D5 = 1'b1;
  assign CLBLM_L_X50Y107_SLICE_X77Y107_D6 = 1'b1;
  assign CLBLM_L_X50Y107_SLICE_X77Y107_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X50Y107_SLICE_X76Y107_A1 = CLBLL_R_X57Y97_SLICE_X86Y97_AQ;
  assign CLBLM_L_X50Y107_SLICE_X76Y107_A2 = CLBLM_L_X50Y109_SLICE_X77Y109_D_XOR;
  assign CLBLM_L_X50Y107_SLICE_X76Y107_A3 = CLBLM_R_X49Y108_SLICE_X75Y108_A_XOR;
  assign CLBLM_L_X50Y107_SLICE_X76Y107_A4 = CLBLM_L_X50Y109_SLICE_X76Y109_D_XOR;
  assign CLBLM_L_X50Y107_SLICE_X76Y107_A5 = CLBLM_R_X53Y101_SLICE_X80Y101_BQ;
  assign CLBLM_L_X50Y107_SLICE_X76Y107_A6 = 1'b1;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_A1 = 1'b1;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_A2 = 1'b1;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_A3 = 1'b1;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_A4 = 1'b1;
  assign CLBLM_L_X50Y107_SLICE_X76Y107_B1 = 1'b1;
  assign CLBLM_L_X50Y107_SLICE_X76Y107_B2 = CLBLM_R_X53Y101_SLICE_X81Y101_AQ;
  assign CLBLM_L_X50Y107_SLICE_X76Y107_B3 = CLBLM_L_X50Y111_SLICE_X76Y111_CO6;
  assign CLBLM_L_X50Y107_SLICE_X76Y107_B4 = CLBLL_L_X52Y107_SLICE_X78Y107_BO5;
  assign CLBLM_L_X50Y107_SLICE_X76Y107_B5 = CLBLM_R_X53Y100_SLICE_X81Y100_AQ;
  assign CLBLM_L_X50Y107_SLICE_X76Y107_B6 = CLBLM_R_X49Y106_SLICE_X75Y106_CO6;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_B2 = 1'b1;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_B3 = 1'b1;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_B4 = 1'b1;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_A6 = CLBLM_R_X59Y98_SLICE_X88Y98_DQ;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_AX = CLBLM_R_X59Y96_SLICE_X88Y96_BQ;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_B1 = 1'b1;
  assign CLBLM_L_X50Y107_SLICE_X76Y107_C1 = CLBLL_L_X54Y100_SLICE_X82Y100_BQ;
  assign CLBLM_L_X50Y107_SLICE_X76Y107_C2 = CLBLM_L_X50Y108_SLICE_X76Y108_A_XOR;
  assign CLBLM_L_X50Y107_SLICE_X76Y107_C3 = CLBLL_R_X57Y97_SLICE_X86Y97_AQ;
  assign CLBLM_L_X50Y107_SLICE_X76Y107_C4 = CLBLM_R_X49Y108_SLICE_X75Y108_A_XOR;
  assign CLBLM_L_X50Y107_SLICE_X76Y107_C5 = CLBLM_L_X50Y108_SLICE_X77Y108_A_XOR;
  assign CLBLM_L_X50Y107_SLICE_X76Y107_C6 = CLBLM_R_X53Y101_SLICE_X80Y101_BQ;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_C5 = 1'b1;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_C6 = CLBLM_R_X59Y97_SLICE_X88Y97_AQ;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_CE = CLBLL_R_X57Y97_SLICE_X87Y97_AO6;
  assign CLBLM_L_X50Y107_SLICE_X76Y107_CE = CLBLM_L_X56Y98_SLICE_X84Y98_DO6;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X50Y107_SLICE_X76Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_C2 = 1'b1;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_C3 = 1'b1;
  assign CLBLM_L_X50Y107_SLICE_X76Y107_D1 = CLBLM_R_X49Y109_SLICE_X75Y109_C_XOR;
  assign CLBLM_L_X50Y107_SLICE_X76Y107_D2 = CLBLM_R_X49Y109_SLICE_X75Y109_D_XOR;
  assign CLBLM_L_X50Y107_SLICE_X76Y107_D3 = CLBLL_L_X54Y100_SLICE_X82Y100_BQ;
  assign CLBLM_L_X50Y107_SLICE_X76Y107_D4 = CLBLM_L_X50Y107_SLICE_X76Y107_AO5;
  assign CLBLM_L_X50Y107_SLICE_X76Y107_D5 = CLBLM_R_X49Y109_SLICE_X75Y109_B_XOR;
  assign CLBLM_L_X50Y107_SLICE_X76Y107_D6 = CLBLM_R_X49Y107_SLICE_X74Y107_DO6;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_CX = CLBLM_R_X59Y98_SLICE_X89Y98_BQ;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_D1 = 1'b1;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_D2 = 1'b1;
  assign CLBLM_L_X50Y107_SLICE_X76Y107_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_D3 = 1'b1;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_D4 = 1'b1;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_D5 = 1'b1;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_D6 = CLBLM_R_X59Y97_SLICE_X88Y97_BQ;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_DX = CLBLM_R_X59Y98_SLICE_X89Y98_B5Q;
  assign CLBLM_R_X59Y97_SLICE_X88Y97_A1 = CLBLM_L_X60Y99_SLICE_X91Y99_DO6;
  assign CLBLM_R_X59Y97_SLICE_X88Y97_A2 = CLBLM_R_X59Y97_SLICE_X88Y97_AQ;
  assign CLBLM_R_X59Y97_SLICE_X88Y97_A3 = CLBLL_R_X57Y98_SLICE_X86Y98_BO6;
  assign CLBLM_R_X59Y97_SLICE_X88Y97_A4 = CLBLM_L_X50Y105_SLICE_X77Y105_AQ;
  assign CLBLM_R_X59Y97_SLICE_X88Y97_A5 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X59Y97_SLICE_X88Y97_A6 = CLBLM_R_X59Y97_SLICE_X88Y97_CO6;
  assign CLBLM_R_X59Y97_SLICE_X88Y97_B1 = CLBLM_R_X59Y97_SLICE_X88Y97_DO6;
  assign CLBLM_R_X59Y97_SLICE_X88Y97_B2 = CLBLM_R_X59Y97_SLICE_X88Y97_BQ;
  assign CLBLM_R_X59Y97_SLICE_X88Y97_B3 = CLBLM_R_X49Y105_SLICE_X75Y105_CQ;
  assign CLBLM_R_X59Y97_SLICE_X88Y97_B4 = CLBLM_L_X60Y99_SLICE_X91Y99_DO6;
  assign CLBLM_R_X59Y97_SLICE_X88Y97_B5 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X59Y97_SLICE_X88Y97_B6 = CLBLL_R_X57Y98_SLICE_X86Y98_DO6;
  assign CLBLM_R_X59Y97_SLICE_X88Y97_C1 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X59Y97_SLICE_X88Y97_C2 = CLBLL_R_X57Y97_SLICE_X86Y97_CO6;
  assign CLBLM_R_X59Y97_SLICE_X88Y97_C3 = CLBLM_R_X59Y97_SLICE_X88Y97_AQ;
  assign CLBLM_R_X59Y97_SLICE_X88Y97_C4 = CLBLM_R_X59Y97_SLICE_X89Y97_CQ;
  assign CLBLM_R_X59Y97_SLICE_X88Y97_C5 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X59Y97_SLICE_X88Y97_C6 = CLBLM_L_X50Y106_SLICE_X76Y106_AQ;
  assign CLBLM_R_X59Y97_SLICE_X88Y97_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X59Y97_SLICE_X88Y97_D1 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X59Y97_SLICE_X88Y97_D2 = CLBLL_R_X57Y97_SLICE_X86Y97_CO6;
  assign CLBLM_R_X59Y97_SLICE_X88Y97_D3 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X59Y97_SLICE_X88Y97_D4 = CLBLM_R_X59Y97_SLICE_X88Y97_BQ;
  assign CLBLM_R_X59Y97_SLICE_X88Y97_D5 = CLBLM_R_X59Y97_SLICE_X89Y97_DQ;
  assign CLBLM_R_X59Y97_SLICE_X88Y97_D6 = CLBLM_L_X60Y97_SLICE_X90Y97_BO6;
  assign CLBLM_R_X59Y97_SLICE_X88Y97_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_A5 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_A6 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_C2 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_C3 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_C4 = 1'b1;
  assign CLBLM_L_X50Y108_SLICE_X77Y108_A1 = 1'b1;
  assign CLBLM_L_X50Y108_SLICE_X77Y108_A2 = 1'b1;
  assign CLBLM_L_X50Y108_SLICE_X77Y108_A3 = CLBLL_R_X57Y97_SLICE_X86Y97_AQ;
  assign CLBLM_L_X50Y108_SLICE_X77Y108_A4 = CLBLL_R_X57Y100_SLICE_X86Y100_AQ;
  assign CLBLM_L_X50Y108_SLICE_X77Y108_A5 = CLBLL_R_X57Y100_SLICE_X86Y100_DQ;
  assign CLBLM_L_X50Y108_SLICE_X77Y108_A6 = 1'b1;
  assign CLBLM_L_X50Y108_SLICE_X77Y108_AX = 1'b1;
  assign CLBLM_L_X50Y108_SLICE_X77Y108_B1 = CLBLL_R_X57Y97_SLICE_X86Y97_AQ;
  assign CLBLM_L_X50Y108_SLICE_X77Y108_B2 = CLBLL_R_X57Y100_SLICE_X86Y100_AQ;
  assign CLBLM_L_X50Y108_SLICE_X77Y108_B3 = CLBLL_R_X57Y100_SLICE_X86Y100_BQ;
  assign CLBLM_L_X50Y108_SLICE_X77Y108_B4 = CLBLL_R_X57Y100_SLICE_X86Y100_CQ;
  assign CLBLM_L_X50Y108_SLICE_X77Y108_B5 = CLBLL_R_X57Y100_SLICE_X86Y100_DQ;
  assign CLBLM_L_X50Y108_SLICE_X77Y108_B6 = 1'b1;
  assign CLBLM_L_X50Y108_SLICE_X77Y108_C1 = CLBLM_L_X56Y101_SLICE_X85Y101_AQ;
  assign CLBLM_L_X50Y108_SLICE_X77Y108_C2 = CLBLL_R_X57Y100_SLICE_X86Y100_CQ;
  assign CLBLM_L_X50Y108_SLICE_X77Y108_C3 = CLBLM_L_X56Y101_SLICE_X85Y101_CQ;
  assign CLBLM_L_X50Y108_SLICE_X77Y108_C4 = 1'b1;
  assign CLBLM_L_X50Y108_SLICE_X77Y108_C5 = CLBLL_R_X57Y100_SLICE_X86Y100_BQ;
  assign CLBLM_L_X50Y108_SLICE_X77Y108_C6 = 1'b1;
  assign CLBLM_L_X50Y108_SLICE_X77Y108_D1 = CLBLM_L_X56Y101_SLICE_X85Y101_AQ;
  assign CLBLM_L_X50Y108_SLICE_X77Y108_D2 = 1'b1;
  assign CLBLM_L_X50Y108_SLICE_X77Y108_D3 = CLBLL_R_X57Y100_SLICE_X87Y100_AQ;
  assign CLBLM_L_X50Y108_SLICE_X77Y108_D4 = CLBLM_L_X56Y101_SLICE_X85Y101_CQ;
  assign CLBLM_L_X50Y108_SLICE_X77Y108_D5 = CLBLL_R_X57Y100_SLICE_X87Y100_CQ;
  assign CLBLM_L_X50Y108_SLICE_X77Y108_D6 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_D4 = 1'b1;
  assign CLBLM_L_X50Y108_SLICE_X76Y108_A1 = 1'b1;
  assign CLBLM_L_X50Y108_SLICE_X76Y108_A2 = 1'b1;
  assign CLBLM_L_X50Y108_SLICE_X76Y108_A3 = CLBLL_R_X57Y100_SLICE_X86Y100_DQ;
  assign CLBLM_L_X50Y108_SLICE_X76Y108_A4 = CLBLL_R_X57Y100_SLICE_X86Y100_AQ;
  assign CLBLM_L_X50Y108_SLICE_X76Y108_A5 = 1'b1;
  assign CLBLM_L_X50Y108_SLICE_X76Y108_A6 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_D5 = 1'b1;
  assign CLBLM_R_X59Y98_SLICE_X89Y98_A1 = CLBLM_L_X60Y98_SLICE_X90Y98_DO6;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_D6 = 1'b1;
  assign CLBLM_L_X50Y108_SLICE_X76Y108_AX = CLBLL_R_X57Y100_SLICE_X86Y100_DQ;
  assign CLBLM_R_X59Y98_SLICE_X89Y98_A2 = CLBLM_L_X50Y104_SLICE_X76Y104_AQ;
  assign CLBLM_R_X59Y98_SLICE_X89Y98_A6 = 1'b1;
  assign CLBLM_L_X50Y108_SLICE_X76Y108_B1 = 1'b1;
  assign CLBLM_L_X50Y108_SLICE_X76Y108_B2 = CLBLL_R_X57Y100_SLICE_X86Y100_CQ;
  assign CLBLM_L_X50Y108_SLICE_X76Y108_B3 = 1'b1;
  assign CLBLM_L_X50Y108_SLICE_X76Y108_B4 = 1'b1;
  assign CLBLM_R_X59Y98_SLICE_X89Y98_B1 = CLBLM_L_X60Y98_SLICE_X90Y98_DO6;
  assign CLBLM_R_X59Y98_SLICE_X89Y98_B2 = CLBLM_R_X49Y105_SLICE_X75Y105_CQ;
  assign CLBLM_R_X59Y98_SLICE_X89Y98_B3 = CLBLM_R_X59Y97_SLICE_X89Y97_D5Q;
  assign CLBLM_R_X59Y98_SLICE_X89Y98_B4 = CLBLM_R_X59Y97_SLICE_X89Y97_C5Q;
  assign CLBLM_L_X50Y108_SLICE_X76Y108_B5 = CLBLL_R_X57Y100_SLICE_X86Y100_BQ;
  assign CLBLM_L_X50Y108_SLICE_X76Y108_B6 = 1'b1;
  assign CLBLM_L_X50Y108_SLICE_X76Y108_BX = CLBLL_R_X57Y100_SLICE_X86Y100_CQ;
  assign CLBLM_L_X50Y108_SLICE_X76Y108_C1 = CLBLM_L_X56Y101_SLICE_X85Y101_AQ;
  assign CLBLM_L_X50Y108_SLICE_X76Y108_C2 = 1'b1;
  assign CLBLM_L_X50Y108_SLICE_X76Y108_C3 = CLBLM_L_X56Y101_SLICE_X85Y101_CQ;
  assign CLBLM_L_X50Y108_SLICE_X76Y108_C4 = 1'b1;
  assign CLBLM_L_X50Y108_SLICE_X76Y108_C5 = 1'b1;
  assign CLBLM_L_X50Y108_SLICE_X76Y108_C6 = 1'b1;
  assign CLBLM_R_X59Y98_SLICE_X89Y98_C5 = CLBLM_L_X50Y106_SLICE_X76Y106_AQ;
  assign CLBLM_R_X59Y98_SLICE_X89Y98_C6 = 1'b1;
  assign CLBLM_R_X59Y98_SLICE_X89Y98_CE = CLBLM_R_X59Y98_SLICE_X89Y98_DO6;
  assign CLBLM_R_X59Y98_SLICE_X89Y98_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X59Y98_SLICE_X89Y98_C1 = CLBLM_L_X50Y106_SLICE_X76Y106_CQ;
  assign CLBLM_R_X59Y98_SLICE_X89Y98_C2 = CLBLL_R_X57Y98_SLICE_X87Y98_CQ;
  assign CLBLM_R_X59Y98_SLICE_X89Y98_C3 = CLBLL_R_X57Y98_SLICE_X87Y98_DQ;
  assign CLBLM_L_X50Y108_SLICE_X76Y108_CX = CLBLM_L_X56Y101_SLICE_X85Y101_CQ;
  assign CLBLM_L_X50Y108_SLICE_X76Y108_D1 = CLBLL_R_X57Y100_SLICE_X87Y100_AQ;
  assign CLBLM_L_X50Y108_SLICE_X76Y108_D2 = 1'b1;
  assign CLBLM_L_X50Y108_SLICE_X76Y108_D3 = CLBLL_R_X57Y100_SLICE_X87Y100_CQ;
  assign CLBLM_L_X50Y108_SLICE_X76Y108_D4 = 1'b1;
  assign CLBLM_L_X50Y108_SLICE_X76Y108_D5 = 1'b1;
  assign CLBLM_L_X50Y108_SLICE_X76Y108_D6 = 1'b1;
  assign CLBLM_R_X59Y98_SLICE_X89Y98_D5 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X59Y98_SLICE_X89Y98_D1 = CLBLM_L_X56Y98_SLICE_X85Y98_BQ;
  assign CLBLM_R_X59Y98_SLICE_X89Y98_D6 = CLBLM_L_X56Y98_SLICE_X85Y98_CQ;
  assign CLBLM_L_X50Y108_SLICE_X76Y108_DX = CLBLL_R_X57Y100_SLICE_X87Y100_CQ;
  assign CLBLM_R_X59Y98_SLICE_X89Y98_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X59Y98_SLICE_X89Y98_D3 = CLBLM_L_X60Y98_SLICE_X91Y98_DQ;
  assign CLBLM_R_X59Y98_SLICE_X89Y98_D4 = CLBLM_L_X60Y98_SLICE_X90Y98_DO6;
  assign CLBLM_R_X59Y98_SLICE_X88Y98_A1 = CLBLM_L_X50Y105_SLICE_X77Y105_AQ;
  assign CLBLM_R_X59Y98_SLICE_X88Y98_A2 = CLBLM_L_X62Y100_SLICE_X92Y100_BQ;
  assign CLBLM_R_X59Y98_SLICE_X88Y98_A3 = CLBLM_L_X60Y99_SLICE_X91Y99_AO5;
  assign CLBLM_R_X59Y98_SLICE_X88Y98_A4 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X59Y98_SLICE_X88Y98_A5 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X59Y98_SLICE_X88Y98_A6 = CLBLM_R_X59Y97_SLICE_X89Y97_BQ;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_A4 = 1'b1;
  assign CLBLM_R_X59Y98_SLICE_X88Y98_B1 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X59Y98_SLICE_X88Y98_B2 = CLBLM_L_X62Y101_SLICE_X93Y101_AQ;
  assign CLBLM_R_X59Y98_SLICE_X88Y98_B3 = CLBLM_L_X60Y99_SLICE_X91Y99_AO5;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_A5 = 1'b1;
  assign CLBLM_R_X59Y98_SLICE_X88Y98_B4 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X59Y98_SLICE_X88Y98_B5 = CLBLM_R_X59Y100_SLICE_X88Y100_AQ;
  assign CLBLM_R_X59Y98_SLICE_X88Y98_B6 = CLBLM_R_X49Y105_SLICE_X75Y105_CQ;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_A6 = 1'b1;
  assign CLBLM_R_X59Y98_SLICE_X88Y98_C1 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X59Y98_SLICE_X88Y98_C2 = CLBLM_R_X59Y100_SLICE_X88Y100_CQ;
  assign CLBLM_R_X59Y98_SLICE_X88Y98_C3 = CLBLM_L_X50Y106_SLICE_X76Y106_AQ;
  assign CLBLM_R_X59Y98_SLICE_X88Y98_C4 = CLBLM_L_X60Y99_SLICE_X91Y99_AO5;
  assign CLBLM_R_X59Y98_SLICE_X88Y98_C5 = CLBLM_L_X64Y100_SLICE_X97Y100_AQ;
  assign CLBLM_R_X59Y98_SLICE_X88Y98_C6 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X59Y98_SLICE_X88Y98_CE = CLBLL_R_X57Y101_SLICE_X86Y101_BO6;
  assign CLBLM_R_X59Y98_SLICE_X88Y98_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X65Y98_SLICE_X99Y98_A5 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_R_X59Y98_SLICE_X88Y98_D1 = CLBLM_L_X50Y104_SLICE_X76Y104_AQ;
  assign CLBLM_R_X59Y98_SLICE_X88Y98_D2 = CLBLM_L_X60Y99_SLICE_X91Y99_AO5;
  assign CLBLM_R_X59Y98_SLICE_X88Y98_D3 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X59Y98_SLICE_X88Y98_D4 = CLBLM_L_X62Y100_SLICE_X92Y100_AQ;
  assign CLBLM_R_X59Y98_SLICE_X88Y98_D5 = CLBLM_R_X59Y97_SLICE_X89Y97_AQ;
  assign CLBLM_R_X59Y98_SLICE_X88Y98_D6 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X65Y98_SLICE_X99Y98_A6 = CLBLM_L_X56Y97_SLICE_X85Y97_AQ;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_D1 = CLBLM_L_X50Y107_SLICE_X76Y107_BQ;
  assign CLBLM_R_X59Y98_SLICE_X88Y98_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_B1 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_T1 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_B3 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_B4 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_D1 = CLBLM_L_X50Y106_SLICE_X76Y106_CQ;
  assign CLBLM_R_X65Y98_SLICE_X99Y98_B1 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_B5 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_B6 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_T1 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_C1 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_C2 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_C3 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_C4 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_D1 = CLBLM_L_X60Y110_SLICE_X91Y110_AQ;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_C5 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_T1 = 1'b1;
  assign CLBLM_R_X65Y98_SLICE_X99Y98_C6 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_D1 = CLBLM_R_X59Y102_SLICE_X89Y102_AQ;
  assign CLBLM_R_X65Y98_SLICE_X99Y98_CE = CLBLM_L_X60Y98_SLICE_X91Y98_BQ;
  assign CLBLM_R_X65Y98_SLICE_X99Y98_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_T1 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_D1 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_D2 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_D3 = 1'b1;
  assign CLBLM_L_X56Y98_SLICE_X85Y98_B6 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_D4 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_D5 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_D6 = 1'b1;
  assign CLBLM_L_X50Y109_SLICE_X77Y109_A1 = 1'b1;
  assign CLBLM_L_X50Y109_SLICE_X77Y109_A2 = CLBLL_R_X57Y101_SLICE_X87Y101_AQ;
  assign CLBLM_L_X50Y109_SLICE_X77Y109_A3 = CLBLL_R_X57Y100_SLICE_X87Y100_AQ;
  assign CLBLM_L_X50Y109_SLICE_X77Y109_A4 = CLBLL_R_X57Y101_SLICE_X87Y101_CQ;
  assign CLBLM_L_X50Y109_SLICE_X77Y109_A5 = CLBLL_R_X57Y100_SLICE_X87Y100_CQ;
  assign CLBLM_L_X50Y109_SLICE_X77Y109_A6 = 1'b1;
  assign CLBLM_L_X56Y98_SLICE_X85Y98_C1 = CLBLL_R_X57Y103_SLICE_X86Y103_AQ;
  assign CLBLM_L_X50Y109_SLICE_X77Y109_B1 = 1'b1;
  assign CLBLM_L_X50Y109_SLICE_X77Y109_B2 = CLBLL_R_X57Y101_SLICE_X87Y101_AQ;
  assign CLBLM_L_X50Y109_SLICE_X77Y109_B3 = CLBLM_L_X56Y101_SLICE_X85Y101_BQ;
  assign CLBLM_L_X50Y109_SLICE_X77Y109_B4 = CLBLM_L_X56Y101_SLICE_X85Y101_DQ;
  assign CLBLM_L_X50Y109_SLICE_X77Y109_B5 = CLBLL_R_X57Y101_SLICE_X87Y101_CQ;
  assign CLBLM_L_X50Y109_SLICE_X77Y109_B6 = 1'b1;
  assign CLBLM_L_X50Y109_SLICE_X77Y109_C1 = CLBLL_R_X57Y100_SLICE_X87Y100_BQ;
  assign CLBLM_L_X50Y109_SLICE_X77Y109_C2 = CLBLM_L_X56Y101_SLICE_X85Y101_BQ;
  assign CLBLM_L_X50Y109_SLICE_X77Y109_C3 = CLBLL_R_X57Y101_SLICE_X87Y101_DQ;
  assign CLBLM_L_X50Y109_SLICE_X77Y109_C4 = 1'b1;
  assign CLBLM_L_X50Y109_SLICE_X77Y109_C5 = CLBLM_L_X56Y101_SLICE_X85Y101_DQ;
  assign CLBLM_L_X50Y109_SLICE_X77Y109_C6 = 1'b1;
  assign CLBLM_R_X65Y98_SLICE_X99Y98_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X50Y109_SLICE_X77Y109_CIN = CLBLM_L_X50Y108_SLICE_X77Y108_COUT;
  assign CLBLM_L_X56Y98_SLICE_X85Y98_C5 = 1'b1;
  assign CLBLM_L_X50Y109_SLICE_X77Y109_D1 = CLBLL_R_X57Y100_SLICE_X87Y100_BQ;
  assign CLBLM_L_X50Y109_SLICE_X77Y109_D2 = CLBLL_R_X57Y99_SLICE_X86Y99_AQ;
  assign CLBLM_L_X50Y109_SLICE_X77Y109_D3 = 1'b1;
  assign CLBLM_L_X50Y109_SLICE_X77Y109_D4 = CLBLL_R_X57Y99_SLICE_X86Y99_BQ;
  assign CLBLM_L_X50Y109_SLICE_X77Y109_D5 = CLBLL_R_X57Y101_SLICE_X87Y101_DQ;
  assign CLBLM_L_X56Y98_SLICE_X85Y98_CE = CLBLM_L_X60Y98_SLICE_X91Y98_DQ;
  assign CLBLM_L_X50Y109_SLICE_X77Y109_D6 = 1'b1;
  assign CLBLM_L_X50Y109_SLICE_X76Y109_A1 = 1'b1;
  assign CLBLM_L_X50Y109_SLICE_X76Y109_A2 = CLBLL_R_X57Y101_SLICE_X87Y101_CQ;
  assign CLBLM_L_X56Y98_SLICE_X85Y98_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X50Y109_SLICE_X76Y109_A3 = 1'b1;
  assign CLBLM_L_X50Y109_SLICE_X76Y109_A4 = CLBLL_R_X57Y101_SLICE_X87Y101_AQ;
  assign CLBLM_L_X50Y109_SLICE_X76Y109_A5 = 1'b1;
  assign CLBLM_L_X50Y109_SLICE_X76Y109_A6 = 1'b1;
  assign CLBLM_L_X62Y108_SLICE_X92Y108_C3 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_R_X59Y99_SLICE_X89Y99_A1 = 1'b1;
  assign CLBLM_R_X59Y99_SLICE_X89Y99_A2 = CLBLM_R_X59Y100_SLICE_X89Y100_CQ;
  assign CLBLM_L_X50Y109_SLICE_X76Y109_AX = CLBLL_R_X57Y101_SLICE_X87Y101_CQ;
  assign CLBLM_L_X62Y108_SLICE_X92Y108_C4 = CLBLM_R_X59Y103_SLICE_X89Y103_CQ;
  assign CLBLM_L_X50Y109_SLICE_X76Y109_B1 = 1'b1;
  assign CLBLM_L_X50Y109_SLICE_X76Y109_B2 = 1'b1;
  assign CLBLM_L_X50Y109_SLICE_X76Y109_B3 = CLBLM_L_X56Y101_SLICE_X85Y101_BQ;
  assign CLBLM_L_X50Y109_SLICE_X76Y109_B4 = 1'b1;
  assign CLBLM_L_X50Y109_SLICE_X76Y109_B5 = CLBLM_L_X56Y101_SLICE_X85Y101_DQ;
  assign CLBLM_L_X50Y109_SLICE_X76Y109_B6 = 1'b1;
  assign CLBLM_L_X62Y108_SLICE_X92Y108_C5 = CLBLM_R_X59Y108_SLICE_X89Y108_AQ;
  assign CLBLM_R_X59Y99_SLICE_X89Y99_A5 = CLBLM_R_X49Y107_SLICE_X75Y107_CQ;
  assign CLBLM_L_X50Y109_SLICE_X76Y109_BX = CLBLM_L_X56Y101_SLICE_X85Y101_DQ;
  assign CLBLM_R_X59Y99_SLICE_X89Y99_B5 = CLBLM_R_X49Y107_SLICE_X75Y107_CQ;
  assign CLBLM_L_X50Y109_SLICE_X76Y109_C1 = CLBLL_R_X57Y100_SLICE_X87Y100_BQ;
  assign CLBLM_L_X50Y109_SLICE_X76Y109_C2 = 1'b1;
  assign CLBLM_L_X50Y109_SLICE_X76Y109_C3 = CLBLL_R_X57Y101_SLICE_X87Y101_DQ;
  assign CLBLM_L_X50Y109_SLICE_X76Y109_C4 = 1'b1;
  assign CLBLM_L_X50Y109_SLICE_X76Y109_C5 = 1'b1;
  assign CLBLM_L_X50Y109_SLICE_X76Y109_C6 = 1'b1;
  assign CLBLM_R_X59Y99_SLICE_X89Y99_C1 = CLBLM_L_X62Y99_SLICE_X92Y99_AO6;
  assign CLBLM_L_X50Y109_SLICE_X76Y109_CIN = CLBLM_L_X50Y108_SLICE_X76Y108_COUT;
  assign CLBLM_R_X59Y99_SLICE_X89Y99_C2 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X59Y99_SLICE_X89Y99_C3 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X59Y99_SLICE_X89Y99_C4 = CLBLM_L_X56Y99_SLICE_X84Y99_BQ;
  assign CLBLM_R_X59Y99_SLICE_X89Y99_C5 = 1'b1;
  assign CLBLM_R_X59Y99_SLICE_X89Y99_C6 = CLBLM_L_X56Y99_SLICE_X84Y99_AQ;
  assign CLBLM_L_X50Y109_SLICE_X76Y109_CX = CLBLL_R_X57Y101_SLICE_X87Y101_DQ;
  assign CLBLM_L_X56Y98_SLICE_X85Y98_D1 = CLBLL_R_X57Y102_SLICE_X86Y102_CO6;
  assign CLBLM_L_X50Y109_SLICE_X76Y109_D1 = 1'b1;
  assign CLBLM_L_X50Y109_SLICE_X76Y109_D2 = 1'b1;
  assign CLBLM_L_X50Y109_SLICE_X76Y109_D3 = 1'b1;
  assign CLBLM_L_X50Y109_SLICE_X76Y109_D4 = CLBLL_R_X57Y99_SLICE_X86Y99_BQ;
  assign CLBLM_L_X50Y109_SLICE_X76Y109_D5 = 1'b1;
  assign CLBLM_L_X50Y109_SLICE_X76Y109_D6 = CLBLL_R_X57Y99_SLICE_X86Y99_AQ;
  assign CLBLM_L_X56Y98_SLICE_X85Y98_D2 = CLBLM_L_X56Y98_SLICE_X84Y98_CO6;
  assign CLBLM_R_X59Y99_SLICE_X89Y99_D1 = 1'b1;
  assign CLBLM_L_X50Y109_SLICE_X76Y109_DX = CLBLL_R_X57Y99_SLICE_X86Y99_BQ;
  assign CLBLM_L_X56Y98_SLICE_X85Y98_D3 = CLBLM_L_X56Y98_SLICE_X84Y98_BO6;
  assign CLBLM_R_X59Y99_SLICE_X89Y99_D2 = 1'b1;
  assign CLBLM_R_X59Y99_SLICE_X89Y99_D3 = 1'b1;
  assign CLBLM_R_X59Y99_SLICE_X89Y99_D4 = 1'b1;
  assign CLBLM_L_X56Y98_SLICE_X85Y98_D4 = CLBLM_R_X49Y104_SLICE_X74Y104_AQ;
  assign CLBLM_R_X59Y99_SLICE_X89Y99_D5 = 1'b1;
  assign CLBLM_R_X59Y99_SLICE_X88Y99_A1 = CLBLM_R_X49Y107_SLICE_X75Y107_CQ;
  assign CLBLM_R_X59Y99_SLICE_X88Y99_A2 = CLBLM_L_X56Y99_SLICE_X84Y99_AQ;
  assign CLBLM_R_X59Y99_SLICE_X88Y99_A3 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLM_L_X56Y98_SLICE_X85Y98_D5 = CLBLM_R_X49Y104_SLICE_X75Y104_AQ;
  assign CLBLM_R_X59Y99_SLICE_X88Y99_A4 = CLBLM_R_X59Y100_SLICE_X89Y100_AQ;
  assign CLBLM_R_X59Y99_SLICE_X88Y99_A5 = 1'b1;
  assign CLBLM_R_X59Y99_SLICE_X88Y99_A6 = CLBLM_L_X56Y99_SLICE_X84Y99_BQ;
  assign CLBLM_L_X56Y98_SLICE_X85Y98_D6 = CLBLM_L_X56Y100_SLICE_X85Y100_BO6;
  assign CLBLM_R_X59Y99_SLICE_X88Y99_B1 = CLBLM_R_X49Y107_SLICE_X75Y107_CQ;
  assign CLBLM_R_X59Y99_SLICE_X88Y99_B2 = CLBLM_R_X59Y100_SLICE_X89Y100_BQ;
  assign CLBLM_R_X59Y99_SLICE_X88Y99_B3 = CLBLM_R_X59Y98_SLICE_X88Y98_CQ;
  assign CLBLM_R_X59Y99_SLICE_X88Y99_B4 = CLBLM_L_X56Y99_SLICE_X84Y99_AQ;
  assign CLBLM_R_X59Y99_SLICE_X88Y99_B5 = 1'b1;
  assign CLBLM_R_X59Y99_SLICE_X88Y99_B6 = 1'b1;
  assign CLBLM_R_X59Y99_SLICE_X88Y99_C1 = CLBLM_R_X59Y98_SLICE_X88Y98_DQ;
  assign CLBLM_R_X59Y99_SLICE_X88Y99_C2 = CLBLM_L_X56Y99_SLICE_X84Y99_BQ;
  assign CLBLM_R_X59Y99_SLICE_X88Y99_C3 = 1'b1;
  assign CLBLM_R_X59Y99_SLICE_X88Y99_C4 = CLBLM_R_X49Y108_SLICE_X75Y108_DQ;
  assign CLBLM_R_X59Y99_SLICE_X88Y99_C5 = CLBLM_R_X49Y107_SLICE_X75Y107_CQ;
  assign CLBLM_L_X56Y98_SLICE_X85Y98_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X59Y99_SLICE_X88Y99_C6 = CLBLM_L_X56Y99_SLICE_X84Y99_AQ;
  assign CLBLM_R_X59Y99_SLICE_X88Y99_CE = CLBLL_R_X57Y99_SLICE_X87Y99_BO6;
  assign CLBLM_R_X59Y99_SLICE_X88Y99_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X59Y99_SLICE_X88Y99_D1 = 1'b1;
  assign CLBLM_R_X59Y99_SLICE_X88Y99_D2 = CLBLM_R_X49Y107_SLICE_X75Y107_DQ;
  assign CLBLM_R_X59Y99_SLICE_X88Y99_D3 = CLBLM_R_X49Y107_SLICE_X75Y107_CQ;
  assign CLBLM_R_X59Y99_SLICE_X88Y99_D4 = CLBLM_L_X56Y99_SLICE_X84Y99_BQ;
  assign CLBLM_R_X59Y99_SLICE_X88Y99_D5 = CLBLM_R_X59Y98_SLICE_X88Y98_AQ;
  assign CLBLM_R_X59Y99_SLICE_X88Y99_D6 = CLBLM_L_X56Y99_SLICE_X84Y99_AQ;
  assign CLBLM_L_X56Y98_SLICE_X84Y98_A1 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLM_R_X59Y99_SLICE_X88Y99_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X56Y98_SLICE_X84Y98_A2 = 1'b1;
  assign CLBLM_L_X56Y98_SLICE_X84Y98_A3 = CLBLM_R_X49Y107_SLICE_X75Y107_DQ;
  assign CLBLM_L_X56Y98_SLICE_X84Y98_A4 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLM_L_X56Y98_SLICE_X84Y98_A5 = 1'b1;
  assign CLBLM_L_X62Y108_SLICE_X92Y108_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X56Y98_SLICE_X84Y98_A6 = 1'b1;
  assign CLBLM_L_X56Y98_SLICE_X84Y98_B1 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLM_L_X56Y98_SLICE_X84Y98_B2 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign CLBLM_L_X56Y98_SLICE_X84Y98_B3 = CLBLM_L_X56Y98_SLICE_X85Y98_BO5;
  assign CLBLM_L_X56Y98_SLICE_X84Y98_B4 = CLBLM_L_X56Y98_SLICE_X84Y98_DO5;
  assign CLBLM_L_X56Y98_SLICE_X84Y98_B5 = CLBLM_L_X56Y97_SLICE_X84Y97_AO6;
  assign CLBLM_L_X56Y98_SLICE_X84Y98_B6 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLL_R_X57Y105_SLICE_X86Y105_A6 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X56Y98_SLICE_X84Y98_C1 = CLBLM_R_X49Y107_SLICE_X75Y107_DQ;
  assign CLBLM_L_X56Y98_SLICE_X84Y98_C2 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLM_L_X56Y98_SLICE_X84Y98_C3 = CLBLM_R_X49Y108_SLICE_X75Y108_DQ;
  assign CLBLL_R_X57Y105_SLICE_X86Y105_B1 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X56Y98_SLICE_X84Y98_C4 = CLBLM_L_X56Y97_SLICE_X84Y97_CO5;
  assign CLBLL_R_X57Y105_SLICE_X86Y105_B2 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLL_R_X57Y105_SLICE_X86Y105_B4 = CLBLL_R_X57Y106_SLICE_X86Y106_C_XOR;
  assign CLBLL_R_X57Y105_SLICE_X86Y105_B5 = CLBLM_L_X62Y98_SLICE_X92Y98_AO6;
  assign CLBLL_R_X57Y105_SLICE_X86Y105_B6 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X50Y110_SLICE_X77Y110_A1 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X77Y110_A2 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X77Y110_A3 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X77Y110_A4 = CLBLL_R_X57Y99_SLICE_X86Y99_AQ;
  assign CLBLM_L_X50Y110_SLICE_X77Y110_A5 = CLBLL_R_X57Y99_SLICE_X86Y99_BQ;
  assign CLBLM_L_X50Y110_SLICE_X77Y110_A6 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X77Y110_AX = 1'b0;
  assign CLBLM_L_X50Y110_SLICE_X77Y110_B1 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X77Y110_B2 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X77Y110_B3 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X77Y110_B4 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X77Y110_B5 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X77Y110_B6 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X77Y110_BX = 1'b0;
  assign CLBLM_L_X50Y110_SLICE_X77Y110_C1 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X77Y110_C2 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X77Y110_C3 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X77Y110_C4 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X77Y110_C5 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X77Y110_C6 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X77Y110_CIN = CLBLM_L_X50Y109_SLICE_X77Y109_COUT;
  assign CLBLL_R_X57Y105_SLICE_X86Y105_C6 = CLBLL_R_X57Y109_SLICE_X86Y109_AQ;
  assign CLBLM_L_X50Y110_SLICE_X77Y110_CX = 1'b0;
  assign CLBLM_L_X50Y110_SLICE_X77Y110_D1 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X77Y110_D2 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X77Y110_D3 = 1'b1;
  assign CLBLL_R_X57Y105_SLICE_X86Y105_CE = CLBLM_L_X60Y100_SLICE_X90Y100_BO6;
  assign CLBLM_L_X50Y110_SLICE_X77Y110_D4 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X77Y110_D5 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X77Y110_D6 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X77Y110_DX = 1'b0;
  assign CLBLM_L_X50Y110_SLICE_X76Y110_A1 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X76Y110_A2 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X76Y110_A3 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X76Y110_A4 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X76Y110_A5 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X76Y110_A6 = 1'b1;
  assign CLBLM_R_X59Y100_SLICE_X89Y100_A1 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X59Y100_SLICE_X89Y100_A2 = CLBLM_L_X60Y99_SLICE_X91Y99_AO5;
  assign CLBLM_R_X59Y100_SLICE_X89Y100_A3 = CLBLM_R_X49Y106_SLICE_X74Y106_AQ;
  assign CLBLM_L_X50Y110_SLICE_X76Y110_AX = 1'b0;
  assign CLBLM_R_X59Y100_SLICE_X89Y100_A4 = CLBLM_R_X59Y100_SLICE_X88Y100_BQ;
  assign CLBLM_L_X50Y110_SLICE_X76Y110_B1 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X76Y110_B2 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X76Y110_B3 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X76Y110_B4 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X76Y110_B5 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X76Y110_B6 = 1'b1;
  assign CLBLM_R_X59Y100_SLICE_X89Y100_A5 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X59Y100_SLICE_X89Y100_A6 = CLBLM_L_X62Y100_SLICE_X92Y100_CQ;
  assign CLBLM_R_X59Y100_SLICE_X89Y100_B4 = CLBLM_R_X59Y100_SLICE_X88Y100_DQ;
  assign CLBLM_L_X50Y110_SLICE_X76Y110_BX = 1'b0;
  assign CLBLM_R_X59Y100_SLICE_X89Y100_B6 = CLBLM_L_X64Y100_SLICE_X97Y100_BQ;
  assign CLBLM_L_X50Y110_SLICE_X76Y110_C1 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X76Y110_C2 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X76Y110_C3 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X76Y110_C4 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X76Y110_C5 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X76Y110_C6 = 1'b1;
  assign CLBLM_R_X59Y100_SLICE_X89Y100_B5 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X59Y100_SLICE_X89Y100_C5 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X59Y100_SLICE_X89Y100_C6 = CLBLM_L_X50Y107_SLICE_X76Y107_BQ;
  assign CLBLM_R_X59Y100_SLICE_X89Y100_CE = CLBLL_R_X57Y101_SLICE_X86Y101_BO6;
  assign CLBLM_L_X50Y110_SLICE_X76Y110_CIN = CLBLM_L_X50Y109_SLICE_X76Y109_COUT;
  assign CLBLM_R_X59Y100_SLICE_X89Y100_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X59Y100_SLICE_X89Y100_C1 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X59Y100_SLICE_X89Y100_C2 = CLBLM_L_X60Y99_SLICE_X91Y99_AO5;
  assign CLBLM_R_X59Y100_SLICE_X89Y100_C3 = CLBLM_R_X59Y100_SLICE_X88Y100_B5Q;
  assign CLBLM_L_X50Y110_SLICE_X76Y110_CX = 1'b0;
  assign CLBLM_L_X50Y110_SLICE_X76Y110_D1 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X76Y110_D2 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X76Y110_D3 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X76Y110_D4 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X76Y110_D5 = 1'b1;
  assign CLBLM_L_X50Y110_SLICE_X76Y110_D6 = 1'b1;
  assign CLBLM_R_X59Y100_SLICE_X89Y100_D6 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X59Y100_SLICE_X89Y100_D1 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X50Y110_SLICE_X76Y110_DX = 1'b0;
  assign CLBLM_R_X59Y100_SLICE_X89Y100_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X59Y100_SLICE_X89Y100_D2 = CLBLM_L_X60Y99_SLICE_X91Y99_AO5;
  assign CLBLM_R_X59Y100_SLICE_X89Y100_D3 = CLBLM_L_X50Y107_SLICE_X77Y107_AQ;
  assign CLBLL_R_X57Y105_SLICE_X86Y105_D4 = CLBLL_R_X57Y109_SLICE_X86Y109_CQ;
  assign CLBLM_R_X59Y100_SLICE_X89Y100_D5 = CLBLM_R_X59Y100_SLICE_X88Y100_C5Q;
  assign CLBLM_R_X59Y100_SLICE_X88Y100_A1 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLL_R_X57Y105_SLICE_X86Y105_D5 = CLBLM_L_X56Y105_SLICE_X84Y105_AQ;
  assign CLBLM_R_X59Y100_SLICE_X88Y100_A3 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X59Y100_SLICE_X88Y100_A4 = CLBLM_L_X50Y104_SLICE_X76Y104_AQ;
  assign CLBLM_R_X59Y100_SLICE_X88Y100_A5 = CLBLM_R_X49Y104_SLICE_X74Y104_AQ;
  assign CLBLM_R_X59Y100_SLICE_X88Y100_A6 = 1'b1;
  assign CLBLM_R_X59Y100_SLICE_X88Y100_A2 = CLBLM_L_X60Y100_SLICE_X90Y100_AQ;
  assign CLBLM_R_X59Y100_SLICE_X88Y100_AX = CLBLM_R_X59Y98_SLICE_X88Y98_BQ;
  assign CLBLM_R_X59Y100_SLICE_X88Y100_B1 = 1'b1;
  assign CLBLM_R_X59Y100_SLICE_X88Y100_B2 = 1'b1;
  assign CLBLM_R_X59Y100_SLICE_X88Y100_B3 = 1'b1;
  assign CLBLM_R_X59Y100_SLICE_X88Y100_B4 = 1'b1;
  assign CLBLM_R_X59Y100_SLICE_X88Y100_B5 = 1'b1;
  assign CLBLM_R_X59Y100_SLICE_X88Y100_B6 = CLBLM_R_X59Y100_SLICE_X89Y100_AQ;
  assign CLBLM_R_X59Y100_SLICE_X88Y100_BX = CLBLM_R_X59Y100_SLICE_X89Y100_CQ;
  assign CLBLM_R_X59Y100_SLICE_X88Y100_C1 = 1'b1;
  assign CLBLM_R_X59Y100_SLICE_X88Y100_C2 = 1'b1;
  assign CLBLM_R_X59Y100_SLICE_X88Y100_C3 = 1'b1;
  assign CLBLM_R_X59Y100_SLICE_X88Y100_C4 = 1'b1;
  assign CLBLM_R_X59Y100_SLICE_X88Y100_C5 = 1'b1;
  assign CLBLM_R_X59Y100_SLICE_X88Y100_C6 = CLBLM_R_X59Y98_SLICE_X88Y98_CQ;
  assign CLBLM_R_X59Y100_SLICE_X88Y100_CE = CLBLL_R_X57Y97_SLICE_X87Y97_AO6;
  assign CLBLM_R_X59Y100_SLICE_X88Y100_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X59Y100_SLICE_X88Y100_CX = CLBLM_R_X59Y100_SLICE_X89Y100_DQ;
  assign CLBLM_R_X59Y100_SLICE_X88Y100_D1 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X59Y100_SLICE_X88Y100_D2 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X59Y100_SLICE_X88Y100_D3 = CLBLL_L_X54Y101_SLICE_X83Y101_AO6;
  assign CLBLM_R_X59Y100_SLICE_X88Y100_D4 = CLBLM_L_X64Y100_SLICE_X97Y100_BQ;
  assign CLBLM_R_X59Y100_SLICE_X88Y100_D5 = CLBLM_R_X59Y101_SLICE_X88Y101_CO6;
  assign CLBLM_R_X59Y100_SLICE_X88Y100_D6 = CLBLM_L_X64Y100_SLICE_X97Y100_AQ;
  assign CLBLM_R_X59Y100_SLICE_X88Y100_DX = CLBLM_R_X59Y100_SLICE_X89Y100_BQ;
  assign CLBLM_R_X59Y100_SLICE_X88Y100_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X59Y101_SLICE_X89Y101_C5 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_D1 = CLBLM_R_X49Y111_SLICE_X75Y111_AQ;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_T1 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_D1 = CLBLM_L_X50Y107_SLICE_X77Y107_AQ;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_T1 = 1'b1;
  assign CLBLL_R_X57Y105_SLICE_X87Y105_B1 = 1'b1;
  assign CLBLL_R_X57Y105_SLICE_X87Y105_B2 = 1'b1;
  assign CLBLM_L_X50Y111_SLICE_X77Y111_A1 = 1'b1;
  assign CLBLM_L_X50Y111_SLICE_X77Y111_A2 = 1'b1;
  assign CLBLM_L_X50Y111_SLICE_X77Y111_A3 = 1'b1;
  assign CLBLM_L_X50Y111_SLICE_X77Y111_A4 = 1'b1;
  assign CLBLL_R_X57Y105_SLICE_X87Y105_B3 = 1'b1;
  assign CLBLM_L_X50Y111_SLICE_X77Y111_A5 = 1'b1;
  assign CLBLM_L_X50Y111_SLICE_X77Y111_A6 = 1'b1;
  assign CLBLL_R_X57Y105_SLICE_X87Y105_B4 = 1'b1;
  assign CLBLM_L_X50Y111_SLICE_X77Y111_B1 = 1'b1;
  assign CLBLM_L_X50Y111_SLICE_X77Y111_B2 = 1'b1;
  assign CLBLM_L_X50Y111_SLICE_X77Y111_B3 = 1'b1;
  assign CLBLM_L_X50Y111_SLICE_X77Y111_B4 = 1'b1;
  assign CLBLM_L_X50Y111_SLICE_X77Y111_B5 = 1'b1;
  assign CLBLL_R_X57Y105_SLICE_X87Y105_B5 = CLBLL_R_X57Y105_SLICE_X86Y105_AQ;
  assign CLBLM_L_X50Y111_SLICE_X77Y111_B6 = 1'b1;
  assign CLBLL_R_X57Y105_SLICE_X87Y105_B6 = 1'b1;
  assign CLBLM_L_X50Y111_SLICE_X77Y111_C1 = 1'b1;
  assign CLBLM_L_X50Y111_SLICE_X77Y111_C2 = 1'b1;
  assign CLBLM_L_X50Y111_SLICE_X77Y111_C3 = 1'b1;
  assign CLBLM_L_X50Y111_SLICE_X77Y111_C4 = 1'b1;
  assign CLBLM_L_X50Y111_SLICE_X77Y111_C5 = 1'b1;
  assign CLBLM_L_X50Y111_SLICE_X77Y111_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_D1 = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_T1 = 1'b1;
  assign CLBLM_L_X50Y111_SLICE_X77Y111_D1 = 1'b1;
  assign CLBLM_L_X50Y111_SLICE_X77Y111_D2 = 1'b1;
  assign CLBLM_L_X50Y111_SLICE_X77Y111_D3 = 1'b1;
  assign CLBLM_L_X50Y111_SLICE_X77Y111_D4 = 1'b1;
  assign CLBLM_L_X50Y111_SLICE_X77Y111_D5 = 1'b1;
  assign CLBLM_L_X50Y111_SLICE_X77Y111_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_D1 = CLBLM_L_X56Y111_SLICE_X84Y111_AQ;
  assign CLBLM_L_X50Y111_SLICE_X76Y111_A1 = CLBLM_R_X49Y107_SLICE_X74Y107_DO6;
  assign CLBLM_L_X50Y111_SLICE_X76Y111_A2 = CLBLM_R_X49Y109_SLICE_X75Y109_C_XOR;
  assign CLBLM_L_X50Y111_SLICE_X76Y111_A3 = CLBLM_R_X49Y109_SLICE_X75Y109_B_XOR;
  assign CLBLM_L_X50Y111_SLICE_X76Y111_A4 = CLBLM_R_X49Y109_SLICE_X75Y109_D_XOR;
  assign CLBLM_L_X50Y111_SLICE_X76Y111_A5 = CLBLM_R_X49Y110_SLICE_X75Y110_A_CY;
  assign CLBLM_L_X50Y111_SLICE_X76Y111_A6 = CLBLL_L_X54Y100_SLICE_X82Y100_BQ;
  assign CLBLM_R_X59Y101_SLICE_X89Y101_A1 = CLBLM_R_X49Y107_SLICE_X75Y107_CQ;
  assign CLBLM_R_X59Y101_SLICE_X89Y101_A2 = CLBLM_R_X49Y106_SLICE_X75Y106_DQ;
  assign CLBLM_R_X59Y101_SLICE_X89Y101_A3 = CLBLM_L_X56Y102_SLICE_X85Y102_BO6;
  assign CLBLM_R_X59Y101_SLICE_X89Y101_A4 = CLBLM_R_X49Y104_SLICE_X75Y104_CQ;
  assign CLBLM_L_X50Y111_SLICE_X76Y111_B1 = 1'b1;
  assign CLBLM_L_X50Y111_SLICE_X76Y111_B2 = CLBLM_R_X53Y101_SLICE_X80Y101_BQ;
  assign CLBLM_L_X50Y111_SLICE_X76Y111_B3 = CLBLM_L_X50Y110_SLICE_X77Y110_A_XOR;
  assign CLBLM_L_X50Y111_SLICE_X76Y111_B4 = CLBLL_L_X54Y100_SLICE_X82Y100_BQ;
  assign CLBLM_L_X50Y111_SLICE_X76Y111_B5 = CLBLM_R_X53Y100_SLICE_X81Y100_AQ;
  assign CLBLM_L_X50Y111_SLICE_X76Y111_B6 = CLBLM_L_X50Y110_SLICE_X76Y110_A_CY;
  assign CLBLM_R_X59Y101_SLICE_X89Y101_B2 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_R_X59Y101_SLICE_X89Y101_B3 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X59Y101_SLICE_X89Y101_A5 = CLBLM_R_X49Y106_SLICE_X75Y106_CQ;
  assign CLBLM_R_X59Y101_SLICE_X89Y101_A6 = CLBLM_R_X49Y104_SLICE_X75Y104_DQ;
  assign CLBLM_R_X59Y101_SLICE_X89Y101_B1 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X50Y111_SLICE_X76Y111_C1 = CLBLM_R_X49Y109_SLICE_X75Y109_B_XOR;
  assign CLBLM_L_X50Y111_SLICE_X76Y111_C2 = CLBLM_R_X49Y107_SLICE_X74Y107_DO6;
  assign CLBLM_L_X50Y111_SLICE_X76Y111_C3 = CLBLM_R_X49Y109_SLICE_X75Y109_C_XOR;
  assign CLBLM_L_X50Y111_SLICE_X76Y111_C4 = CLBLL_L_X54Y100_SLICE_X82Y100_BQ;
  assign CLBLM_L_X50Y111_SLICE_X76Y111_C5 = CLBLM_L_X50Y111_SLICE_X76Y111_DO6;
  assign CLBLM_L_X50Y111_SLICE_X76Y111_C6 = 1'b1;
  assign CLBLM_R_X59Y101_SLICE_X89Y101_B6 = CLBLM_R_X59Y103_SLICE_X89Y103_CQ;
  assign CLBLM_R_X59Y101_SLICE_X89Y101_C6 = CLBLM_R_X59Y98_SLICE_X89Y98_BQ;
  assign CLBLM_R_X59Y101_SLICE_X89Y101_CE = CLBLM_L_X60Y98_SLICE_X91Y98_DQ;
  assign CLBLM_R_X59Y101_SLICE_X89Y101_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X59Y101_SLICE_X89Y101_C1 = CLBLM_R_X59Y98_SLICE_X88Y98_BQ;
  assign CLBLM_R_X59Y101_SLICE_X89Y101_C2 = CLBLM_R_X59Y111_SLICE_X89Y111_BQ;
  assign CLBLM_R_X59Y101_SLICE_X89Y101_C3 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_R_X59Y101_SLICE_X89Y101_C4 = CLBLM_R_X59Y105_SLICE_X89Y105_CQ;
  assign CLBLM_L_X50Y111_SLICE_X76Y111_D1 = CLBLM_L_X50Y109_SLICE_X77Y109_C_XOR;
  assign CLBLM_L_X50Y111_SLICE_X76Y111_D2 = CLBLM_L_X50Y109_SLICE_X76Y109_C_XOR;
  assign CLBLM_L_X50Y111_SLICE_X76Y111_D3 = 1'b1;
  assign CLBLM_L_X50Y111_SLICE_X76Y111_D4 = 1'b1;
  assign CLBLM_L_X50Y111_SLICE_X76Y111_D5 = 1'b1;
  assign CLBLM_L_X50Y111_SLICE_X76Y111_D6 = CLBLM_R_X53Y101_SLICE_X80Y101_BQ;
  assign CLBLM_R_X59Y101_SLICE_X89Y101_D1 = CLBLM_R_X59Y100_SLICE_X89Y100_AQ;
  assign CLBLM_R_X59Y101_SLICE_X89Y101_D2 = CLBLM_R_X59Y110_SLICE_X89Y110_AQ;
  assign CLBLM_R_X59Y101_SLICE_X89Y101_D3 = CLBLM_R_X59Y104_SLICE_X89Y104_CQ;
  assign CLBLM_R_X59Y101_SLICE_X89Y101_D4 = CLBLM_R_X59Y98_SLICE_X89Y98_B5Q;
  assign CLBLM_R_X59Y101_SLICE_X89Y101_D5 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_R_X59Y101_SLICE_X89Y101_D6 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_R_X59Y101_SLICE_X89Y101_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X59Y101_SLICE_X88Y101_A1 = CLBLM_L_X64Y100_SLICE_X97Y100_AQ;
  assign CLBLM_R_X59Y101_SLICE_X88Y101_A2 = CLBLL_L_X54Y101_SLICE_X83Y101_AO6;
  assign CLBLM_R_X59Y101_SLICE_X88Y101_A3 = CLBLM_L_X64Y100_SLICE_X97Y100_BQ;
  assign CLBLM_R_X59Y101_SLICE_X88Y101_A4 = CLBLM_R_X59Y101_SLICE_X88Y101_BO6;
  assign CLBLM_R_X59Y101_SLICE_X88Y101_A5 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X59Y101_SLICE_X88Y101_A6 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X59Y101_SLICE_X88Y101_B1 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X59Y101_SLICE_X88Y101_B2 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X59Y101_SLICE_X88Y101_B3 = CLBLM_R_X59Y103_SLICE_X89Y103_DQ;
  assign CLBLM_R_X59Y101_SLICE_X88Y101_B4 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_R_X59Y101_SLICE_X88Y101_B5 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_R_X59Y101_SLICE_X88Y101_B6 = CLBLM_R_X59Y103_SLICE_X89Y103_CQ;
  assign CLBLM_R_X59Y101_SLICE_X88Y101_C1 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_R_X59Y101_SLICE_X88Y101_C2 = CLBLM_R_X59Y103_SLICE_X89Y103_CQ;
  assign CLBLM_R_X59Y101_SLICE_X88Y101_C3 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X59Y101_SLICE_X88Y101_C4 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X59Y101_SLICE_X88Y101_C5 = CLBLM_R_X59Y103_SLICE_X89Y103_DQ;
  assign CLBLM_R_X59Y101_SLICE_X88Y101_C6 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_R_X59Y101_SLICE_X88Y101_D1 = CLBLM_R_X59Y111_SLICE_X89Y111_AQ;
  assign CLBLM_R_X59Y101_SLICE_X88Y101_D2 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_R_X59Y101_SLICE_X88Y101_D3 = CLBLM_R_X59Y106_SLICE_X89Y106_CQ;
  assign CLBLM_R_X59Y101_SLICE_X88Y101_D4 = CLBLM_R_X59Y98_SLICE_X89Y98_A5Q;
  assign CLBLM_R_X59Y101_SLICE_X88Y101_D5 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_R_X59Y101_SLICE_X88Y101_D6 = CLBLM_R_X59Y98_SLICE_X88Y98_AQ;
  assign CLBLM_R_X65Y107_SLICE_X99Y107_D5 = 1'b1;
  assign CLBLM_R_X59Y102_SLICE_X89Y102_A1 = CLBLM_R_X59Y103_SLICE_X89Y103_DQ;
  assign CLBLM_R_X59Y102_SLICE_X89Y102_A2 = CLBLM_R_X49Y104_SLICE_X75Y104_CQ;
  assign CLBLM_R_X59Y102_SLICE_X89Y102_A3 = CLBLM_R_X59Y106_SLICE_X89Y106_DO6;
  assign CLBLM_R_X59Y102_SLICE_X89Y102_A4 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X59Y102_SLICE_X89Y102_A5 = 1'b1;
  assign CLBLM_R_X59Y102_SLICE_X89Y102_A6 = CLBLM_L_X60Y102_SLICE_X90Y102_DO6;
  assign CLBLM_R_X59Y102_SLICE_X89Y102_B1 = CLBLL_R_X57Y105_SLICE_X86Y105_DO6;
  assign CLBLM_R_X59Y102_SLICE_X89Y102_B2 = CLBLM_R_X59Y101_SLICE_X89Y101_DO6;
  assign CLBLM_R_X59Y102_SLICE_X89Y102_B3 = CLBLM_L_X62Y106_SLICE_X93Y106_CO6;
  assign CLBLM_R_X59Y102_SLICE_X89Y102_B4 = CLBLM_R_X59Y102_SLICE_X89Y102_DO6;
  assign CLBLM_R_X59Y102_SLICE_X89Y102_B5 = CLBLM_L_X62Y103_SLICE_X93Y103_BO6;
  assign CLBLM_R_X59Y102_SLICE_X89Y102_B6 = CLBLM_L_X62Y107_SLICE_X93Y107_CO6;
  assign CLBLM_R_X59Y102_SLICE_X89Y102_C1 = CLBLM_R_X59Y97_SLICE_X88Y97_AQ;
  assign CLBLM_R_X59Y102_SLICE_X89Y102_C2 = CLBLM_L_X60Y109_SLICE_X91Y109_AQ;
  assign CLBLM_R_X59Y102_SLICE_X89Y102_C3 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_R_X59Y102_SLICE_X89Y102_C4 = 1'b1;
  assign CLBLM_R_X59Y102_SLICE_X89Y102_C5 = CLBLM_L_X60Y102_SLICE_X90Y102_CQ;
  assign CLBLM_R_X59Y102_SLICE_X89Y102_C6 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_R_X59Y102_SLICE_X89Y102_CE = CLBLM_R_X59Y99_SLICE_X89Y99_CO6;
  assign CLBLM_R_X59Y102_SLICE_X89Y102_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X59Y102_SLICE_X89Y102_D1 = CLBLM_L_X60Y102_SLICE_X90Y102_AQ;
  assign CLBLM_R_X59Y102_SLICE_X89Y102_D2 = 1'b1;
  assign CLBLM_R_X59Y102_SLICE_X89Y102_D3 = CLBLM_R_X59Y96_SLICE_X88Y96_BQ;
  assign CLBLM_R_X59Y102_SLICE_X89Y102_D4 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_R_X59Y102_SLICE_X89Y102_D5 = CLBLM_L_X60Y109_SLICE_X91Y109_BQ;
  assign CLBLM_R_X59Y102_SLICE_X89Y102_D6 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_R_X59Y102_SLICE_X89Y102_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X59Y102_SLICE_X88Y102_A1 = CLBLM_R_X59Y103_SLICE_X89Y103_DQ;
  assign CLBLM_R_X59Y102_SLICE_X88Y102_A2 = CLBLM_R_X49Y104_SLICE_X74Y104_AQ;
  assign CLBLM_R_X59Y102_SLICE_X88Y102_A3 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X59Y102_SLICE_X88Y102_A4 = CLBLM_R_X59Y102_SLICE_X88Y102_BO6;
  assign CLBLM_R_X59Y102_SLICE_X88Y102_A5 = CLBLM_L_X62Y106_SLICE_X92Y106_AO5;
  assign CLBLM_R_X59Y102_SLICE_X88Y102_A6 = CLBLM_R_X59Y103_SLICE_X88Y103_F7AMUX_O;
  assign CLBLM_R_X59Y102_SLICE_X88Y102_B1 = CLBLL_R_X57Y109_SLICE_X87Y109_A_XOR;
  assign CLBLM_R_X59Y102_SLICE_X88Y102_B2 = CLBLL_R_X57Y101_SLICE_X86Y101_AQ;
  assign CLBLM_R_X59Y102_SLICE_X88Y102_B3 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_R_X59Y102_SLICE_X88Y102_B4 = CLBLM_R_X59Y103_SLICE_X88Y103_BQ;
  assign CLBLM_R_X59Y102_SLICE_X88Y102_B5 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_R_X59Y102_SLICE_X88Y102_B6 = CLBLM_R_X59Y103_SLICE_X89Y103_CQ;
  assign CLBLM_R_X59Y102_SLICE_X88Y102_C1 = CLBLM_R_X63Y100_SLICE_X94Y100_AQ;
  assign CLBLM_R_X59Y102_SLICE_X88Y102_C2 = CLBLM_L_X60Y101_SLICE_X90Y101_AQ;
  assign CLBLM_R_X59Y102_SLICE_X88Y102_C3 = CLBLL_R_X57Y97_SLICE_X86Y97_AQ;
  assign CLBLM_R_X59Y102_SLICE_X88Y102_C4 = CLBLM_L_X62Y102_SLICE_X92Y102_BQ;
  assign CLBLM_R_X59Y102_SLICE_X88Y102_C5 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_R_X59Y102_SLICE_X88Y102_C6 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_R_X59Y102_SLICE_X88Y102_CE = CLBLM_R_X59Y99_SLICE_X89Y99_CO6;
  assign CLBLM_R_X59Y102_SLICE_X88Y102_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X59Y102_SLICE_X88Y102_D1 = CLBLM_R_X59Y101_SLICE_X88Y101_DO6;
  assign CLBLM_R_X59Y102_SLICE_X88Y102_D2 = CLBLM_R_X59Y102_SLICE_X89Y102_CO6;
  assign CLBLM_R_X59Y102_SLICE_X88Y102_D3 = CLBLM_R_X63Y103_SLICE_X94Y103_AO6;
  assign CLBLM_R_X59Y102_SLICE_X88Y102_D4 = CLBLM_L_X62Y103_SLICE_X93Y103_BO6;
  assign CLBLM_R_X59Y102_SLICE_X88Y102_D5 = CLBLL_R_X57Y105_SLICE_X86Y105_CO6;
  assign CLBLM_R_X59Y102_SLICE_X88Y102_D6 = CLBLM_L_X62Y106_SLICE_X93Y106_CO6;
  assign CLBLM_R_X59Y102_SLICE_X88Y102_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_D1 = CLBLM_L_X62Y110_SLICE_X92Y110_BQ;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_D1 = CLBLM_L_X60Y111_SLICE_X90Y111_AQ;
  assign CLBLM_R_X59Y103_SLICE_X89Y103_A1 = CLBLM_R_X59Y103_SLICE_X88Y103_DQ;
  assign CLBLM_R_X59Y103_SLICE_X89Y103_A2 = CLBLM_R_X59Y104_SLICE_X89Y104_DO6;
  assign CLBLM_R_X59Y103_SLICE_X89Y103_A3 = CLBLM_R_X59Y103_SLICE_X88Y103_BQ;
  assign CLBLM_R_X59Y103_SLICE_X89Y103_A4 = CLBLM_R_X59Y103_SLICE_X88Y103_CQ;
  assign CLBLM_R_X59Y103_SLICE_X89Y103_A5 = CLBLM_R_X59Y104_SLICE_X88Y104_AO6;
  assign CLBLM_R_X59Y103_SLICE_X89Y103_A6 = CLBLM_R_X59Y104_SLICE_X88Y104_AO5;
  assign CLBLM_R_X59Y103_SLICE_X89Y103_AX = CLBLL_R_X57Y102_SLICE_X86Y102_AO5;
  assign CLBLM_R_X59Y103_SLICE_X89Y103_B1 = CLBLM_R_X59Y103_SLICE_X88Y103_DQ;
  assign CLBLM_R_X59Y103_SLICE_X89Y103_B2 = CLBLM_R_X59Y104_SLICE_X89Y104_DO6;
  assign CLBLM_R_X59Y103_SLICE_X89Y103_B3 = CLBLM_R_X59Y104_SLICE_X88Y104_AO6;
  assign CLBLM_R_X59Y103_SLICE_X89Y103_B4 = CLBLM_R_X59Y103_SLICE_X88Y103_BQ;
  assign CLBLM_R_X59Y103_SLICE_X89Y103_B5 = CLBLM_R_X59Y103_SLICE_X88Y103_CQ;
  assign CLBLM_R_X59Y103_SLICE_X89Y103_B6 = CLBLM_R_X59Y104_SLICE_X88Y104_AO5;
  assign CLBLM_R_X59Y103_SLICE_X89Y103_C1 = CLBLM_R_X59Y104_SLICE_X88Y104_AO6;
  assign CLBLM_R_X59Y103_SLICE_X89Y103_C2 = CLBLM_R_X59Y104_SLICE_X88Y104_AO5;
  assign CLBLM_R_X59Y103_SLICE_X89Y103_C3 = CLBLM_R_X59Y104_SLICE_X89Y104_DO6;
  assign CLBLM_R_X59Y103_SLICE_X89Y103_C4 = CLBLM_R_X59Y103_SLICE_X88Y103_CQ;
  assign CLBLM_R_X59Y103_SLICE_X89Y103_C5 = CLBLM_R_X59Y103_SLICE_X88Y103_DQ;
  assign CLBLM_R_X59Y103_SLICE_X89Y103_C6 = CLBLM_R_X59Y103_SLICE_X88Y103_BQ;
  assign CLBLM_R_X59Y103_SLICE_X89Y103_CE = CLBLM_L_X60Y98_SLICE_X91Y98_DQ;
  assign CLBLM_R_X59Y103_SLICE_X89Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X59Y103_SLICE_X89Y103_D1 = CLBLM_R_X59Y104_SLICE_X88Y104_AO6;
  assign CLBLM_R_X59Y103_SLICE_X89Y103_D2 = CLBLM_R_X59Y104_SLICE_X88Y104_AO5;
  assign CLBLM_R_X59Y103_SLICE_X89Y103_D3 = 1'b1;
  assign CLBLM_R_X59Y103_SLICE_X89Y103_D4 = CLBLM_R_X59Y103_SLICE_X88Y103_CQ;
  assign CLBLM_R_X59Y103_SLICE_X89Y103_D5 = CLBLM_R_X59Y103_SLICE_X88Y103_DQ;
  assign CLBLM_R_X59Y103_SLICE_X89Y103_D6 = CLBLM_R_X59Y103_SLICE_X88Y103_BQ;
  assign CLBLM_R_X59Y103_SLICE_X89Y103_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X59Y103_SLICE_X88Y103_A1 = CLBLM_L_X60Y105_SLICE_X90Y105_A_XOR;
  assign CLBLM_R_X59Y103_SLICE_X88Y103_A2 = CLBLM_L_X62Y102_SLICE_X92Y102_BQ;
  assign CLBLM_R_X59Y103_SLICE_X88Y103_A3 = CLBLM_L_X60Y100_SLICE_X90Y100_AQ;
  assign CLBLM_R_X59Y103_SLICE_X88Y103_A4 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_R_X59Y103_SLICE_X88Y103_A5 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_R_X59Y103_SLICE_X88Y103_A6 = CLBLM_R_X59Y103_SLICE_X89Y103_CQ;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_T1 = 1'b1;
  assign CLBLM_R_X59Y103_SLICE_X88Y103_AX = CLBLM_R_X59Y103_SLICE_X89Y103_DQ;
  assign CLBLM_R_X59Y103_SLICE_X88Y103_B1 = CLBLM_R_X59Y108_SLICE_X88Y108_A_XOR;
  assign CLBLM_R_X59Y103_SLICE_X88Y103_B2 = 1'b1;
  assign CLBLM_R_X59Y103_SLICE_X88Y103_B3 = CLBLM_L_X60Y100_SLICE_X90Y100_AQ;
  assign CLBLM_R_X59Y103_SLICE_X88Y103_B4 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_R_X59Y103_SLICE_X88Y103_B5 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_R_X59Y103_SLICE_X88Y103_B6 = CLBLM_R_X59Y103_SLICE_X89Y103_CQ;
  assign CLBLM_R_X59Y103_SLICE_X88Y103_BX = CLBLM_R_X49Y104_SLICE_X74Y104_AQ;
  assign CLBLM_R_X59Y103_SLICE_X88Y103_C1 = CLBLM_L_X62Y106_SLICE_X93Y106_CO6;
  assign CLBLM_R_X59Y103_SLICE_X88Y103_C2 = CLBLM_R_X59Y102_SLICE_X88Y102_CO6;
  assign CLBLM_R_X59Y103_SLICE_X88Y103_C3 = CLBLL_R_X57Y104_SLICE_X86Y104_DO6;
  assign CLBLM_R_X59Y103_SLICE_X88Y103_C4 = CLBLM_R_X59Y104_SLICE_X88Y104_DO6;
  assign CLBLM_R_X59Y103_SLICE_X88Y103_C5 = CLBLM_R_X59Y103_SLICE_X88Y103_DO6;
  assign CLBLM_R_X59Y103_SLICE_X88Y103_C6 = CLBLM_L_X62Y103_SLICE_X93Y103_BO6;
  assign CLBLM_R_X59Y103_SLICE_X88Y103_CE = CLBLL_R_X57Y99_SLICE_X87Y99_BO6;
  assign CLBLM_R_X59Y103_SLICE_X88Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X59Y103_SLICE_X88Y103_CX = CLBLM_R_X49Y104_SLICE_X75Y104_AQ;
  assign CLBLM_R_X59Y103_SLICE_X88Y103_D1 = CLBLM_L_X60Y100_SLICE_X90Y100_AQ;
  assign CLBLM_R_X59Y103_SLICE_X88Y103_D2 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_R_X59Y103_SLICE_X88Y103_D3 = CLBLM_R_X59Y111_SLICE_X89Y111_CQ;
  assign CLBLM_R_X59Y103_SLICE_X88Y103_D4 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_R_X59Y103_SLICE_X88Y103_D5 = CLBLM_R_X59Y98_SLICE_X88Y98_DQ;
  assign CLBLM_R_X59Y103_SLICE_X88Y103_D6 = CLBLM_R_X59Y98_SLICE_X89Y98_AQ;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_A4 = CLBLM_R_X65Y99_SLICE_X99Y99_BO6;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_A5 = CLBLM_R_X65Y97_SLICE_X98Y97_AO6;
  assign CLBLM_R_X59Y103_SLICE_X88Y103_DX = CLBLM_R_X49Y104_SLICE_X75Y104_BQ;
  assign CLBLM_R_X59Y103_SLICE_X88Y103_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_D1 = CLBLM_L_X50Y105_SLICE_X77Y105_AQ;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_B3 = 1'b1;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_B4 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_B6 = CLBLM_L_X56Y97_SLICE_X85Y97_AQ;
  assign CLBLM_L_X62Y109_SLICE_X93Y109_D4 = 1'b1;
  assign CLBLM_L_X62Y109_SLICE_X93Y109_D5 = 1'b1;
  assign CLBLM_L_X62Y109_SLICE_X93Y109_D6 = 1'b1;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_C1 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_T1 = 1'b1;
  assign CLBLM_R_X65Y99_SLICE_X99Y99_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign RIOB33_X105Y107_IOB_X1Y108_O = CLBLM_R_X65Y100_SLICE_X99Y100_CQ;
  assign RIOB33_X105Y107_IOB_X1Y107_O = 1'b0;
  assign CLBLM_L_X62Y109_SLICE_X92Y109_B1 = CLBLL_R_X57Y102_SLICE_X86Y102_AQ;
  assign CLBLM_L_X62Y109_SLICE_X92Y109_B2 = CLBLM_L_X60Y98_SLICE_X90Y98_BQ;
  assign CLBLM_L_X62Y109_SLICE_X92Y109_B3 = CLBLM_R_X59Y102_SLICE_X88Y102_AQ;
  assign CLBLM_L_X62Y109_SLICE_X92Y109_B4 = CLBLM_L_X56Y103_SLICE_X85Y103_CO6;
  assign CLBLM_L_X62Y109_SLICE_X92Y109_B5 = CLBLL_R_X57Y102_SLICE_X86Y102_BQ;
  assign CLBLM_L_X56Y99_SLICE_X85Y99_C1 = CLBLM_R_X49Y106_SLICE_X75Y106_CQ;
  assign CLBLM_L_X62Y109_SLICE_X92Y109_B6 = CLBLM_L_X62Y109_SLICE_X92Y109_CO6;
  assign CLBLM_L_X56Y99_SLICE_X85Y99_C5 = CLBLM_R_X49Y104_SLICE_X75Y104_AQ;
  assign CLBLM_L_X56Y99_SLICE_X85Y99_CE = CLBLM_L_X60Y98_SLICE_X91Y98_DQ;
  assign CLBLM_L_X62Y109_SLICE_X92Y109_C1 = CLBLM_L_X62Y103_SLICE_X92Y103_AQ;
  assign CLBLM_R_X59Y104_SLICE_X89Y104_A1 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_R_X59Y104_SLICE_X89Y104_A2 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_R_X59Y104_SLICE_X89Y104_A3 = CLBLM_R_X59Y106_SLICE_X88Y106_AQ;
  assign CLBLM_L_X62Y109_SLICE_X92Y109_C2 = CLBLM_L_X62Y106_SLICE_X93Y106_AQ;
  assign CLBLM_R_X59Y104_SLICE_X89Y104_A4 = CLBLL_R_X57Y104_SLICE_X87Y104_BQ;
  assign CLBLM_L_X56Y99_SLICE_X85Y99_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X59Y104_SLICE_X89Y104_A5 = CLBLM_L_X60Y107_SLICE_X90Y107_AQ;
  assign CLBLM_R_X59Y104_SLICE_X89Y104_A6 = CLBLM_L_X56Y104_SLICE_X85Y104_AQ;
  assign CLBLM_L_X62Y109_SLICE_X92Y109_C3 = CLBLM_L_X62Y104_SLICE_X93Y104_AQ;
  assign CLBLM_R_X59Y104_SLICE_X89Y104_AX = CLBLM_L_X62Y106_SLICE_X93Y106_CO6;
  assign CLBLM_R_X59Y104_SLICE_X89Y104_B1 = CLBLM_L_X64Y106_SLICE_X96Y106_BQ;
  assign CLBLM_R_X59Y104_SLICE_X89Y104_B2 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_R_X59Y104_SLICE_X89Y104_B3 = 1'b1;
  assign CLBLM_R_X59Y104_SLICE_X89Y104_B4 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_R_X59Y104_SLICE_X89Y104_B5 = CLBLM_L_X64Y108_SLICE_X96Y108_BQ;
  assign CLBLM_R_X59Y104_SLICE_X89Y104_B6 = CLBLM_R_X49Y109_SLICE_X74Y109_CQ;
  assign CLBLM_L_X62Y109_SLICE_X92Y109_C4 = CLBLM_L_X60Y110_SLICE_X91Y110_AQ;
  assign CLBLM_L_X62Y109_SLICE_X92Y109_C5 = CLBLM_L_X62Y110_SLICE_X92Y110_DO6;
  assign CLBLM_R_X59Y104_SLICE_X89Y104_C1 = CLBLM_L_X60Y108_SLICE_X90Y108_C_XOR;
  assign CLBLM_R_X59Y104_SLICE_X89Y104_C2 = CLBLM_L_X62Y98_SLICE_X92Y98_AO6;
  assign CLBLM_R_X59Y104_SLICE_X89Y104_C3 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_R_X59Y104_SLICE_X89Y104_C4 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X59Y104_SLICE_X89Y104_C5 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X59Y104_SLICE_X89Y104_C6 = CLBLM_R_X59Y107_SLICE_X89Y107_C_XOR;
  assign CLBLM_R_X59Y104_SLICE_X89Y104_CE = CLBLM_L_X60Y99_SLICE_X90Y99_DO6;
  assign CLBLM_L_X62Y109_SLICE_X92Y109_C6 = CLBLM_R_X59Y102_SLICE_X89Y102_AQ;
  assign CLBLM_R_X59Y104_SLICE_X89Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X59Y104_SLICE_X89Y104_D1 = 1'b1;
  assign CLBLM_R_X59Y104_SLICE_X89Y104_D2 = CLBLM_R_X59Y107_SLICE_X89Y107_BQ;
  assign CLBLM_R_X59Y104_SLICE_X89Y104_D3 = CLBLM_R_X59Y104_SLICE_X88Y104_BO6;
  assign CLBLM_R_X59Y104_SLICE_X89Y104_D4 = 1'b1;
  assign CLBLM_R_X59Y104_SLICE_X89Y104_D5 = 1'b1;
  assign CLBLM_R_X59Y104_SLICE_X89Y104_D6 = CLBLM_R_X59Y104_SLICE_X88Y104_BQ;
  assign CLBLM_L_X56Y99_SLICE_X85Y99_D1 = 1'b1;
  assign CLBLM_R_X59Y104_SLICE_X89Y104_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X56Y99_SLICE_X85Y99_D2 = 1'b1;
  assign CLBLM_R_X59Y104_SLICE_X88Y104_A1 = CLBLM_R_X59Y107_SLICE_X89Y107_BQ;
  assign CLBLM_R_X59Y104_SLICE_X88Y104_A2 = CLBLM_R_X59Y104_SLICE_X88Y104_BQ;
  assign CLBLM_R_X59Y104_SLICE_X88Y104_A3 = CLBLM_R_X59Y104_SLICE_X88Y104_AQ;
  assign CLBLM_L_X56Y99_SLICE_X85Y99_D3 = 1'b1;
  assign CLBLM_R_X59Y104_SLICE_X88Y104_A5 = CLBLM_R_X59Y104_SLICE_X88Y104_CO6;
  assign CLBLM_R_X59Y104_SLICE_X88Y104_A6 = 1'b1;
  assign CLBLM_R_X59Y104_SLICE_X88Y104_A4 = CLBLM_R_X59Y104_SLICE_X88Y104_BO6;
  assign CLBLM_L_X56Y99_SLICE_X85Y99_D4 = 1'b1;
  assign CLBLM_R_X59Y104_SLICE_X88Y104_AX = CLBLM_R_X49Y104_SLICE_X75Y104_CQ;
  assign CLBLM_R_X59Y104_SLICE_X88Y104_B1 = CLBLM_R_X59Y106_SLICE_X88Y106_DO6;
  assign CLBLM_R_X59Y104_SLICE_X88Y104_B2 = CLBLM_R_X59Y99_SLICE_X89Y99_AQ;
  assign CLBLM_R_X59Y104_SLICE_X88Y104_B3 = CLBLM_R_X59Y104_SLICE_X88Y104_AQ;
  assign CLBLM_R_X59Y104_SLICE_X88Y104_B4 = CLBLM_R_X59Y99_SLICE_X89Y99_A5Q;
  assign CLBLM_R_X59Y104_SLICE_X88Y104_B5 = CLBLM_R_X59Y99_SLICE_X88Y99_BQ;
  assign CLBLM_R_X59Y104_SLICE_X88Y104_B6 = CLBLM_R_X59Y99_SLICE_X88Y99_B5Q;
  assign CLBLM_L_X56Y99_SLICE_X85Y99_D5 = 1'b1;
  assign CLBLM_L_X56Y99_SLICE_X85Y99_D6 = 1'b1;
  assign CLBLM_R_X59Y104_SLICE_X88Y104_BX = CLBLM_R_X49Y106_SLICE_X75Y106_CQ;
  assign CLBLM_R_X59Y104_SLICE_X88Y104_C1 = CLBLM_R_X59Y99_SLICE_X88Y99_BQ;
  assign CLBLM_R_X59Y104_SLICE_X88Y104_C2 = 1'b1;
  assign CLBLM_R_X59Y104_SLICE_X88Y104_C3 = CLBLM_R_X59Y99_SLICE_X89Y99_A5Q;
  assign CLBLM_R_X59Y104_SLICE_X88Y104_C4 = CLBLM_R_X59Y99_SLICE_X88Y99_B5Q;
  assign CLBLM_R_X59Y104_SLICE_X88Y104_C5 = CLBLM_R_X59Y106_SLICE_X88Y106_DO6;
  assign CLBLM_R_X59Y104_SLICE_X88Y104_C6 = CLBLM_R_X59Y99_SLICE_X89Y99_AQ;
  assign CLBLM_R_X59Y104_SLICE_X88Y104_CE = CLBLL_R_X57Y99_SLICE_X87Y99_BO6;
  assign CLBLM_R_X59Y104_SLICE_X88Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X62Y109_SLICE_X92Y109_D1 = 1'b1;
  assign CLBLM_L_X62Y109_SLICE_X92Y109_D2 = 1'b1;
  assign CLBLM_R_X59Y104_SLICE_X88Y104_D1 = 1'b1;
  assign CLBLM_R_X59Y104_SLICE_X88Y104_D2 = CLBLM_L_X62Y105_SLICE_X92Y105_CQ;
  assign CLBLM_R_X59Y104_SLICE_X88Y104_D3 = CLBLM_R_X49Y109_SLICE_X74Y109_DQ;
  assign CLBLM_R_X59Y104_SLICE_X88Y104_D4 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_R_X59Y104_SLICE_X88Y104_D5 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_R_X59Y104_SLICE_X88Y104_D6 = CLBLM_L_X64Y107_SLICE_X97Y107_BQ;
  assign CLBLM_L_X56Y99_SLICE_X85Y99_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X62Y109_SLICE_X92Y109_D3 = 1'b1;
  assign CLBLM_L_X62Y109_SLICE_X92Y109_D4 = 1'b1;
  assign CLBLM_R_X59Y104_SLICE_X88Y104_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X62Y109_SLICE_X92Y109_D5 = 1'b1;
  assign CLBLM_L_X62Y109_SLICE_X92Y109_D6 = 1'b1;
  assign CLBLM_L_X56Y99_SLICE_X84Y99_A2 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLM_L_X56Y99_SLICE_X84Y99_A3 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLM_L_X56Y99_SLICE_X84Y99_A4 = CLBLL_L_X54Y98_SLICE_X82Y98_AO6;
  assign CLBLM_L_X56Y99_SLICE_X84Y99_A5 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign CLBLM_L_X56Y99_SLICE_X84Y99_A6 = CLBLM_R_X49Y108_SLICE_X75Y108_DQ;
  assign CLBLM_L_X56Y99_SLICE_X84Y99_B1 = 1'b1;
  assign CLBLM_L_X56Y99_SLICE_X84Y99_B2 = CLBLL_L_X54Y98_SLICE_X82Y98_AO6;
  assign CLBLM_L_X56Y99_SLICE_X84Y99_B3 = 1'b1;
  assign CLBLL_R_X57Y106_SLICE_X86Y106_A5 = 1'b1;
  assign CLBLM_L_X56Y99_SLICE_X84Y99_B4 = 1'b1;
  assign CLBLL_R_X57Y106_SLICE_X86Y106_A6 = 1'b1;
  assign CLBLM_L_X56Y99_SLICE_X84Y99_B5 = 1'b1;
  assign CLBLM_L_X56Y99_SLICE_X84Y99_B6 = 1'b1;
  assign RIOB33_X105Y109_IOB_X1Y110_O = CLBLM_R_X65Y106_SLICE_X98Y106_CQ;
  assign RIOB33_X105Y109_IOB_X1Y109_O = CLBLM_R_X65Y100_SLICE_X99Y100_AQ;
  assign CLBLL_R_X57Y106_SLICE_X86Y106_B6 = CLBLL_R_X57Y105_SLICE_X86Y105_AQ;
  assign CLBLM_L_X56Y99_SLICE_X84Y99_C6 = CLBLM_R_X49Y108_SLICE_X75Y108_DQ;
  assign CLBLM_L_X56Y99_SLICE_X84Y99_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X59Y105_SLICE_X89Y105_A1 = CLBLM_L_X56Y105_SLICE_X85Y105_CQ;
  assign CLBLM_R_X59Y105_SLICE_X89Y105_A2 = CLBLM_L_X56Y105_SLICE_X84Y105_CQ;
  assign CLBLM_R_X59Y105_SLICE_X89Y105_A3 = CLBLL_R_X57Y108_SLICE_X87Y108_BQ;
  assign CLBLM_R_X59Y105_SLICE_X89Y105_A4 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_R_X59Y105_SLICE_X89Y105_A5 = CLBLM_R_X59Y108_SLICE_X88Y108_AQ;
  assign CLBLM_R_X59Y105_SLICE_X89Y105_A6 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_R_X59Y105_SLICE_X89Y105_AX = CLBLM_L_X62Y106_SLICE_X93Y106_CO6;
  assign CLBLM_R_X59Y105_SLICE_X89Y105_B1 = CLBLM_R_X49Y111_SLICE_X74Y111_CQ;
  assign CLBLM_R_X59Y105_SLICE_X89Y105_B2 = 1'b1;
  assign CLBLM_R_X59Y105_SLICE_X89Y105_B3 = CLBLM_R_X63Y110_SLICE_X94Y110_AQ;
  assign CLBLM_R_X59Y105_SLICE_X89Y105_B4 = CLBLM_L_X64Y106_SLICE_X96Y106_AQ;
  assign CLBLM_R_X59Y105_SLICE_X89Y105_B5 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_R_X59Y105_SLICE_X89Y105_B6 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLL_R_X57Y106_SLICE_X86Y106_D2 = 1'b1;
  assign CLBLM_R_X59Y105_SLICE_X89Y105_C1 = CLBLM_L_X60Y108_SLICE_X90Y108_B_XOR;
  assign CLBLM_R_X59Y105_SLICE_X89Y105_C2 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X59Y105_SLICE_X89Y105_C3 = CLBLM_R_X59Y107_SLICE_X89Y107_B_XOR;
  assign CLBLM_R_X59Y105_SLICE_X89Y105_C4 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X59Y105_SLICE_X89Y105_C5 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_R_X59Y105_SLICE_X89Y105_C6 = CLBLM_L_X62Y105_SLICE_X92Y105_AO6;
  assign CLBLM_R_X59Y105_SLICE_X89Y105_CE = CLBLM_L_X60Y99_SLICE_X90Y99_DO6;
  assign CLBLM_R_X59Y105_SLICE_X89Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X59Y105_SLICE_X89Y105_D1 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_R_X59Y105_SLICE_X89Y105_D2 = CLBLM_R_X59Y108_SLICE_X89Y108_AQ;
  assign CLBLM_R_X59Y105_SLICE_X89Y105_D3 = CLBLM_R_X59Y96_SLICE_X89Y96_AQ;
  assign CLBLM_R_X59Y105_SLICE_X89Y105_D4 = CLBLM_R_X59Y100_SLICE_X89Y100_CQ;
  assign CLBLM_R_X59Y105_SLICE_X89Y105_D5 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_R_X59Y105_SLICE_X89Y105_D6 = CLBLM_R_X59Y112_SLICE_X89Y112_BQ;
  assign CLBLM_R_X59Y105_SLICE_X89Y105_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X59Y105_SLICE_X88Y105_A1 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_R_X59Y105_SLICE_X88Y105_A2 = CLBLM_R_X59Y105_SLICE_X88Y105_BQ;
  assign CLBLM_R_X59Y105_SLICE_X88Y105_A3 = CLBLM_L_X56Y105_SLICE_X85Y105_BQ;
  assign CLBLM_R_X59Y105_SLICE_X88Y105_A4 = CLBLL_R_X57Y108_SLICE_X87Y108_AQ;
  assign CLBLM_R_X59Y105_SLICE_X88Y105_A5 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_R_X59Y105_SLICE_X88Y105_A6 = CLBLM_L_X56Y105_SLICE_X84Y105_BQ;
  assign CLBLM_R_X59Y105_SLICE_X88Y105_AX = CLBLM_L_X62Y106_SLICE_X93Y106_CO6;
  assign CLBLM_R_X59Y105_SLICE_X88Y105_B1 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_R_X59Y105_SLICE_X88Y105_B2 = CLBLM_R_X49Y109_SLICE_X74Y109_BQ;
  assign CLBLM_R_X59Y105_SLICE_X88Y105_B3 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_R_X59Y105_SLICE_X88Y105_B4 = CLBLM_L_X62Y105_SLICE_X93Y105_BQ;
  assign CLBLM_R_X59Y105_SLICE_X88Y105_B5 = 1'b1;
  assign CLBLM_R_X59Y105_SLICE_X88Y105_B6 = CLBLM_L_X64Y108_SLICE_X97Y108_AQ;
  assign CLBLM_R_X59Y105_SLICE_X88Y105_BX = CLBLM_L_X62Y106_SLICE_X93Y106_BO6;
  assign CLBLM_R_X59Y105_SLICE_X88Y105_C1 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_R_X59Y105_SLICE_X88Y105_C2 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_R_X59Y105_SLICE_X88Y105_C3 = CLBLM_R_X59Y103_SLICE_X89Y103_DQ;
  assign CLBLM_R_X59Y105_SLICE_X88Y105_C4 = CLBLM_R_X59Y103_SLICE_X89Y103_CQ;
  assign CLBLM_R_X59Y105_SLICE_X88Y105_C5 = CLBLM_R_X59Y105_SLICE_X88Y105_BQ;
  assign CLBLM_R_X59Y105_SLICE_X88Y105_C6 = CLBLM_R_X59Y99_SLICE_X88Y99_B5Q;
  assign CLBLM_R_X59Y105_SLICE_X88Y105_CE = CLBLM_L_X60Y100_SLICE_X90Y100_CO6;
  assign CLBLM_R_X59Y105_SLICE_X88Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X59Y105_SLICE_X88Y105_D1 = 1'b1;
  assign CLBLM_R_X59Y105_SLICE_X88Y105_D2 = 1'b1;
  assign CLBLM_R_X59Y105_SLICE_X88Y105_D3 = 1'b1;
  assign CLBLM_R_X59Y105_SLICE_X88Y105_D4 = 1'b1;
  assign CLBLM_R_X59Y105_SLICE_X88Y105_D5 = 1'b1;
  assign CLBLM_R_X59Y105_SLICE_X88Y105_D6 = 1'b1;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_D = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X59Y105_SLICE_X88Y105_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign RIOI3_X105Y109_OLOGIC_X1Y110_D1 = CLBLM_R_X65Y106_SLICE_X98Y106_CQ;
  assign RIOI3_X105Y109_OLOGIC_X1Y110_T1 = 1'b1;
  assign RIOB33_X105Y111_IOB_X1Y112_O = CLBLM_R_X65Y100_SLICE_X99Y100_BQ;
  assign RIOB33_X105Y111_IOB_X1Y111_O = CLBLM_L_X64Y106_SLICE_X97Y106_DQ;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_A1 = 1'b1;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_A2 = 1'b1;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_A3 = 1'b1;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_A5 = CLBLL_R_X57Y108_SLICE_X87Y108_AQ;
  assign RIOI3_X105Y109_OLOGIC_X1Y109_D1 = CLBLM_R_X65Y100_SLICE_X99Y100_AQ;
  assign RIOI3_X105Y109_OLOGIC_X1Y109_T1 = 1'b1;
  assign CLBLM_R_X59Y106_SLICE_X89Y106_A1 = CLBLM_L_X60Y106_SLICE_X90Y106_A_XOR;
  assign CLBLM_R_X59Y106_SLICE_X89Y106_A2 = CLBLM_L_X60Y104_SLICE_X90Y104_AQ;
  assign CLBLM_R_X59Y106_SLICE_X89Y106_A3 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_R_X59Y106_SLICE_X89Y106_A4 = CLBLM_R_X59Y103_SLICE_X89Y103_CQ;
  assign CLBLM_R_X59Y106_SLICE_X89Y106_A5 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_R_X59Y106_SLICE_X89Y106_A6 = 1'b1;
  assign CLBLM_R_X59Y106_SLICE_X89Y106_B1 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X59Y106_SLICE_X89Y106_B2 = CLBLM_L_X60Y109_SLICE_X90Y109_C_XOR;
  assign CLBLM_R_X59Y106_SLICE_X89Y106_B3 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X59Y106_SLICE_X89Y106_B4 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_R_X59Y106_SLICE_X89Y106_B5 = CLBLM_R_X59Y108_SLICE_X89Y108_C_XOR;
  assign CLBLM_R_X59Y106_SLICE_X89Y106_B6 = CLBLM_L_X62Y107_SLICE_X92Y107_BO5;
  assign CLBLM_R_X59Y106_SLICE_X89Y106_C1 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X59Y106_SLICE_X89Y106_C2 = CLBLM_R_X59Y107_SLICE_X89Y107_A_XOR;
  assign CLBLM_R_X59Y106_SLICE_X89Y106_C3 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_R_X59Y106_SLICE_X89Y106_C4 = CLBLM_L_X62Y103_SLICE_X93Y103_AO6;
  assign CLBLM_R_X59Y106_SLICE_X89Y106_C5 = CLBLM_L_X60Y108_SLICE_X90Y108_A_XOR;
  assign CLBLM_R_X59Y106_SLICE_X89Y106_C6 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X59Y106_SLICE_X89Y106_CE = CLBLM_L_X60Y99_SLICE_X90Y99_DO6;
  assign CLBLM_R_X59Y106_SLICE_X89Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1 = CLBLM_R_X49Y111_SLICE_X75Y111_A5Q;
  assign CLBLM_R_X59Y106_SLICE_X89Y106_D1 = CLBLM_R_X59Y106_SLICE_X89Y106_AO6;
  assign CLBLM_R_X59Y106_SLICE_X89Y106_D2 = CLBLM_R_X59Y106_SLICE_X88Y106_CO6;
  assign CLBLM_R_X59Y106_SLICE_X89Y106_D3 = CLBLM_L_X60Y108_SLICE_X90Y108_C_XOR;
  assign CLBLM_R_X59Y106_SLICE_X89Y106_D4 = CLBLL_R_X57Y105_SLICE_X86Y105_BQ;
  assign CLBLM_R_X59Y106_SLICE_X89Y106_D5 = CLBLM_L_X62Y106_SLICE_X92Y106_AO5;
  assign CLBLM_R_X59Y106_SLICE_X89Y106_D6 = CLBLM_R_X59Y108_SLICE_X88Y108_D_XOR;
  assign CLBLM_R_X59Y106_SLICE_X89Y106_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1 = 1'b1;
  assign CLBLM_R_X59Y106_SLICE_X88Y106_A1 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_R_X59Y106_SLICE_X88Y106_A2 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X59Y106_SLICE_X88Y106_A3 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X59Y106_SLICE_X88Y106_A4 = CLBLL_R_X57Y107_SLICE_X86Y107_C_XOR;
  assign CLBLM_R_X59Y106_SLICE_X88Y106_A5 = CLBLL_R_X57Y106_SLICE_X87Y106_C_XOR;
  assign CLBLM_R_X59Y106_SLICE_X88Y106_A6 = CLBLM_L_X62Y107_SLICE_X92Y107_BO5;
  assign CLBLM_R_X59Y106_SLICE_X88Y106_B1 = CLBLL_R_X57Y105_SLICE_X87Y105_A_XOR;
  assign CLBLM_R_X59Y106_SLICE_X88Y106_B2 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X59Y106_SLICE_X88Y106_B3 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_R_X59Y106_SLICE_X88Y106_B4 = CLBLM_L_X62Y103_SLICE_X93Y103_AO6;
  assign CLBLM_R_X59Y106_SLICE_X88Y106_B5 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X59Y106_SLICE_X88Y106_B6 = CLBLL_R_X57Y106_SLICE_X86Y106_A_XOR;
  assign CLBLM_R_X59Y106_SLICE_X88Y106_C1 = CLBLM_R_X59Y104_SLICE_X88Y104_AQ;
  assign CLBLM_R_X59Y106_SLICE_X88Y106_C2 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_R_X59Y106_SLICE_X88Y106_C3 = CLBLL_R_X57Y106_SLICE_X86Y106_C_XOR;
  assign CLBLM_R_X59Y106_SLICE_X88Y106_C4 = CLBLL_R_X57Y105_SLICE_X86Y105_BQ;
  assign CLBLM_R_X59Y106_SLICE_X88Y106_C5 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_R_X59Y106_SLICE_X88Y106_C6 = CLBLL_R_X57Y109_SLICE_X87Y109_D_XOR;
  assign CLBLM_R_X59Y106_SLICE_X88Y106_CE = CLBLM_L_X60Y100_SLICE_X90Y100_BO6;
  assign CLBLM_R_X59Y106_SLICE_X88Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X59Y106_SLICE_X88Y106_D1 = CLBLL_R_X57Y106_SLICE_X87Y106_AQ;
  assign CLBLM_R_X59Y106_SLICE_X88Y106_D2 = CLBLM_R_X59Y107_SLICE_X88Y107_AQ;
  assign CLBLM_R_X59Y106_SLICE_X88Y106_D3 = CLBLM_R_X59Y99_SLICE_X89Y99_BQ;
  assign CLBLM_R_X59Y106_SLICE_X88Y106_D4 = CLBLM_R_X59Y99_SLICE_X88Y99_CQ;
  assign CLBLM_R_X59Y106_SLICE_X88Y106_D5 = CLBLM_R_X59Y99_SLICE_X88Y99_AQ;
  assign CLBLM_R_X59Y106_SLICE_X88Y106_D6 = CLBLM_R_X59Y99_SLICE_X88Y99_DQ;
  assign CLBLM_R_X59Y106_SLICE_X88Y106_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_B2 = 1'b1;
  assign RIOB33_X105Y113_IOB_X1Y114_O = CLBLM_R_X63Y103_SLICE_X95Y103_BQ;
  assign RIOB33_X105Y113_IOB_X1Y113_O = CLBLM_R_X65Y106_SLICE_X98Y106_DQ;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_B5 = CLBLM_L_X56Y98_SLICE_X85Y98_DQ;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_B6 = CLBLM_L_X50Y105_SLICE_X77Y105_AQ;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_A1 = 1'b1;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_A2 = 1'b1;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_A3 = 1'b1;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_A4 = CLBLM_R_X59Y106_SLICE_X89Y106_CQ;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_A5 = 1'b1;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_A6 = 1'b1;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_AX = CLBLM_L_X60Y100_SLICE_X90Y100_AQ;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_B1 = 1'b1;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_B2 = CLBLM_R_X49Y104_SLICE_X75Y104_DQ;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_B3 = 1'b1;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_B4 = 1'b1;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_B5 = CLBLM_R_X59Y105_SLICE_X89Y105_CQ;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_B6 = 1'b1;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_BX = CLBLM_R_X59Y105_SLICE_X89Y105_CQ;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_C1 = 1'b1;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_C2 = CLBLM_R_X59Y104_SLICE_X89Y104_CQ;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_C3 = 1'b1;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_C4 = 1'b1;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_C5 = 1'b1;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_C6 = 1'b1;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_CE = CLBLL_R_X57Y99_SLICE_X87Y99_BO6;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_CX = CLBLM_R_X59Y104_SLICE_X89Y104_CQ;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_D1 = 1'b1;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_D2 = 1'b1;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_D3 = 1'b1;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_D4 = CLBLM_L_X60Y104_SLICE_X90Y104_AQ;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_D5 = 1'b1;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_D6 = 1'b1;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_DX = CLBLM_L_X60Y104_SLICE_X90Y104_AQ;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X59Y107_SLICE_X88Y107_A1 = CLBLM_R_X59Y108_SLICE_X88Y108_B_XOR;
  assign CLBLM_R_X59Y107_SLICE_X88Y107_A2 = CLBLM_L_X62Y106_SLICE_X92Y106_AO5;
  assign CLBLM_R_X59Y107_SLICE_X88Y107_A3 = CLBLM_R_X59Y106_SLICE_X88Y106_BQ;
  assign CLBLM_R_X59Y107_SLICE_X88Y107_A4 = CLBLM_R_X59Y107_SLICE_X88Y107_BO6;
  assign CLBLM_R_X59Y107_SLICE_X88Y107_A5 = CLBLM_L_X60Y108_SLICE_X90Y108_A_XOR;
  assign CLBLM_R_X59Y107_SLICE_X88Y107_A6 = CLBLM_R_X59Y106_SLICE_X89Y106_AO6;
  assign CLBLM_R_X59Y107_SLICE_X88Y107_AX = CLBLM_R_X49Y107_SLICE_X75Y107_CQ;
  assign CLBLM_R_X59Y107_SLICE_X88Y107_B1 = CLBLL_R_X57Y109_SLICE_X87Y109_B_XOR;
  assign CLBLM_R_X59Y107_SLICE_X88Y107_B2 = CLBLL_R_X57Y106_SLICE_X86Y106_A_XOR;
  assign CLBLM_R_X59Y107_SLICE_X88Y107_B3 = CLBLM_R_X59Y103_SLICE_X88Y103_CQ;
  assign CLBLM_R_X59Y107_SLICE_X88Y107_B4 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_R_X59Y107_SLICE_X88Y107_B5 = CLBLM_R_X59Y106_SLICE_X88Y106_BQ;
  assign CLBLM_R_X59Y107_SLICE_X88Y107_B6 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_R_X59Y107_SLICE_X88Y107_C1 = CLBLM_R_X59Y106_SLICE_X88Y106_AQ;
  assign CLBLM_R_X59Y107_SLICE_X88Y107_C2 = CLBLM_R_X59Y109_SLICE_X88Y109_D_XOR;
  assign CLBLM_R_X59Y107_SLICE_X88Y107_C3 = CLBLM_L_X62Y106_SLICE_X92Y106_AO5;
  assign CLBLM_R_X59Y107_SLICE_X88Y107_C4 = CLBLM_R_X59Y106_SLICE_X89Y106_AO6;
  assign CLBLM_R_X59Y107_SLICE_X88Y107_C5 = CLBLM_R_X59Y107_SLICE_X88Y107_DO6;
  assign CLBLM_R_X59Y107_SLICE_X88Y107_C6 = CLBLM_L_X60Y109_SLICE_X90Y109_C_XOR;
  assign CLBLM_R_X59Y107_SLICE_X88Y107_CE = CLBLL_R_X57Y99_SLICE_X87Y99_BO6;
  assign CLBLM_R_X59Y107_SLICE_X88Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X59Y107_SLICE_X88Y107_D1 = CLBLL_R_X57Y107_SLICE_X86Y107_C_XOR;
  assign CLBLM_R_X59Y107_SLICE_X88Y107_D2 = CLBLM_R_X59Y106_SLICE_X88Y106_AQ;
  assign CLBLM_R_X59Y107_SLICE_X88Y107_D3 = CLBLL_R_X57Y110_SLICE_X87Y110_D_XOR;
  assign CLBLM_R_X59Y107_SLICE_X88Y107_D4 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_R_X59Y107_SLICE_X88Y107_D5 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_R_X59Y107_SLICE_X88Y107_D6 = CLBLM_R_X59Y107_SLICE_X88Y107_AQ;
  assign CLBLM_R_X59Y107_SLICE_X88Y107_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign RIOB33_X105Y115_IOB_X1Y116_O = CLBLM_R_X63Y103_SLICE_X95Y103_CQ;
  assign RIOB33_X105Y115_IOB_X1Y115_O = CLBLM_R_X63Y101_SLICE_X95Y101_AQ;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_A1 = 1'b1;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_A2 = 1'b1;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_A3 = CLBLM_R_X59Y112_SLICE_X89Y112_AQ;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_A4 = CLBLM_L_X62Y108_SLICE_X92Y108_BO6;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_A5 = 1'b1;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_A6 = 1'b1;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_AX = CLBLM_R_X59Y112_SLICE_X89Y112_AQ;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_B1 = 1'b1;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_B2 = CLBLM_R_X59Y112_SLICE_X89Y112_BQ;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_B3 = 1'b1;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_B4 = 1'b1;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_B5 = 1'b1;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_B6 = 1'b1;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_BX = CLBLM_R_X59Y112_SLICE_X89Y112_BQ;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_C1 = CLBLM_R_X59Y106_SLICE_X89Y106_BQ;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_C2 = 1'b1;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_C3 = 1'b1;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_C4 = 1'b1;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_C5 = 1'b1;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_C6 = 1'b1;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_CE = CLBLM_L_X60Y100_SLICE_X90Y100_DO6;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_CIN = CLBLM_R_X59Y107_SLICE_X89Y107_COUT;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_CX = CLBLM_R_X59Y106_SLICE_X89Y106_BQ;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_D1 = 1'b1;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_D2 = CLBLM_R_X59Y111_SLICE_X89Y111_CQ;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_D3 = 1'b1;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_D4 = 1'b1;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_D5 = 1'b1;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_D6 = 1'b1;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_DX = CLBLM_R_X59Y111_SLICE_X89Y111_CQ;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_A1 = 1'b1;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_A2 = CLBLM_R_X59Y98_SLICE_X89Y98_AQ;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_A3 = CLBLM_L_X62Y108_SLICE_X92Y108_BO6;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_A4 = 1'b1;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_A5 = CLBLM_L_X60Y100_SLICE_X90Y100_AQ;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_A6 = 1'b1;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_AX = CLBLM_L_X60Y100_SLICE_X90Y100_AQ;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_B1 = 1'b1;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_B2 = CLBLM_R_X59Y106_SLICE_X89Y106_CQ;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_B3 = 1'b1;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_B4 = 1'b1;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_B5 = 1'b1;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_B6 = CLBLM_R_X59Y98_SLICE_X89Y98_A5Q;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_BX = CLBLM_R_X59Y106_SLICE_X89Y106_CQ;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_C1 = CLBLM_R_X59Y98_SLICE_X89Y98_BQ;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_C2 = 1'b1;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_C3 = 1'b1;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_C4 = CLBLM_R_X59Y105_SLICE_X89Y105_CQ;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_C5 = 1'b1;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_C6 = 1'b1;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_CE = CLBLM_L_X60Y100_SLICE_X90Y100_CO6;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOB33_X105Y117_IOB_X1Y118_O = CLBLM_R_X65Y107_SLICE_X98Y107_AQ;
  assign RIOB33_X105Y117_IOB_X1Y117_O = CLBLM_R_X65Y107_SLICE_X98Y107_DQ;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_CX = CLBLM_R_X59Y105_SLICE_X89Y105_CQ;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_D1 = CLBLM_R_X59Y104_SLICE_X89Y104_CQ;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_D2 = 1'b1;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_D3 = 1'b1;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_D4 = 1'b1;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_D5 = 1'b1;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_D6 = CLBLM_R_X59Y98_SLICE_X89Y98_B5Q;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_DX = CLBLM_R_X59Y104_SLICE_X89Y104_CQ;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X65Y100_SLICE_X99Y100_A4 = CLBLM_L_X64Y105_SLICE_X96Y105_AQ;
  assign CLBLM_L_X56Y100_SLICE_X85Y100_C2 = 1'b1;
  assign CLBLM_L_X56Y100_SLICE_X85Y100_C5 = 1'b1;
  assign CLBLM_R_X59Y109_SLICE_X89Y109_A1 = 1'b1;
  assign CLBLM_R_X59Y109_SLICE_X89Y109_A2 = 1'b1;
  assign CLBLM_R_X59Y109_SLICE_X89Y109_A3 = 1'b1;
  assign CLBLM_R_X59Y109_SLICE_X89Y109_A4 = CLBLM_R_X59Y111_SLICE_X89Y111_AQ;
  assign CLBLM_R_X59Y109_SLICE_X89Y109_A5 = 1'b1;
  assign CLBLM_R_X59Y109_SLICE_X89Y109_A6 = 1'b1;
  assign CLBLM_L_X56Y100_SLICE_X85Y100_C6 = 1'b1;
  assign CLBLM_L_X56Y100_SLICE_X85Y100_CE = CLBLM_L_X56Y98_SLICE_X84Y98_DO6;
  assign CLBLM_R_X59Y109_SLICE_X89Y109_AX = CLBLM_R_X59Y111_SLICE_X89Y111_AQ;
  assign CLBLM_R_X59Y109_SLICE_X89Y109_B1 = 1'b1;
  assign CLBLM_R_X59Y109_SLICE_X89Y109_B2 = 1'b1;
  assign CLBLM_R_X59Y109_SLICE_X89Y109_B3 = 1'b1;
  assign CLBLM_R_X59Y109_SLICE_X89Y109_B4 = 1'b1;
  assign CLBLM_R_X59Y109_SLICE_X89Y109_B5 = 1'b1;
  assign CLBLM_R_X59Y109_SLICE_X89Y109_B6 = CLBLM_R_X59Y111_SLICE_X89Y111_BQ;
  assign CLBLM_R_X59Y109_SLICE_X89Y109_BX = CLBLM_R_X59Y111_SLICE_X89Y111_BQ;
  assign CLBLM_R_X59Y109_SLICE_X89Y109_C1 = 1'b1;
  assign CLBLM_R_X59Y109_SLICE_X89Y109_C2 = CLBLM_R_X59Y110_SLICE_X89Y110_AQ;
  assign CLBLM_R_X59Y109_SLICE_X89Y109_C3 = 1'b1;
  assign CLBLM_R_X59Y109_SLICE_X89Y109_C4 = 1'b1;
  assign CLBLM_R_X59Y109_SLICE_X89Y109_C5 = 1'b1;
  assign CLBLM_R_X59Y109_SLICE_X89Y109_C6 = 1'b1;
  assign CLBLM_R_X59Y109_SLICE_X89Y109_CIN = CLBLM_R_X59Y108_SLICE_X89Y108_COUT;
  assign CLBLM_R_X59Y109_SLICE_X89Y109_CX = 1'b0;
  assign CLBLM_R_X59Y109_SLICE_X89Y109_D1 = 1'b1;
  assign CLBLM_R_X59Y109_SLICE_X89Y109_D2 = 1'b1;
  assign CLBLM_R_X59Y109_SLICE_X89Y109_D3 = 1'b1;
  assign CLBLM_R_X59Y109_SLICE_X89Y109_D4 = 1'b1;
  assign CLBLM_R_X59Y109_SLICE_X89Y109_D5 = 1'b1;
  assign CLBLM_R_X59Y109_SLICE_X89Y109_D6 = 1'b1;
  assign CLBLM_R_X59Y109_SLICE_X89Y109_DX = 1'b0;
  assign CLBLM_R_X59Y109_SLICE_X88Y109_A1 = 1'b1;
  assign CLBLM_R_X59Y109_SLICE_X88Y109_A2 = CLBLM_R_X59Y98_SLICE_X89Y98_CQ;
  assign CLBLM_R_X59Y109_SLICE_X88Y109_A3 = 1'b1;
  assign CLBLM_R_X59Y109_SLICE_X88Y109_A4 = 1'b1;
  assign CLBLM_R_X59Y109_SLICE_X88Y109_A5 = CLBLM_L_X60Y104_SLICE_X90Y104_AQ;
  assign CLBLM_R_X59Y109_SLICE_X88Y109_A6 = 1'b1;
  assign RIOB33_X105Y119_IOB_X1Y119_O = CLBLM_R_X65Y107_SLICE_X98Y107_BQ;
  assign RIOB33_X105Y119_IOB_X1Y120_O = CLBLM_R_X65Y107_SLICE_X98Y107_CQ;
  assign CLBLM_L_X56Y100_SLICE_X85Y100_D2 = 1'b1;
  assign CLBLM_R_X59Y109_SLICE_X88Y109_AX = CLBLM_L_X60Y104_SLICE_X90Y104_AQ;
  assign CLBLM_R_X59Y109_SLICE_X88Y109_B1 = 1'b1;
  assign CLBLM_R_X59Y109_SLICE_X88Y109_B2 = 1'b1;
  assign CLBLM_R_X59Y109_SLICE_X88Y109_B3 = CLBLM_R_X59Y98_SLICE_X89Y98_C5Q;
  assign CLBLM_L_X56Y100_SLICE_X85Y100_D3 = 1'b1;
  assign CLBLM_R_X59Y109_SLICE_X88Y109_B4 = 1'b1;
  assign CLBLM_R_X59Y109_SLICE_X88Y109_B5 = CLBLM_R_X59Y112_SLICE_X89Y112_AQ;
  assign CLBLM_R_X59Y109_SLICE_X88Y109_B6 = 1'b1;
  assign CLBLM_L_X56Y100_SLICE_X85Y100_D4 = 1'b1;
  assign CLBLM_R_X59Y109_SLICE_X88Y109_BX = CLBLM_R_X59Y112_SLICE_X89Y112_AQ;
  assign CLBLM_R_X59Y109_SLICE_X88Y109_C1 = 1'b1;
  assign CLBLM_R_X59Y109_SLICE_X88Y109_C2 = 1'b1;
  assign CLBLM_R_X59Y109_SLICE_X88Y109_C3 = CLBLM_R_X59Y96_SLICE_X89Y96_AQ;
  assign CLBLM_R_X59Y109_SLICE_X88Y109_C4 = 1'b1;
  assign CLBLM_R_X59Y109_SLICE_X88Y109_C5 = 1'b1;
  assign CLBLM_R_X59Y109_SLICE_X88Y109_C6 = CLBLM_R_X59Y112_SLICE_X89Y112_BQ;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_T1 = 1'b1;
  assign CLBLM_R_X59Y109_SLICE_X88Y109_CIN = CLBLM_R_X59Y108_SLICE_X88Y108_COUT;
  assign CLBLM_R_X59Y109_SLICE_X88Y109_CX = CLBLM_R_X59Y112_SLICE_X89Y112_BQ;
  assign CLBLM_R_X59Y109_SLICE_X88Y109_D1 = CLBLM_R_X59Y106_SLICE_X89Y106_BQ;
  assign CLBLM_R_X59Y109_SLICE_X88Y109_D2 = 1'b1;
  assign CLBLM_R_X59Y109_SLICE_X88Y109_D3 = CLBLM_R_X59Y96_SLICE_X89Y96_A5Q;
  assign CLBLM_R_X59Y109_SLICE_X88Y109_D4 = 1'b1;
  assign CLBLM_R_X59Y109_SLICE_X88Y109_D5 = 1'b1;
  assign CLBLM_L_X56Y100_SLICE_X85Y100_DX = CLBLM_L_X56Y97_SLICE_X84Y97_AO6;
  assign CLBLM_R_X59Y109_SLICE_X88Y109_D6 = 1'b1;
  assign CLBLM_R_X59Y109_SLICE_X88Y109_DX = CLBLM_R_X59Y106_SLICE_X89Y106_BQ;
  assign CLBLM_L_X56Y100_SLICE_X84Y100_A1 = CLBLM_L_X56Y102_SLICE_X85Y102_A5Q;
  assign CLBLM_L_X56Y100_SLICE_X84Y100_A2 = 1'b1;
  assign CLBLM_L_X56Y100_SLICE_X84Y100_A3 = CLBLM_L_X56Y100_SLICE_X84Y100_AQ;
  assign CLBLM_L_X56Y100_SLICE_X84Y100_A4 = 1'b1;
  assign CLBLM_L_X56Y100_SLICE_X84Y100_A5 = CLBLM_L_X56Y102_SLICE_X85Y102_AQ;
  assign CLBLM_L_X56Y100_SLICE_X84Y100_A6 = 1'b1;
  assign CLBLM_L_X56Y100_SLICE_X84Y100_B1 = CLBLM_L_X56Y102_SLICE_X85Y102_A5Q;
  assign CLBLM_L_X56Y100_SLICE_X84Y100_B2 = CLBLM_L_X56Y100_SLICE_X84Y100_BQ;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_D1 = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X56Y100_SLICE_X84Y100_B4 = 1'b1;
  assign CLBLM_L_X56Y100_SLICE_X84Y100_B5 = 1'b1;
  assign CLBLM_L_X56Y100_SLICE_X84Y100_B6 = 1'b1;
  assign CLBLM_R_X59Y110_SLICE_X89Y110_A1 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X59Y110_SLICE_X89Y110_A2 = CLBLM_L_X60Y110_SLICE_X90Y110_C_XOR;
  assign CLBLM_R_X59Y110_SLICE_X89Y110_A3 = CLBLM_R_X59Y109_SLICE_X89Y109_C_XOR;
  assign CLBLM_R_X59Y110_SLICE_X89Y110_A4 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_R_X59Y110_SLICE_X89Y110_A5 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X59Y110_SLICE_X89Y110_A6 = CLBLM_L_X62Y100_SLICE_X93Y100_BO6;
  assign CLBLM_R_X59Y110_SLICE_X89Y110_B1 = CLBLM_R_X59Y106_SLICE_X89Y106_AO6;
  assign CLBLM_R_X59Y110_SLICE_X89Y110_B2 = CLBLM_L_X62Y106_SLICE_X92Y106_AO5;
  assign CLBLM_R_X59Y110_SLICE_X89Y110_B3 = CLBLM_R_X59Y110_SLICE_X88Y110_C_XOR;
  assign CLBLM_R_X59Y110_SLICE_X89Y110_B4 = CLBLL_R_X57Y109_SLICE_X86Y109_DO6;
  assign CLBLM_R_X59Y110_SLICE_X89Y110_B5 = CLBLL_R_X57Y109_SLICE_X86Y109_BQ;
  assign CLBLM_R_X59Y110_SLICE_X89Y110_B6 = CLBLM_L_X60Y110_SLICE_X90Y110_B_XOR;
  assign RIOB33_X105Y121_IOB_X1Y122_O = CLBLM_L_X64Y106_SLICE_X97Y106_AQ;
  assign CLBLM_R_X59Y110_SLICE_X89Y110_C1 = CLBLL_R_X57Y108_SLICE_X87Y108_AQ;
  assign CLBLM_R_X59Y110_SLICE_X89Y110_C2 = CLBLM_L_X60Y109_SLICE_X90Y109_A_XOR;
  assign CLBLM_R_X59Y110_SLICE_X89Y110_C3 = CLBLM_R_X59Y106_SLICE_X89Y106_AO6;
  assign CLBLM_R_X59Y110_SLICE_X89Y110_C4 = CLBLM_L_X62Y106_SLICE_X92Y106_AO5;
  assign CLBLM_R_X59Y110_SLICE_X89Y110_C5 = CLBLM_R_X59Y109_SLICE_X88Y109_B_XOR;
  assign CLBLM_R_X59Y110_SLICE_X89Y110_C6 = CLBLM_R_X59Y110_SLICE_X89Y110_DO6;
  assign CLBLM_R_X59Y110_SLICE_X89Y110_CE = CLBLM_L_X60Y100_SLICE_X90Y100_DO6;
  assign RIOB33_X105Y121_IOB_X1Y121_O = CLBLM_R_X65Y106_SLICE_X98Y106_AQ;
  assign CLBLM_R_X59Y110_SLICE_X89Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X59Y110_SLICE_X89Y110_D1 = CLBLL_R_X57Y108_SLICE_X87Y108_AQ;
  assign CLBLM_R_X59Y110_SLICE_X89Y110_D2 = CLBLL_R_X57Y107_SLICE_X86Y107_A_XOR;
  assign CLBLM_R_X59Y110_SLICE_X89Y110_D3 = CLBLL_R_X57Y110_SLICE_X87Y110_B_XOR;
  assign CLBLM_R_X59Y110_SLICE_X89Y110_D4 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_R_X59Y110_SLICE_X89Y110_D5 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_R_X59Y110_SLICE_X89Y110_D6 = CLBLM_R_X59Y104_SLICE_X88Y104_BQ;
  assign CLBLM_R_X59Y110_SLICE_X89Y110_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X59Y110_SLICE_X88Y110_A1 = 1'b1;
  assign CLBLM_R_X59Y110_SLICE_X88Y110_A2 = 1'b1;
  assign CLBLM_R_X59Y110_SLICE_X88Y110_A3 = 1'b1;
  assign CLBLM_R_X59Y110_SLICE_X88Y110_A4 = 1'b1;
  assign CLBLM_R_X59Y110_SLICE_X88Y110_A5 = 1'b1;
  assign CLBLM_R_X59Y110_SLICE_X88Y110_A6 = CLBLM_R_X59Y111_SLICE_X89Y111_CQ;
  assign CLBLM_R_X59Y110_SLICE_X88Y110_AX = 1'b0;
  assign CLBLM_R_X59Y110_SLICE_X88Y110_B1 = 1'b1;
  assign CLBLM_R_X59Y110_SLICE_X88Y110_B2 = 1'b1;
  assign CLBLM_R_X59Y110_SLICE_X88Y110_B3 = 1'b1;
  assign CLBLM_R_X59Y110_SLICE_X88Y110_B4 = 1'b1;
  assign CLBLM_R_X59Y110_SLICE_X88Y110_B5 = 1'b1;
  assign CLBLM_R_X59Y110_SLICE_X88Y110_B6 = CLBLM_R_X59Y111_SLICE_X89Y111_AQ;
  assign CLBLM_R_X59Y110_SLICE_X88Y110_BX = 1'b0;
  assign CLBLM_R_X59Y110_SLICE_X88Y110_C1 = 1'b1;
  assign CLBLM_R_X59Y110_SLICE_X88Y110_C2 = 1'b1;
  assign CLBLM_R_X59Y110_SLICE_X88Y110_C3 = 1'b1;
  assign CLBLM_R_X59Y110_SLICE_X88Y110_C4 = 1'b1;
  assign CLBLM_R_X59Y110_SLICE_X88Y110_C5 = 1'b1;
  assign CLBLM_R_X59Y110_SLICE_X88Y110_C6 = CLBLM_R_X59Y111_SLICE_X89Y111_BQ;
  assign CLBLM_R_X59Y110_SLICE_X88Y110_CIN = CLBLM_R_X59Y109_SLICE_X88Y109_COUT;
  assign CLBLM_R_X59Y110_SLICE_X88Y110_CX = 1'b0;
  assign CLBLM_R_X59Y110_SLICE_X88Y110_D1 = 1'b1;
  assign CLBLM_R_X59Y110_SLICE_X88Y110_D2 = 1'b1;
  assign CLBLM_R_X59Y110_SLICE_X88Y110_D3 = 1'b1;
  assign CLBLM_R_X59Y110_SLICE_X88Y110_D4 = 1'b1;
  assign CLBLM_R_X59Y110_SLICE_X88Y110_D5 = 1'b1;
  assign CLBLM_R_X59Y110_SLICE_X88Y110_D6 = CLBLM_R_X59Y110_SLICE_X89Y110_AQ;
  assign CLBLM_R_X59Y110_SLICE_X88Y110_DX = 1'b0;
  assign RIOB33_X105Y123_IOB_X1Y124_O = CLBLM_R_X65Y106_SLICE_X98Y106_BQ;
  assign RIOB33_X105Y123_IOB_X1Y123_O = CLBLM_R_X63Y103_SLICE_X95Y103_AQ;
  assign CLBLM_R_X59Y111_SLICE_X89Y111_A1 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X59Y111_SLICE_X89Y111_A2 = CLBLM_L_X60Y110_SLICE_X90Y110_A_XOR;
  assign CLBLM_R_X59Y111_SLICE_X89Y111_A3 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_R_X59Y111_SLICE_X89Y111_A4 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X59Y111_SLICE_X89Y111_A5 = CLBLM_L_X62Y97_SLICE_X92Y97_BO6;
  assign CLBLM_R_X59Y111_SLICE_X89Y111_A6 = CLBLM_R_X59Y109_SLICE_X89Y109_A_XOR;
  assign CLBLM_R_X59Y111_SLICE_X89Y111_B1 = CLBLM_R_X59Y109_SLICE_X89Y109_B_XOR;
  assign CLBLM_R_X59Y111_SLICE_X89Y111_B2 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X59Y111_SLICE_X89Y111_B3 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_R_X59Y111_SLICE_X89Y111_B4 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X59Y111_SLICE_X89Y111_B5 = CLBLM_L_X62Y100_SLICE_X93Y100_AO6;
  assign CLBLM_R_X59Y111_SLICE_X89Y111_B6 = CLBLM_L_X60Y110_SLICE_X90Y110_B_XOR;
  assign CLBLM_R_X59Y111_SLICE_X89Y111_C1 = CLBLM_R_X59Y108_SLICE_X89Y108_D_XOR;
  assign CLBLM_R_X59Y111_SLICE_X89Y111_C2 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_R_X59Y111_SLICE_X89Y111_C3 = CLBLM_L_X62Y97_SLICE_X92Y97_AO6;
  assign CLBLM_R_X59Y111_SLICE_X89Y111_C4 = CLBLM_L_X60Y109_SLICE_X90Y109_D_XOR;
  assign CLBLM_R_X59Y111_SLICE_X89Y111_C5 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X59Y111_SLICE_X89Y111_C6 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X59Y111_SLICE_X89Y111_CE = CLBLM_L_X60Y100_SLICE_X90Y100_DO6;
  assign CLBLM_R_X59Y111_SLICE_X89Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X59Y111_SLICE_X89Y111_D1 = CLBLM_L_X60Y110_SLICE_X90Y110_C_XOR;
  assign CLBLM_R_X59Y111_SLICE_X89Y111_D2 = CLBLM_R_X59Y111_SLICE_X88Y111_AO6;
  assign CLBLM_R_X59Y111_SLICE_X89Y111_D3 = CLBLL_R_X57Y109_SLICE_X86Y109_CQ;
  assign CLBLM_R_X59Y111_SLICE_X89Y111_D4 = CLBLM_L_X62Y106_SLICE_X92Y106_AO5;
  assign CLBLM_R_X59Y111_SLICE_X89Y111_D5 = CLBLM_R_X59Y106_SLICE_X89Y106_AO6;
  assign CLBLM_R_X59Y111_SLICE_X89Y111_D6 = CLBLM_R_X59Y110_SLICE_X88Y110_D_XOR;
  assign CLBLM_R_X59Y111_SLICE_X89Y111_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X59Y111_SLICE_X88Y111_A1 = CLBLL_R_X57Y111_SLICE_X87Y111_D_XOR;
  assign CLBLM_R_X59Y111_SLICE_X88Y111_A2 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_R_X59Y111_SLICE_X88Y111_A3 = CLBLL_R_X57Y108_SLICE_X86Y108_C_XOR;
  assign CLBLM_R_X59Y111_SLICE_X88Y111_A4 = CLBLL_R_X57Y109_SLICE_X86Y109_CQ;
  assign CLBLM_R_X59Y111_SLICE_X88Y111_A5 = CLBLM_R_X59Y99_SLICE_X88Y99_AQ;
  assign CLBLM_R_X59Y111_SLICE_X88Y111_A6 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_R_X59Y111_SLICE_X88Y111_B1 = CLBLM_R_X59Y99_SLICE_X88Y99_CQ;
  assign CLBLM_R_X59Y111_SLICE_X88Y111_B2 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_R_X59Y111_SLICE_X88Y111_B3 = CLBLL_R_X57Y107_SLICE_X86Y107_D_XOR;
  assign CLBLM_R_X59Y111_SLICE_X88Y111_B4 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_R_X59Y111_SLICE_X88Y111_B5 = CLBLM_L_X60Y108_SLICE_X91Y108_AQ;
  assign CLBLM_R_X59Y111_SLICE_X88Y111_B6 = CLBLL_R_X57Y111_SLICE_X87Y111_A_XOR;
  assign CLBLM_R_X59Y111_SLICE_X88Y111_C1 = CLBLL_R_X57Y109_SLICE_X86Y109_AQ;
  assign CLBLM_R_X59Y111_SLICE_X88Y111_C2 = CLBLM_L_X62Y106_SLICE_X92Y106_AO5;
  assign CLBLM_R_X59Y111_SLICE_X88Y111_C3 = CLBLM_R_X59Y110_SLICE_X88Y110_B_XOR;
  assign CLBLM_R_X59Y111_SLICE_X88Y111_C4 = CLBLM_R_X59Y106_SLICE_X89Y106_AO6;
  assign CLBLM_R_X59Y111_SLICE_X88Y111_C5 = CLBLM_R_X59Y111_SLICE_X88Y111_DO6;
  assign CLBLM_R_X59Y111_SLICE_X88Y111_C6 = CLBLM_L_X60Y110_SLICE_X90Y110_A_XOR;
  assign CLBLM_R_X59Y111_SLICE_X88Y111_D1 = CLBLL_R_X57Y109_SLICE_X86Y109_AQ;
  assign CLBLM_R_X59Y111_SLICE_X88Y111_D2 = CLBLM_R_X59Y99_SLICE_X88Y99_DQ;
  assign CLBLM_R_X59Y111_SLICE_X88Y111_D3 = CLBLL_R_X57Y111_SLICE_X87Y111_B_XOR;
  assign CLBLM_R_X59Y111_SLICE_X88Y111_D4 = CLBLL_R_X57Y108_SLICE_X86Y108_A_XOR;
  assign CLBLM_R_X59Y111_SLICE_X88Y111_D5 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_R_X59Y111_SLICE_X88Y111_D6 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign RIOB33_X105Y125_IOB_X1Y126_O = CLBLM_L_X64Y106_SLICE_X97Y106_CQ;
  assign RIOB33_X105Y125_IOB_X1Y125_O = CLBLM_L_X64Y106_SLICE_X97Y106_BQ;
  assign CLBLM_R_X59Y112_SLICE_X89Y112_A1 = CLBLM_L_X62Y106_SLICE_X93Y106_BO5;
  assign CLBLM_R_X59Y112_SLICE_X89Y112_A2 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_R_X59Y112_SLICE_X89Y112_A3 = CLBLM_L_X60Y109_SLICE_X90Y109_A_XOR;
  assign CLBLM_R_X59Y112_SLICE_X89Y112_A4 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X59Y112_SLICE_X89Y112_A5 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X59Y112_SLICE_X89Y112_A6 = CLBLM_R_X59Y108_SLICE_X89Y108_A_XOR;
  assign CLBLM_R_X59Y112_SLICE_X89Y112_B1 = CLBLM_L_X60Y109_SLICE_X90Y109_B_XOR;
  assign CLBLM_R_X59Y112_SLICE_X89Y112_B2 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_R_X59Y112_SLICE_X89Y112_B3 = CLBLM_L_X62Y108_SLICE_X92Y108_BO5;
  assign CLBLM_R_X59Y112_SLICE_X89Y112_B4 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X59Y112_SLICE_X89Y112_B5 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X59Y112_SLICE_X89Y112_B6 = CLBLM_R_X59Y108_SLICE_X89Y108_B_XOR;
  assign CLBLM_R_X59Y112_SLICE_X89Y112_C1 = CLBLM_R_X59Y109_SLICE_X88Y109_C_XOR;
  assign CLBLM_R_X59Y112_SLICE_X89Y112_C2 = CLBLM_L_X62Y106_SLICE_X92Y106_AO5;
  assign CLBLM_R_X59Y112_SLICE_X89Y112_C3 = CLBLL_R_X57Y108_SLICE_X87Y108_DO6;
  assign CLBLM_R_X59Y112_SLICE_X89Y112_C4 = CLBLM_R_X59Y106_SLICE_X89Y106_AO6;
  assign CLBLM_R_X59Y112_SLICE_X89Y112_C5 = CLBLM_L_X60Y109_SLICE_X90Y109_B_XOR;
  assign CLBLM_R_X59Y112_SLICE_X89Y112_C6 = CLBLL_R_X57Y108_SLICE_X87Y108_BQ;
  assign CLBLM_R_X59Y112_SLICE_X89Y112_CE = CLBLM_L_X60Y99_SLICE_X90Y99_DO6;
  assign CLBLM_R_X59Y112_SLICE_X89Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X59Y112_SLICE_X89Y112_D1 = 1'b1;
  assign CLBLM_R_X59Y112_SLICE_X89Y112_D2 = 1'b1;
  assign CLBLM_R_X59Y112_SLICE_X89Y112_D3 = 1'b1;
  assign CLBLM_R_X59Y112_SLICE_X89Y112_D4 = 1'b1;
  assign CLBLM_R_X59Y112_SLICE_X89Y112_D5 = 1'b1;
  assign CLBLM_R_X59Y112_SLICE_X89Y112_D6 = 1'b1;
  assign CLBLM_R_X59Y112_SLICE_X89Y112_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X59Y112_SLICE_X88Y112_A1 = 1'b1;
  assign CLBLM_R_X59Y112_SLICE_X88Y112_A2 = 1'b1;
  assign CLBLM_R_X59Y112_SLICE_X88Y112_A3 = 1'b1;
  assign CLBLM_R_X59Y112_SLICE_X88Y112_A4 = 1'b1;
  assign CLBLM_R_X59Y112_SLICE_X88Y112_A5 = 1'b1;
  assign CLBLM_R_X59Y112_SLICE_X88Y112_A6 = 1'b1;
  assign CLBLM_R_X59Y112_SLICE_X88Y112_B1 = 1'b1;
  assign CLBLM_R_X59Y112_SLICE_X88Y112_B2 = 1'b1;
  assign CLBLM_R_X59Y112_SLICE_X88Y112_B3 = 1'b1;
  assign CLBLM_R_X59Y112_SLICE_X88Y112_B4 = 1'b1;
  assign CLBLM_R_X59Y112_SLICE_X88Y112_B5 = 1'b1;
  assign CLBLM_R_X59Y112_SLICE_X88Y112_B6 = 1'b1;
  assign CLBLM_R_X59Y112_SLICE_X88Y112_C1 = 1'b1;
  assign CLBLM_R_X59Y112_SLICE_X88Y112_C2 = 1'b1;
  assign CLBLM_R_X59Y112_SLICE_X88Y112_C3 = 1'b1;
  assign CLBLM_R_X59Y112_SLICE_X88Y112_C4 = 1'b1;
  assign CLBLM_R_X59Y112_SLICE_X88Y112_C5 = 1'b1;
  assign CLBLM_R_X59Y112_SLICE_X88Y112_C6 = 1'b1;
  assign CLBLM_R_X59Y112_SLICE_X88Y112_D1 = 1'b1;
  assign CLBLM_R_X59Y112_SLICE_X88Y112_D2 = 1'b1;
  assign CLBLM_R_X59Y112_SLICE_X88Y112_D3 = 1'b1;
  assign CLBLM_R_X59Y112_SLICE_X88Y112_D4 = 1'b1;
  assign CLBLM_R_X59Y112_SLICE_X88Y112_D5 = 1'b1;
  assign CLBLM_R_X59Y112_SLICE_X88Y112_D6 = 1'b1;
  assign RIOB33_X105Y127_IOB_X1Y127_O = CLBLM_R_X59Y102_SLICE_X88Y102_AQ;
  assign RIOB33_X105Y129_IOB_X1Y130_O = CLBLM_L_X62Y103_SLICE_X92Y103_AQ;
  assign RIOB33_X105Y129_IOB_X1Y129_O = CLBLM_L_X62Y104_SLICE_X93Y104_AQ;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_C6 = 1'b1;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_CE = CLBLM_L_X60Y98_SLICE_X91Y98_BQ;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X65Y101_SLICE_X99Y101_D1 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_L_X56Y101_SLICE_X85Y101_CE = CLBLL_R_X57Y100_SLICE_X87Y100_DO6;
  assign CLBLM_L_X56Y101_SLICE_X85Y101_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X56Y101_SLICE_X85Y101_D3 = CLBLM_L_X56Y99_SLICE_X85Y99_BQ;
  assign CLBLM_L_X56Y101_SLICE_X84Y101_A6 = 1'b1;
  assign RIOB33_X105Y131_IOB_X1Y132_O = CLBLM_L_X60Y110_SLICE_X91Y110_AQ;
  assign RIOB33_X105Y131_IOB_X1Y131_O = CLBLM_R_X59Y102_SLICE_X89Y102_AQ;
  assign CLBLM_L_X56Y101_SLICE_X84Y101_B1 = CLBLM_L_X56Y102_SLICE_X85Y102_A5Q;
  assign CLBLM_L_X56Y101_SLICE_X84Y101_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign RIOB33_X105Y133_IOB_X1Y134_O = CLBLM_L_X62Y110_SLICE_X92Y110_AQ;
  assign RIOB33_X105Y133_IOB_X1Y133_O = CLBLM_L_X62Y106_SLICE_X93Y106_AQ;
  assign CLBLM_L_X60Y96_SLICE_X91Y96_D5 = 1'b1;
  assign CLBLM_L_X60Y96_SLICE_X91Y96_D6 = 1'b1;
  assign CLBLM_L_X60Y96_SLICE_X90Y96_A1 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X75Y104_A1 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X75Y104_A2 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X49Y104_SLICE_X75Y104_A3 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X49Y104_SLICE_X75Y104_A4 = CLBLM_R_X49Y119_SLICE_X74Y119_BQ;
  assign CLBLM_R_X49Y104_SLICE_X75Y104_A5 = CLBLM_R_X49Y119_SLICE_X74Y119_AQ;
  assign CLBLM_R_X49Y104_SLICE_X75Y104_A6 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X75Y104_AX = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X49Y104_SLICE_X75Y104_B1 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X75Y104_B2 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X75Y104_B3 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X75Y104_B4 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X75Y104_B5 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X75Y104_B6 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X75Y104_BX = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X49Y104_SLICE_X75Y104_C1 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X75Y104_C2 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X75Y104_C3 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X75Y104_C4 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X75Y104_C5 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X75Y104_C6 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X75Y104_CE = CLBLM_R_X49Y104_SLICE_X75Y104_AO6;
  assign CLBLM_R_X49Y104_SLICE_X75Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X49Y104_SLICE_X75Y104_CX = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X49Y104_SLICE_X75Y104_D1 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X75Y104_D2 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X75Y104_D3 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X75Y104_D4 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X75Y104_D5 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X75Y104_D6 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X75Y104_DX = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X49Y104_SLICE_X75Y104_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X49Y104_SLICE_X74Y104_A1 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X74Y104_A2 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X74Y104_A3 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X74Y104_A4 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X74Y104_A5 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X74Y104_A6 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X74Y104_AX = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X49Y104_SLICE_X74Y104_B1 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X74Y104_B2 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X74Y104_B3 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X74Y104_B4 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X74Y104_B5 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X74Y104_B6 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X74Y104_BX = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X49Y104_SLICE_X74Y104_C1 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X74Y104_C2 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X74Y104_C3 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X74Y104_C4 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X74Y104_C5 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X74Y104_C6 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X74Y104_CE = CLBLM_R_X49Y104_SLICE_X75Y104_AO6;
  assign CLBLM_R_X49Y104_SLICE_X74Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X49Y104_SLICE_X74Y104_D1 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X74Y104_D2 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X74Y104_D3 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X74Y104_D4 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X74Y104_D5 = 1'b1;
  assign CLBLM_R_X49Y104_SLICE_X74Y104_D6 = 1'b1;
  assign RIOB33_X105Y135_IOB_X1Y136_O = CLBLM_L_X60Y111_SLICE_X91Y111_BQ;
  assign RIOB33_X105Y135_IOB_X1Y135_O = CLBLM_L_X62Y108_SLICE_X93Y108_AQ;
  assign CLBLM_R_X49Y104_SLICE_X74Y104_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X49Y105_SLICE_X75Y105_A1 = CLBLM_L_X56Y101_SLICE_X85Y101_CQ;
  assign CLBLM_R_X49Y105_SLICE_X75Y105_A2 = CLBLM_L_X50Y106_SLICE_X77Y106_AO5;
  assign CLBLM_R_X49Y105_SLICE_X75Y105_A3 = CLBLM_L_X56Y101_SLICE_X85Y101_AQ;
  assign CLBLM_R_X49Y105_SLICE_X75Y105_A4 = CLBLL_R_X57Y100_SLICE_X86Y100_CQ;
  assign CLBLM_R_X49Y105_SLICE_X75Y105_A5 = 1'b1;
  assign CLBLM_R_X49Y105_SLICE_X75Y105_A6 = CLBLL_R_X57Y100_SLICE_X86Y100_DQ;
  assign CLBLM_R_X49Y105_SLICE_X75Y105_AX = CLBLM_R_X49Y106_SLICE_X74Y106_CO6;
  assign CLBLM_R_X49Y105_SLICE_X75Y105_B1 = CLBLM_L_X56Y101_SLICE_X85Y101_CQ;
  assign CLBLM_R_X49Y105_SLICE_X75Y105_B2 = CLBLM_L_X50Y106_SLICE_X77Y106_AO5;
  assign CLBLM_R_X49Y105_SLICE_X75Y105_B3 = CLBLM_L_X56Y101_SLICE_X85Y101_AQ;
  assign CLBLM_R_X49Y105_SLICE_X75Y105_B4 = CLBLL_R_X57Y100_SLICE_X86Y100_CQ;
  assign CLBLM_R_X49Y105_SLICE_X75Y105_B5 = CLBLL_L_X54Y100_SLICE_X82Y100_BQ;
  assign CLBLM_R_X49Y105_SLICE_X75Y105_B6 = CLBLL_R_X57Y100_SLICE_X87Y100_CQ;
  assign CLBLM_R_X49Y105_SLICE_X75Y105_C1 = CLBLM_R_X49Y105_SLICE_X75Y105_F7AMUX_O;
  assign CLBLM_R_X49Y105_SLICE_X75Y105_C2 = CLBLM_R_X49Y107_SLICE_X75Y107_F7AMUX_O;
  assign CLBLM_R_X49Y105_SLICE_X75Y105_C3 = CLBLM_R_X53Y100_SLICE_X81Y100_AQ;
  assign CLBLM_R_X49Y105_SLICE_X75Y105_C4 = 1'b1;
  assign CLBLM_R_X49Y105_SLICE_X75Y105_C5 = 1'b1;
  assign CLBLM_R_X49Y105_SLICE_X75Y105_C6 = 1'b1;
  assign CLBLM_R_X49Y105_SLICE_X75Y105_CE = CLBLM_L_X56Y98_SLICE_X84Y98_DO6;
  assign CLBLM_R_X49Y105_SLICE_X75Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X49Y105_SLICE_X75Y105_D1 = 1'b1;
  assign CLBLM_R_X49Y105_SLICE_X75Y105_D2 = 1'b1;
  assign CLBLM_R_X49Y105_SLICE_X75Y105_D3 = 1'b1;
  assign CLBLM_R_X49Y105_SLICE_X75Y105_D4 = 1'b1;
  assign CLBLM_R_X49Y105_SLICE_X75Y105_D5 = 1'b1;
  assign CLBLM_R_X49Y105_SLICE_X75Y105_D6 = 1'b1;
  assign CLBLM_R_X49Y105_SLICE_X75Y105_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X49Y105_SLICE_X74Y105_A1 = 1'b1;
  assign CLBLM_R_X49Y105_SLICE_X74Y105_A2 = 1'b1;
  assign CLBLM_R_X49Y105_SLICE_X74Y105_A3 = 1'b1;
  assign CLBLM_R_X49Y105_SLICE_X74Y105_A4 = 1'b1;
  assign CLBLM_R_X49Y105_SLICE_X74Y105_A5 = 1'b1;
  assign CLBLM_R_X49Y105_SLICE_X74Y105_A6 = 1'b1;
  assign CLBLM_R_X49Y105_SLICE_X74Y105_B1 = 1'b1;
  assign CLBLM_R_X49Y105_SLICE_X74Y105_B2 = 1'b1;
  assign CLBLM_R_X49Y105_SLICE_X74Y105_B3 = 1'b1;
  assign CLBLM_R_X49Y105_SLICE_X74Y105_B4 = 1'b1;
  assign CLBLM_R_X49Y105_SLICE_X74Y105_B5 = 1'b1;
  assign CLBLM_R_X49Y105_SLICE_X74Y105_B6 = 1'b1;
  assign RIOB33_X105Y137_IOB_X1Y137_O = CLBLM_L_X60Y111_SLICE_X90Y111_AQ;
  assign RIOB33_X105Y137_IOB_X1Y138_O = CLBLM_L_X62Y110_SLICE_X92Y110_BQ;
  assign CLBLM_R_X49Y105_SLICE_X74Y105_C1 = 1'b1;
  assign CLBLM_R_X49Y105_SLICE_X74Y105_C2 = 1'b1;
  assign CLBLM_R_X49Y105_SLICE_X74Y105_C3 = 1'b1;
  assign CLBLM_R_X49Y105_SLICE_X74Y105_C4 = 1'b1;
  assign CLBLM_R_X49Y105_SLICE_X74Y105_C5 = 1'b1;
  assign CLBLM_R_X49Y105_SLICE_X74Y105_C6 = 1'b1;
  assign CLBLM_R_X49Y105_SLICE_X74Y105_D1 = 1'b1;
  assign CLBLM_R_X49Y105_SLICE_X74Y105_D2 = 1'b1;
  assign CLBLM_R_X49Y105_SLICE_X74Y105_D3 = 1'b1;
  assign CLBLM_R_X49Y105_SLICE_X74Y105_D4 = 1'b1;
  assign CLBLM_R_X49Y105_SLICE_X74Y105_D5 = 1'b1;
  assign CLBLM_R_X49Y105_SLICE_X74Y105_D6 = 1'b1;
  assign CLBLM_R_X49Y106_SLICE_X75Y106_A1 = CLBLM_L_X50Y106_SLICE_X77Y106_AO5;
  assign CLBLM_R_X49Y106_SLICE_X75Y106_A2 = CLBLL_R_X57Y100_SLICE_X87Y100_AQ;
  assign CLBLM_R_X49Y106_SLICE_X75Y106_A3 = CLBLM_L_X56Y101_SLICE_X85Y101_CQ;
  assign CLBLM_R_X49Y106_SLICE_X75Y106_A4 = CLBLL_R_X57Y100_SLICE_X86Y100_DQ;
  assign CLBLM_R_X49Y106_SLICE_X75Y106_A5 = CLBLL_R_X57Y100_SLICE_X86Y100_CQ;
  assign CLBLM_R_X49Y106_SLICE_X75Y106_A6 = CLBLL_R_X57Y100_SLICE_X87Y100_CQ;
  assign CLBLM_R_X49Y106_SLICE_X75Y106_AX = CLBLM_R_X49Y106_SLICE_X74Y106_CO6;
  assign CLBLM_R_X49Y106_SLICE_X75Y106_B1 = CLBLM_L_X50Y106_SLICE_X77Y106_AO5;
  assign CLBLM_R_X49Y106_SLICE_X75Y106_B2 = CLBLL_R_X57Y100_SLICE_X87Y100_AQ;
  assign CLBLM_R_X49Y106_SLICE_X75Y106_B3 = CLBLM_L_X56Y101_SLICE_X85Y101_CQ;
  assign CLBLM_R_X49Y106_SLICE_X75Y106_B4 = CLBLL_R_X57Y101_SLICE_X87Y101_CQ;
  assign CLBLM_R_X49Y106_SLICE_X75Y106_B5 = CLBLL_R_X57Y100_SLICE_X87Y100_CQ;
  assign CLBLM_R_X49Y106_SLICE_X75Y106_B6 = CLBLL_L_X54Y100_SLICE_X82Y100_BQ;
  assign CLBLM_R_X49Y106_SLICE_X75Y106_BX = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X49Y106_SLICE_X75Y106_C1 = CLBLM_L_X50Y105_SLICE_X76Y105_BO6;
  assign CLBLM_R_X49Y106_SLICE_X75Y106_C2 = CLBLM_R_X49Y106_SLICE_X74Y106_CO6;
  assign CLBLM_R_X49Y106_SLICE_X75Y106_C3 = CLBLL_R_X57Y100_SLICE_X87Y100_BQ;
  assign CLBLM_R_X49Y106_SLICE_X75Y106_C4 = CLBLL_R_X57Y101_SLICE_X87Y101_DQ;
  assign CLBLM_R_X49Y106_SLICE_X75Y106_C5 = CLBLM_L_X50Y106_SLICE_X77Y106_AO5;
  assign CLBLM_R_X49Y106_SLICE_X75Y106_C6 = CLBLM_R_X49Y106_SLICE_X75Y106_DO6;
  assign CLBLM_R_X49Y106_SLICE_X75Y106_CE = CLBLM_R_X49Y104_SLICE_X75Y104_AO6;
  assign CLBLM_R_X49Y106_SLICE_X75Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOB33_X105Y139_IOB_X1Y140_O = CLBLL_R_X57Y99_SLICE_X87Y99_AQ;
  assign RIOB33_X105Y139_IOB_X1Y139_O = CLBLM_L_X60Y111_SLICE_X91Y111_AQ;
  assign CLBLM_R_X49Y106_SLICE_X75Y106_CX = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X49Y106_SLICE_X75Y106_D1 = CLBLL_R_X57Y100_SLICE_X87Y100_CQ;
  assign CLBLM_R_X49Y106_SLICE_X75Y106_D2 = CLBLM_L_X56Y101_SLICE_X85Y101_DQ;
  assign CLBLM_R_X49Y106_SLICE_X75Y106_D3 = CLBLL_R_X57Y101_SLICE_X87Y101_CQ;
  assign CLBLM_R_X49Y106_SLICE_X75Y106_D4 = CLBLL_R_X57Y100_SLICE_X86Y100_CQ;
  assign CLBLM_R_X49Y106_SLICE_X75Y106_D5 = CLBLM_L_X56Y101_SLICE_X85Y101_CQ;
  assign CLBLM_R_X49Y106_SLICE_X75Y106_D6 = CLBLL_R_X57Y100_SLICE_X86Y100_DQ;
  assign CLBLM_R_X49Y106_SLICE_X75Y106_DX = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X49Y106_SLICE_X75Y106_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X49Y106_SLICE_X74Y106_A1 = CLBLM_R_X49Y107_SLICE_X75Y107_DO6;
  assign CLBLM_R_X49Y106_SLICE_X74Y106_A2 = CLBLM_R_X53Y101_SLICE_X81Y101_AQ;
  assign CLBLM_R_X49Y106_SLICE_X74Y106_A3 = CLBLM_R_X49Y106_SLICE_X75Y106_F7AMUX_O;
  assign CLBLM_R_X49Y106_SLICE_X74Y106_A4 = CLBLM_R_X49Y106_SLICE_X74Y106_BO6;
  assign CLBLM_R_X49Y106_SLICE_X74Y106_A5 = CLBLM_R_X53Y100_SLICE_X81Y100_AQ;
  assign CLBLM_R_X49Y106_SLICE_X74Y106_A6 = 1'b1;
  assign CLBLM_R_X49Y106_SLICE_X74Y106_B1 = CLBLL_R_X57Y99_SLICE_X86Y99_BQ;
  assign CLBLM_R_X49Y106_SLICE_X74Y106_B2 = CLBLL_R_X57Y100_SLICE_X87Y100_CQ;
  assign CLBLM_R_X49Y106_SLICE_X74Y106_B3 = CLBLL_L_X54Y100_SLICE_X82Y100_BQ;
  assign CLBLM_R_X49Y106_SLICE_X74Y106_B4 = CLBLM_R_X53Y101_SLICE_X80Y101_BQ;
  assign CLBLM_R_X49Y106_SLICE_X74Y106_B5 = 1'b1;
  assign CLBLM_R_X49Y106_SLICE_X74Y106_B6 = CLBLL_R_X57Y100_SLICE_X87Y100_AQ;
  assign CLBLM_R_X49Y106_SLICE_X74Y106_C1 = CLBLL_L_X54Y100_SLICE_X82Y100_BQ;
  assign CLBLM_R_X49Y106_SLICE_X74Y106_C2 = 1'b1;
  assign CLBLM_R_X49Y106_SLICE_X74Y106_C3 = 1'b1;
  assign CLBLM_R_X49Y106_SLICE_X74Y106_C4 = 1'b1;
  assign CLBLM_R_X49Y106_SLICE_X74Y106_C5 = CLBLM_R_X53Y101_SLICE_X81Y101_AQ;
  assign CLBLM_R_X49Y106_SLICE_X74Y106_C6 = 1'b1;
  assign CLBLM_R_X49Y106_SLICE_X74Y106_CE = CLBLM_L_X56Y98_SLICE_X84Y98_DO6;
  assign CLBLM_R_X49Y106_SLICE_X74Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X49Y106_SLICE_X74Y106_D1 = 1'b1;
  assign CLBLM_R_X49Y106_SLICE_X74Y106_D2 = 1'b1;
  assign CLBLM_R_X49Y106_SLICE_X74Y106_D3 = 1'b1;
  assign CLBLM_R_X49Y106_SLICE_X74Y106_D4 = 1'b1;
  assign CLBLM_R_X49Y106_SLICE_X74Y106_D5 = 1'b1;
  assign CLBLM_R_X49Y106_SLICE_X74Y106_D6 = 1'b1;
  assign CLBLM_R_X49Y106_SLICE_X74Y106_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_B2 = CLBLM_R_X65Y102_SLICE_X98Y102_D_XOR;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_B3 = 1'b1;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_B6 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_C2 = CLBLM_L_X60Y98_SLICE_X90Y98_AQ;
  assign CLBLM_R_X65Y102_SLICE_X99Y102_C4 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_A1 = CLBLM_L_X62Y98_SLICE_X92Y98_CQ;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_A2 = CLBLM_L_X62Y98_SLICE_X92Y98_AQ;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_A3 = CLBLM_L_X62Y98_SLICE_X92Y98_DQ;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_A4 = CLBLM_L_X56Y98_SLICE_X85Y98_DQ;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_A5 = CLBLM_L_X62Y95_SLICE_X92Y95_AQ;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_A6 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X92Y112_A1 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_AX = CLBLM_L_X62Y95_SLICE_X93Y95_BO5;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_B1 = CLBLM_L_X62Y98_SLICE_X92Y98_DQ;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_B2 = CLBLM_L_X62Y98_SLICE_X92Y98_AQ;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_B3 = CLBLM_L_X62Y95_SLICE_X92Y95_A5Q;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_B4 = CLBLM_L_X62Y98_SLICE_X92Y98_CQ;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_B5 = CLBLM_L_X62Y95_SLICE_X92Y95_AQ;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_B6 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_BX = CLBLM_L_X62Y95_SLICE_X93Y95_AO5;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_C1 = CLBLM_L_X62Y95_SLICE_X92Y95_AQ;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_C2 = CLBLM_L_X62Y95_SLICE_X92Y95_A5Q;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_C3 = CLBLM_L_X62Y98_SLICE_X92Y98_AQ;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_C4 = CLBLM_L_X62Y98_SLICE_X92Y98_CQ;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_C5 = CLBLM_L_X62Y98_SLICE_X92Y98_DQ;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_C6 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_CE = CLBLM_L_X60Y98_SLICE_X91Y98_AQ;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_D1 = CLBLM_L_X62Y95_SLICE_X92Y95_AQ;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_D2 = CLBLM_L_X62Y98_SLICE_X92Y98_CQ;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_D3 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_D4 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_D5 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_D6 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X93Y95_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_A1 = CLBLM_L_X50Y106_SLICE_X76Y106_AQ;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_A2 = CLBLM_L_X50Y104_SLICE_X76Y104_AQ;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_A3 = CLBLM_L_X62Y95_SLICE_X92Y95_AQ;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_A4 = CLBLM_L_X62Y95_SLICE_X92Y95_BO6;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_A5 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_A6 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_B1 = CLBLM_L_X56Y98_SLICE_X85Y98_DQ;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_B2 = CLBLM_L_X62Y98_SLICE_X92Y98_DQ;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_B3 = CLBLM_L_X62Y95_SLICE_X92Y95_AQ;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_B4 = CLBLM_L_X62Y98_SLICE_X92Y98_AQ;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_B5 = CLBLM_L_X62Y95_SLICE_X92Y95_A5Q;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_B6 = CLBLM_L_X62Y98_SLICE_X92Y98_CQ;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_C1 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_C2 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_C3 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_C4 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_C5 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_C6 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_CE = CLBLM_L_X62Y98_SLICE_X93Y98_CO6;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_D1 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_D2 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_D3 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_D4 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_D5 = 1'b1;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_D6 = 1'b1;
  assign CLBLM_L_X56Y102_SLICE_X85Y102_C2 = 1'b1;
  assign CLBLM_L_X56Y102_SLICE_X85Y102_C3 = CLBLM_L_X56Y102_SLICE_X85Y102_AQ;
  assign CLBLM_L_X62Y95_SLICE_X92Y95_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X56Y102_SLICE_X85Y102_C5 = 1'b1;
  assign CLBLM_R_X49Y107_SLICE_X75Y107_A1 = CLBLL_L_X54Y100_SLICE_X82Y100_BQ;
  assign CLBLM_R_X49Y107_SLICE_X75Y107_A2 = CLBLM_R_X49Y108_SLICE_X75Y108_C_XOR;
  assign CLBLM_R_X49Y107_SLICE_X75Y107_A3 = CLBLM_R_X53Y101_SLICE_X80Y101_BQ;
  assign CLBLM_R_X49Y107_SLICE_X75Y107_A4 = CLBLM_L_X50Y108_SLICE_X77Y108_C_XOR;
  assign CLBLM_R_X49Y107_SLICE_X75Y107_A5 = CLBLM_L_X50Y108_SLICE_X76Y108_C_XOR;
  assign CLBLM_R_X49Y107_SLICE_X75Y107_A6 = CLBLM_R_X49Y107_SLICE_X75Y107_CO6;
  assign RIOB33_X105Y141_IOB_X1Y141_O = CLBLM_L_X60Y98_SLICE_X90Y98_BQ;
  assign RIOB33_X105Y141_IOB_X1Y142_O = CLBLM_L_X62Y110_SLICE_X93Y110_AQ;
  assign CLBLM_R_X49Y107_SLICE_X75Y107_AX = CLBLM_R_X53Y101_SLICE_X81Y101_AQ;
  assign CLBLM_R_X49Y107_SLICE_X75Y107_B1 = CLBLL_L_X54Y100_SLICE_X82Y100_BQ;
  assign CLBLM_R_X49Y107_SLICE_X75Y107_B2 = CLBLL_R_X57Y101_SLICE_X87Y101_DQ;
  assign CLBLM_R_X49Y107_SLICE_X75Y107_B3 = 1'b1;
  assign CLBLM_R_X49Y107_SLICE_X75Y107_B4 = CLBLM_L_X56Y101_SLICE_X85Y101_AQ;
  assign CLBLM_R_X49Y107_SLICE_X75Y107_B5 = CLBLM_R_X53Y101_SLICE_X80Y101_BQ;
  assign CLBLM_R_X49Y107_SLICE_X75Y107_B6 = CLBLM_L_X56Y101_SLICE_X85Y101_CQ;
  assign CLBLM_R_X49Y107_SLICE_X75Y107_BX = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X49Y107_SLICE_X75Y107_C1 = CLBLM_R_X53Y101_SLICE_X80Y101_BQ;
  assign CLBLM_R_X49Y107_SLICE_X75Y107_C2 = CLBLM_R_X49Y108_SLICE_X75Y108_C_XOR;
  assign CLBLM_R_X49Y107_SLICE_X75Y107_C3 = CLBLL_R_X57Y97_SLICE_X86Y97_AQ;
  assign CLBLM_R_X49Y107_SLICE_X75Y107_C4 = CLBLM_R_X49Y108_SLICE_X75Y108_A_XOR;
  assign CLBLM_R_X49Y107_SLICE_X75Y107_C5 = CLBLM_R_X49Y108_SLICE_X75Y108_B_XOR;
  assign CLBLM_R_X49Y107_SLICE_X75Y107_C6 = 1'b1;
  assign CLBLM_R_X49Y107_SLICE_X75Y107_CE = CLBLM_R_X49Y104_SLICE_X75Y104_AO6;
  assign CLBLM_R_X49Y107_SLICE_X75Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X49Y107_SLICE_X75Y107_CX = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X49Y107_SLICE_X75Y107_D1 = CLBLM_R_X53Y101_SLICE_X80Y101_BQ;
  assign CLBLM_R_X49Y107_SLICE_X75Y107_D2 = CLBLL_L_X54Y100_SLICE_X82Y100_BQ;
  assign CLBLM_R_X49Y107_SLICE_X75Y107_D3 = CLBLM_L_X50Y108_SLICE_X76Y108_D_XOR;
  assign CLBLM_R_X49Y107_SLICE_X75Y107_D4 = CLBLM_R_X49Y107_SLICE_X75Y107_CO5;
  assign CLBLM_R_X49Y107_SLICE_X75Y107_D5 = CLBLM_R_X49Y108_SLICE_X75Y108_D_XOR;
  assign CLBLM_R_X49Y107_SLICE_X75Y107_D6 = CLBLM_L_X50Y108_SLICE_X77Y108_D_XOR;
  assign CLBLM_R_X49Y107_SLICE_X75Y107_DX = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X49Y107_SLICE_X75Y107_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X56Y102_SLICE_X85Y102_D1 = 1'b1;
  assign CLBLM_R_X49Y107_SLICE_X74Y107_A1 = CLBLM_R_X49Y108_SLICE_X74Y108_A5Q;
  assign CLBLM_R_X49Y107_SLICE_X74Y107_A2 = CLBLL_R_X57Y102_SLICE_X86Y102_AQ;
  assign CLBLM_R_X49Y107_SLICE_X74Y107_A3 = CLBLM_L_X50Y105_SLICE_X77Y105_AQ;
  assign CLBLM_R_X49Y107_SLICE_X74Y107_A4 = CLBLL_R_X57Y102_SLICE_X86Y102_BQ;
  assign CLBLM_R_X49Y107_SLICE_X74Y107_A5 = 1'b1;
  assign CLBLM_R_X49Y107_SLICE_X74Y107_A6 = 1'b1;
  assign CLBLM_L_X56Y102_SLICE_X85Y102_D2 = 1'b1;
  assign CLBLM_R_X49Y107_SLICE_X74Y107_B1 = CLBLM_L_X50Y109_SLICE_X77Y109_A_XOR;
  assign CLBLM_R_X49Y107_SLICE_X74Y107_B2 = CLBLL_L_X54Y100_SLICE_X82Y100_BQ;
  assign CLBLM_R_X49Y107_SLICE_X74Y107_B3 = CLBLM_R_X49Y109_SLICE_X75Y109_A_XOR;
  assign CLBLM_R_X49Y107_SLICE_X74Y107_B4 = CLBLM_L_X50Y109_SLICE_X76Y109_A_XOR;
  assign CLBLM_R_X49Y107_SLICE_X74Y107_B5 = CLBLM_R_X53Y101_SLICE_X80Y101_BQ;
  assign CLBLM_R_X49Y107_SLICE_X74Y107_B6 = CLBLM_R_X49Y107_SLICE_X74Y107_CO6;
  assign CLBLM_R_X49Y107_SLICE_X74Y107_C1 = CLBLL_R_X57Y97_SLICE_X86Y97_AQ;
  assign CLBLM_R_X49Y107_SLICE_X74Y107_C2 = CLBLM_R_X53Y101_SLICE_X80Y101_BQ;
  assign CLBLM_R_X49Y107_SLICE_X74Y107_C3 = CLBLM_R_X49Y108_SLICE_X75Y108_D_XOR;
  assign CLBLM_R_X49Y107_SLICE_X74Y107_C4 = CLBLM_R_X49Y108_SLICE_X75Y108_A_XOR;
  assign CLBLM_R_X49Y107_SLICE_X74Y107_C5 = CLBLM_R_X49Y108_SLICE_X75Y108_B_XOR;
  assign CLBLM_R_X49Y107_SLICE_X74Y107_C6 = CLBLM_R_X49Y108_SLICE_X75Y108_C_XOR;
  assign CLBLM_R_X49Y107_SLICE_X74Y107_CE = CLBLM_L_X62Y109_SLICE_X92Y109_BO6;
  assign CLBLM_R_X49Y107_SLICE_X74Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X49Y107_SLICE_X74Y107_D1 = CLBLM_L_X50Y105_SLICE_X76Y105_CO6;
  assign CLBLM_R_X49Y107_SLICE_X74Y107_D2 = CLBLM_R_X49Y108_SLICE_X75Y108_A_XOR;
  assign CLBLM_R_X49Y107_SLICE_X74Y107_D3 = CLBLM_R_X49Y108_SLICE_X75Y108_D_XOR;
  assign CLBLM_R_X49Y107_SLICE_X74Y107_D4 = CLBLM_R_X49Y109_SLICE_X75Y109_A_XOR;
  assign CLBLM_R_X49Y107_SLICE_X74Y107_D5 = CLBLM_R_X49Y108_SLICE_X75Y108_B_XOR;
  assign CLBLM_R_X49Y107_SLICE_X74Y107_D6 = CLBLM_R_X49Y108_SLICE_X75Y108_C_XOR;
  assign CLBLM_R_X49Y107_SLICE_X74Y107_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X56Y102_SLICE_X84Y102_A4 = CLBLM_L_X56Y102_SLICE_X85Y102_A5Q;
  assign CLBLM_L_X62Y96_SLICE_X93Y96_A1 = CLBLM_L_X62Y97_SLICE_X93Y97_DQ;
  assign CLBLM_L_X62Y96_SLICE_X93Y96_A2 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_L_X62Y96_SLICE_X93Y96_A3 = CLBLM_R_X63Y98_SLICE_X95Y98_D5Q;
  assign CLBLM_L_X62Y96_SLICE_X93Y96_A4 = CLBLM_L_X62Y97_SLICE_X92Y97_D5Q;
  assign CLBLM_L_X62Y96_SLICE_X93Y96_A5 = CLBLM_R_X63Y99_SLICE_X94Y99_C5Q;
  assign CLBLM_L_X62Y96_SLICE_X93Y96_A6 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_L_X62Y96_SLICE_X93Y96_AX = CLBLM_L_X62Y106_SLICE_X93Y106_CO6;
  assign CLBLM_L_X62Y96_SLICE_X93Y96_B1 = CLBLM_L_X62Y98_SLICE_X93Y98_AQ;
  assign CLBLM_L_X62Y96_SLICE_X93Y96_B2 = CLBLM_L_X62Y96_SLICE_X93Y96_BQ;
  assign CLBLM_L_X62Y96_SLICE_X93Y96_B3 = CLBLM_R_X63Y94_SLICE_X94Y94_AQ;
  assign CLBLM_L_X62Y96_SLICE_X93Y96_B4 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_L_X62Y96_SLICE_X93Y96_B5 = CLBLM_R_X63Y95_SLICE_X95Y95_D5Q;
  assign CLBLM_L_X62Y96_SLICE_X93Y96_B6 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_L_X62Y96_SLICE_X93Y96_BX = CLBLM_R_X63Y96_SLICE_X95Y96_AO6;
  assign CLBLM_L_X62Y96_SLICE_X93Y96_C1 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y96_SLICE_X93Y96_C2 = 1'b1;
  assign CLBLM_L_X62Y96_SLICE_X93Y96_C3 = CLBLM_L_X56Y98_SLICE_X85Y98_DQ;
  assign CLBLM_L_X62Y96_SLICE_X93Y96_C4 = CLBLM_R_X49Y106_SLICE_X74Y106_AQ;
  assign CLBLM_L_X62Y96_SLICE_X93Y96_C5 = CLBLM_R_X63Y100_SLICE_X95Y100_A5Q;
  assign CLBLM_L_X62Y96_SLICE_X93Y96_C6 = CLBLM_R_X63Y95_SLICE_X94Y95_AO6;
  assign CLBLM_L_X62Y96_SLICE_X93Y96_CE = CLBLM_L_X62Y99_SLICE_X93Y99_DO6;
  assign CLBLM_L_X62Y96_SLICE_X93Y96_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X62Y96_SLICE_X93Y96_D1 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y96_SLICE_X93Y96_D2 = CLBLM_L_X50Y104_SLICE_X76Y104_AQ;
  assign CLBLM_L_X62Y96_SLICE_X93Y96_D3 = CLBLM_L_X56Y98_SLICE_X85Y98_DQ;
  assign CLBLM_L_X62Y96_SLICE_X93Y96_D4 = CLBLM_L_X64Y97_SLICE_X96Y97_BQ;
  assign CLBLM_L_X62Y96_SLICE_X93Y96_D5 = 1'b1;
  assign CLBLM_L_X62Y96_SLICE_X93Y96_D6 = CLBLM_R_X63Y96_SLICE_X94Y96_CO5;
  assign CLBLM_L_X62Y96_SLICE_X93Y96_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X62Y96_SLICE_X92Y96_A1 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_L_X62Y96_SLICE_X92Y96_A2 = CLBLM_R_X63Y98_SLICE_X94Y98_C5Q;
  assign CLBLM_L_X62Y96_SLICE_X92Y96_A3 = CLBLM_L_X62Y97_SLICE_X92Y97_C5Q;
  assign CLBLM_L_X62Y96_SLICE_X92Y96_A4 = CLBLM_L_X62Y99_SLICE_X93Y99_AQ;
  assign CLBLM_L_X62Y96_SLICE_X92Y96_A5 = CLBLM_R_X63Y98_SLICE_X95Y98_C5Q;
  assign CLBLM_L_X62Y96_SLICE_X92Y96_A6 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_L_X62Y96_SLICE_X92Y96_AX = CLBLM_L_X62Y106_SLICE_X93Y106_CO6;
  assign CLBLM_L_X62Y96_SLICE_X92Y96_B1 = CLBLM_L_X62Y96_SLICE_X92Y96_CQ;
  assign CLBLM_L_X62Y96_SLICE_X92Y96_B2 = 1'b1;
  assign CLBLM_L_X62Y96_SLICE_X92Y96_B3 = CLBLM_R_X63Y95_SLICE_X95Y95_B5Q;
  assign CLBLM_L_X62Y96_SLICE_X92Y96_B4 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_L_X62Y96_SLICE_X92Y96_B5 = CLBLM_R_X63Y96_SLICE_X95Y96_AQ;
  assign CLBLM_L_X62Y96_SLICE_X92Y96_B6 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_L_X62Y96_SLICE_X92Y96_C1 = CLBLM_L_X50Y106_SLICE_X76Y106_CQ;
  assign CLBLM_L_X62Y96_SLICE_X92Y96_C2 = CLBLM_R_X63Y96_SLICE_X94Y96_AO6;
  assign CLBLM_L_X62Y96_SLICE_X92Y96_C3 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y96_SLICE_X92Y96_C4 = CLBLM_R_X63Y98_SLICE_X95Y98_B5Q;
  assign CLBLM_L_X62Y96_SLICE_X92Y96_C5 = CLBLM_L_X56Y98_SLICE_X85Y98_DQ;
  assign CLBLM_L_X62Y96_SLICE_X92Y96_C6 = 1'b1;
  assign CLBLM_L_X62Y96_SLICE_X92Y96_CE = CLBLM_L_X62Y99_SLICE_X93Y99_AO6;
  assign CLBLM_L_X62Y96_SLICE_X92Y96_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign RIOB33_X105Y143_IOB_X1Y143_O = CLBLM_L_X56Y111_SLICE_X84Y111_AQ;
  assign RIOB33_X105Y143_IOB_X1Y144_O = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X62Y96_SLICE_X92Y96_D1 = 1'b1;
  assign CLBLM_L_X62Y96_SLICE_X92Y96_D2 = 1'b1;
  assign CLBLM_L_X62Y96_SLICE_X92Y96_D3 = 1'b1;
  assign CLBLM_L_X62Y96_SLICE_X92Y96_D4 = 1'b1;
  assign CLBLM_L_X62Y96_SLICE_X92Y96_D5 = 1'b1;
  assign CLBLM_L_X62Y96_SLICE_X92Y96_D6 = 1'b1;
  assign CLBLM_L_X62Y96_SLICE_X92Y96_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_A1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_A2 = CLBLL_R_X57Y100_SLICE_X86Y100_DQ;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_A3 = CLBLL_R_X57Y100_SLICE_X86Y100_AQ;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_A4 = 1'b1;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_A5 = 1'b1;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_A6 = 1'b1;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_AX = CLBLL_R_X57Y100_SLICE_X86Y100_AQ;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_B1 = 1'b1;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_B2 = CLBLL_R_X57Y100_SLICE_X86Y100_BQ;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_B3 = CLBLL_R_X57Y100_SLICE_X86Y100_CQ;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_B4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_B5 = 1'b1;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_B6 = 1'b1;
  assign CLBLM_L_X56Y102_SLICE_X84Y102_D6 = 1'b1;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_BX = CLBLL_R_X57Y100_SLICE_X86Y100_BQ;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_C1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_C2 = CLBLM_L_X56Y101_SLICE_X85Y101_CQ;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_C3 = 1'b1;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_C4 = 1'b1;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_C5 = CLBLM_L_X56Y101_SLICE_X85Y101_AQ;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_C6 = 1'b1;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_CE = CLBLM_R_X49Y104_SLICE_X75Y104_AO6;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_CX = CLBLM_L_X56Y101_SLICE_X85Y101_AQ;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_D1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_D2 = 1'b1;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_D3 = CLBLL_R_X57Y100_SLICE_X87Y100_CQ;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_D4 = 1'b1;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_D5 = CLBLL_R_X57Y100_SLICE_X87Y100_AQ;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_D6 = 1'b1;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_DX = CLBLL_R_X57Y100_SLICE_X87Y100_AQ;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X49Y108_SLICE_X74Y108_A1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X49Y108_SLICE_X74Y108_A2 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X49Y108_SLICE_X74Y108_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X49Y108_SLICE_X74Y108_A4 = CLBLM_L_X62Y105_SLICE_X92Y105_CQ;
  assign CLBLM_R_X49Y108_SLICE_X74Y108_A5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X49Y108_SLICE_X74Y108_A6 = 1'b1;
  assign CLBLM_R_X49Y108_SLICE_X74Y108_B1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X49Y108_SLICE_X74Y108_B2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X49Y108_SLICE_X74Y108_B3 = CLBLM_L_X62Y105_SLICE_X92Y105_CQ;
  assign CLBLM_R_X49Y108_SLICE_X74Y108_B4 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X49Y108_SLICE_X74Y108_B5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X49Y108_SLICE_X74Y108_B6 = 1'b1;
  assign CLBLM_R_X49Y108_SLICE_X74Y108_C1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X49Y108_SLICE_X74Y108_C2 = CLBLM_L_X62Y105_SLICE_X92Y105_CQ;
  assign CLBLM_R_X49Y108_SLICE_X74Y108_C3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X49Y108_SLICE_X74Y108_C4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X49Y108_SLICE_X74Y108_C5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X49Y108_SLICE_X74Y108_C6 = 1'b1;
  assign CLBLM_R_X49Y108_SLICE_X74Y108_CE = CLBLM_R_X49Y110_SLICE_X74Y110_BO6;
  assign CLBLM_R_X49Y108_SLICE_X74Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X49Y108_SLICE_X74Y108_D1 = CLBLM_L_X50Y109_SLICE_X77Y109_B_XOR;
  assign CLBLM_R_X49Y108_SLICE_X74Y108_D2 = CLBLL_L_X54Y100_SLICE_X82Y100_BQ;
  assign CLBLM_R_X49Y108_SLICE_X74Y108_D3 = CLBLM_R_X49Y107_SLICE_X74Y107_DO6;
  assign CLBLM_R_X49Y108_SLICE_X74Y108_D4 = CLBLM_L_X50Y109_SLICE_X76Y109_B_XOR;
  assign CLBLM_R_X49Y108_SLICE_X74Y108_D5 = CLBLM_R_X49Y109_SLICE_X75Y109_B_XOR;
  assign CLBLM_R_X49Y108_SLICE_X74Y108_D6 = CLBLM_R_X53Y101_SLICE_X80Y101_BQ;
  assign CLBLM_R_X49Y108_SLICE_X74Y108_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_A1 = CLBLM_L_X62Y97_SLICE_X93Y97_CQ;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_A2 = CLBLM_R_X63Y98_SLICE_X95Y98_DQ;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_A3 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_A4 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_A5 = CLBLM_L_X62Y97_SLICE_X92Y97_DQ;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_A6 = CLBLM_R_X63Y99_SLICE_X94Y99_CQ;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_AX = CLBLM_L_X62Y106_SLICE_X93Y106_CO6;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_B1 = CLBLM_R_X63Y97_SLICE_X94Y97_CQ;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_B2 = CLBLM_R_X63Y95_SLICE_X95Y95_C5Q;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_B3 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_B4 = CLBLM_L_X64Y97_SLICE_X97Y97_BQ;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_B5 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_B6 = CLBLM_L_X62Y98_SLICE_X93Y98_BQ;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_BX = CLBLM_R_X63Y97_SLICE_X94Y97_CO6;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_C1 = CLBLM_L_X50Y107_SLICE_X76Y107_BQ;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_C2 = CLBLM_L_X64Y96_SLICE_X96Y96_AO5;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_C3 = CLBLM_L_X56Y98_SLICE_X85Y98_DQ;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_C4 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_C5 = CLBLM_R_X63Y98_SLICE_X95Y98_DQ;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_C6 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_CE = CLBLM_L_X62Y100_SLICE_X92Y100_DO6;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_D1 = CLBLM_L_X62Y96_SLICE_X92Y96_CQ;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_D2 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_D3 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_D4 = CLBLM_L_X56Y97_SLICE_X85Y97_AQ;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_D5 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_D6 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_DX = CLBLM_R_X63Y96_SLICE_X95Y96_AO6;
  assign CLBLM_L_X62Y97_SLICE_X93Y97_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_A1 = CLBLM_L_X50Y104_SLICE_X76Y104_AQ;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_A2 = CLBLM_L_X62Y100_SLICE_X92Y100_AQ;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_A3 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_A4 = CLBLM_L_X64Y97_SLICE_X96Y97_BQ;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_A5 = CLBLM_L_X62Y100_SLICE_X92Y100_AO6;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_A6 = 1'b1;
  assign RIOB33_X105Y145_IOB_X1Y145_O = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_B1 = CLBLM_L_X50Y105_SLICE_X77Y105_AQ;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_B2 = CLBLM_L_X64Y97_SLICE_X96Y97_B5Q;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_B3 = CLBLM_L_X62Y100_SLICE_X92Y100_BQ;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_B4 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_B5 = CLBLM_L_X62Y100_SLICE_X92Y100_AO6;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_B6 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_C1 = CLBLM_L_X62Y100_SLICE_X92Y100_AO6;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_C2 = CLBLM_L_X50Y106_SLICE_X76Y106_CQ;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_C3 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_C4 = CLBLM_L_X50Y106_SLICE_X76Y106_AQ;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_C5 = CLBLM_L_X60Y97_SLICE_X91Y97_BQ;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_C6 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_CE = CLBLM_L_X62Y100_SLICE_X92Y100_BO6;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_D1 = CLBLM_L_X62Y100_SLICE_X92Y100_AO6;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_D2 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_D3 = CLBLM_L_X50Y107_SLICE_X76Y107_BQ;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_D4 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_D5 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_D6 = 1'b1;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_DX = CLBLM_L_X60Y97_SLICE_X91Y97_AO5;
  assign CLBLM_L_X62Y97_SLICE_X92Y97_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X49Y109_SLICE_X75Y109_A1 = 1'b1;
  assign CLBLM_R_X49Y109_SLICE_X75Y109_A2 = 1'b1;
  assign CLBLM_R_X49Y109_SLICE_X75Y109_A3 = CLBLL_R_X57Y101_SLICE_X87Y101_CQ;
  assign CLBLM_R_X49Y109_SLICE_X75Y109_A4 = 1'b1;
  assign CLBLM_R_X49Y109_SLICE_X75Y109_A5 = CLBLL_R_X57Y101_SLICE_X87Y101_AQ;
  assign CLBLM_R_X49Y109_SLICE_X75Y109_A6 = 1'b1;
  assign CLBLM_R_X49Y109_SLICE_X75Y109_AX = CLBLL_R_X57Y101_SLICE_X87Y101_AQ;
  assign CLBLM_R_X49Y109_SLICE_X75Y109_B1 = 1'b1;
  assign CLBLM_R_X49Y109_SLICE_X75Y109_B2 = 1'b1;
  assign CLBLM_R_X49Y109_SLICE_X75Y109_B3 = 1'b1;
  assign CLBLM_R_X49Y109_SLICE_X75Y109_B4 = CLBLM_L_X56Y101_SLICE_X85Y101_DQ;
  assign CLBLM_R_X49Y109_SLICE_X75Y109_B5 = CLBLM_L_X56Y101_SLICE_X85Y101_BQ;
  assign CLBLM_R_X49Y109_SLICE_X75Y109_B6 = 1'b1;
  assign CLBLM_R_X49Y109_SLICE_X75Y109_BX = CLBLM_L_X56Y101_SLICE_X85Y101_BQ;
  assign CLBLM_R_X49Y109_SLICE_X75Y109_C1 = 1'b1;
  assign CLBLM_R_X49Y109_SLICE_X75Y109_C2 = CLBLL_R_X57Y100_SLICE_X87Y100_BQ;
  assign CLBLM_R_X49Y109_SLICE_X75Y109_C3 = 1'b1;
  assign CLBLM_R_X49Y109_SLICE_X75Y109_C4 = CLBLL_R_X57Y101_SLICE_X87Y101_DQ;
  assign CLBLM_R_X49Y109_SLICE_X75Y109_C5 = 1'b1;
  assign CLBLM_R_X49Y109_SLICE_X75Y109_C6 = 1'b1;
  assign CLBLM_R_X49Y109_SLICE_X75Y109_CIN = CLBLM_R_X49Y108_SLICE_X75Y108_COUT;
  assign CLBLM_R_X49Y109_SLICE_X75Y109_CX = CLBLL_R_X57Y100_SLICE_X87Y100_BQ;
  assign CLBLM_R_X49Y109_SLICE_X75Y109_D1 = CLBLL_R_X57Y99_SLICE_X86Y99_BQ;
  assign CLBLM_R_X49Y109_SLICE_X75Y109_D2 = 1'b1;
  assign CLBLM_R_X49Y109_SLICE_X75Y109_D3 = 1'b1;
  assign CLBLM_R_X49Y109_SLICE_X75Y109_D4 = 1'b1;
  assign CLBLM_R_X49Y109_SLICE_X75Y109_D5 = CLBLL_R_X57Y99_SLICE_X86Y99_AQ;
  assign CLBLM_R_X49Y109_SLICE_X75Y109_D6 = 1'b1;
  assign CLBLM_R_X49Y109_SLICE_X75Y109_DX = CLBLL_R_X57Y99_SLICE_X86Y99_AQ;
  assign CLBLM_R_X49Y109_SLICE_X74Y109_A1 = CLBLL_R_X57Y102_SLICE_X86Y102_AQ;
  assign CLBLM_R_X49Y109_SLICE_X74Y109_A2 = CLBLM_R_X49Y108_SLICE_X74Y108_BQ;
  assign CLBLM_R_X49Y109_SLICE_X74Y109_A3 = 1'b1;
  assign CLBLM_R_X49Y109_SLICE_X74Y109_A4 = CLBLL_R_X57Y102_SLICE_X86Y102_BQ;
  assign CLBLM_R_X49Y109_SLICE_X74Y109_A5 = CLBLM_L_X50Y106_SLICE_X76Y106_AQ;
  assign CLBLM_R_X49Y109_SLICE_X74Y109_A6 = 1'b1;
  assign CLBLM_R_X49Y109_SLICE_X74Y109_B1 = CLBLL_R_X57Y102_SLICE_X86Y102_AQ;
  assign CLBLM_R_X49Y109_SLICE_X74Y109_B2 = 1'b1;
  assign CLBLM_R_X49Y109_SLICE_X74Y109_B3 = CLBLM_L_X50Y106_SLICE_X76Y106_CQ;
  assign CLBLM_R_X49Y109_SLICE_X74Y109_B4 = CLBLL_R_X57Y102_SLICE_X86Y102_BQ;
  assign CLBLM_R_X49Y109_SLICE_X74Y109_B5 = 1'b1;
  assign CLBLM_R_X49Y109_SLICE_X74Y109_B6 = CLBLM_R_X49Y108_SLICE_X74Y108_B5Q;
  assign CLBLM_R_X49Y109_SLICE_X74Y109_C1 = CLBLM_R_X49Y108_SLICE_X74Y108_C5Q;
  assign CLBLM_R_X49Y109_SLICE_X74Y109_C2 = 1'b1;
  assign CLBLM_R_X49Y109_SLICE_X74Y109_C3 = CLBLM_L_X50Y107_SLICE_X77Y107_AQ;
  assign CLBLM_R_X49Y109_SLICE_X74Y109_C4 = CLBLL_R_X57Y102_SLICE_X86Y102_BQ;
  assign CLBLM_R_X49Y109_SLICE_X74Y109_C5 = CLBLL_R_X57Y102_SLICE_X86Y102_AQ;
  assign CLBLM_R_X49Y109_SLICE_X74Y109_C6 = 1'b1;
  assign CLBLM_R_X49Y109_SLICE_X74Y109_CE = CLBLM_L_X62Y109_SLICE_X92Y109_BO6;
  assign CLBLM_R_X49Y109_SLICE_X74Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X49Y109_SLICE_X74Y109_D1 = CLBLM_L_X50Y104_SLICE_X76Y104_AQ;
  assign CLBLM_R_X49Y109_SLICE_X74Y109_D2 = 1'b1;
  assign CLBLM_R_X49Y109_SLICE_X74Y109_D3 = CLBLL_R_X57Y102_SLICE_X86Y102_AQ;
  assign CLBLM_R_X49Y109_SLICE_X74Y109_D4 = 1'b1;
  assign CLBLM_R_X49Y109_SLICE_X74Y109_D5 = CLBLM_R_X49Y108_SLICE_X74Y108_AQ;
  assign CLBLM_R_X49Y109_SLICE_X74Y109_D6 = CLBLL_R_X57Y102_SLICE_X86Y102_BQ;
  assign CLBLM_R_X49Y109_SLICE_X74Y109_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_A1 = CLBLM_R_X49Y119_SLICE_X74Y119_AQ;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_A2 = CLBLM_R_X49Y119_SLICE_X74Y119_BQ;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_A3 = CLBLM_L_X62Y95_SLICE_X93Y95_BO6;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_A4 = CLBLM_L_X62Y98_SLICE_X92Y98_BQ;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_A5 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_A6 = CLBLM_L_X62Y98_SLICE_X93Y98_AQ;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_B1 = CLBLM_R_X49Y119_SLICE_X74Y119_AQ;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_B2 = CLBLM_R_X49Y119_SLICE_X74Y119_BQ;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_B3 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_B4 = CLBLM_L_X62Y98_SLICE_X92Y98_BQ;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_B5 = CLBLM_L_X62Y95_SLICE_X93Y95_CO6;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_B6 = CLBLM_L_X62Y98_SLICE_X93Y98_BQ;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_C1 = CLBLM_L_X62Y99_SLICE_X92Y99_AO6;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_C2 = CLBLM_L_X62Y100_SLICE_X93Y100_CO6;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_C3 = CLBLM_R_X59Y102_SLICE_X88Y102_AQ;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_C4 = CLBLL_R_X57Y101_SLICE_X86Y101_AO5;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_C5 = CLBLM_L_X62Y98_SLICE_X93Y98_DO6;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_C6 = CLBLM_L_X60Y98_SLICE_X90Y98_BQ;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_D1 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_D2 = CLBLM_L_X56Y98_SLICE_X85Y98_A5Q;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_D3 = CLBLM_L_X56Y98_SLICE_X85Y98_DQ;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_D4 = CLBLM_L_X62Y98_SLICE_X93Y98_BQ;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_D5 = CLBLM_L_X62Y98_SLICE_X93Y98_AQ;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_D6 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y98_SLICE_X93Y98_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_A1 = CLBLM_R_X49Y104_SLICE_X75Y104_CQ;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_A2 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_A3 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_A4 = CLBLM_R_X49Y106_SLICE_X74Y106_AQ;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_A5 = CLBLM_L_X62Y95_SLICE_X93Y95_AO6;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_A6 = 1'b1;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_B1 = CLBLM_L_X56Y98_SLICE_X85Y98_DQ;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_B2 = CLBLM_L_X62Y98_SLICE_X92Y98_BQ;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_B3 = CLBLM_L_X62Y95_SLICE_X93Y95_CO6;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_B4 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_B5 = CLBLM_L_X62Y95_SLICE_X93Y95_BO6;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_B6 = CLBLM_L_X50Y106_SLICE_X76Y106_CQ;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_C1 = 1'b1;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_C2 = CLBLM_L_X62Y98_SLICE_X92Y98_CQ;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_C3 = CLBLM_L_X56Y98_SLICE_X85Y98_DQ;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_C4 = CLBLM_L_X50Y105_SLICE_X77Y105_AQ;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_C5 = CLBLM_L_X62Y95_SLICE_X92Y95_AQ;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_C6 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_CE = CLBLM_L_X62Y98_SLICE_X93Y98_CO6;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_D1 = CLBLM_L_X62Y98_SLICE_X92Y98_DQ;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_D2 = CLBLM_L_X62Y98_SLICE_X92Y98_CQ;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_D3 = CLBLM_L_X56Y98_SLICE_X85Y98_DQ;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_D4 = CLBLM_R_X49Y105_SLICE_X75Y105_CQ;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_D5 = CLBLM_L_X62Y95_SLICE_X92Y95_AQ;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_D6 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y98_SLICE_X92Y98_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X49Y110_SLICE_X75Y110_A1 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X75Y110_A2 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X75Y110_A3 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X75Y110_A4 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X75Y110_A5 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X75Y110_A6 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X75Y110_AX = 1'b0;
  assign CLBLM_R_X49Y110_SLICE_X75Y110_B1 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X75Y110_B2 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X75Y110_B3 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X75Y110_B4 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X75Y110_B5 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X75Y110_B6 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X75Y110_BX = 1'b0;
  assign CLBLM_R_X49Y110_SLICE_X75Y110_C1 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X75Y110_C2 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X75Y110_C3 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X75Y110_C4 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X75Y110_C5 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X75Y110_C6 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X75Y110_CIN = CLBLM_R_X49Y109_SLICE_X75Y109_COUT;
  assign CLBLM_R_X49Y110_SLICE_X75Y110_CX = 1'b0;
  assign CLBLM_R_X49Y110_SLICE_X75Y110_D1 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X75Y110_D2 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X75Y110_D3 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X75Y110_D4 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X75Y110_D5 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X75Y110_D6 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X75Y110_DX = 1'b0;
  assign CLBLM_R_X49Y110_SLICE_X74Y110_A1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X49Y110_SLICE_X74Y110_A2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X49Y110_SLICE_X74Y110_A3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X49Y110_SLICE_X74Y110_A4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X49Y110_SLICE_X74Y110_A5 = CLBLM_L_X62Y105_SLICE_X92Y105_CQ;
  assign CLBLM_R_X49Y110_SLICE_X74Y110_A6 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X74Y110_B1 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X74Y110_B2 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X74Y110_B3 = CLBLM_R_X49Y119_SLICE_X74Y119_AQ;
  assign CLBLM_R_X49Y110_SLICE_X74Y110_B4 = CLBLM_R_X49Y119_SLICE_X74Y119_BQ;
  assign CLBLM_R_X49Y110_SLICE_X74Y110_B5 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X49Y110_SLICE_X74Y110_B6 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X49Y110_SLICE_X74Y110_C1 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X74Y110_C2 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X74Y110_C3 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X74Y110_C4 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X74Y110_C5 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X74Y110_C6 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X74Y110_CE = CLBLM_R_X49Y110_SLICE_X74Y110_BO6;
  assign CLBLM_R_X49Y110_SLICE_X74Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X49Y110_SLICE_X74Y110_D1 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X74Y110_D2 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X74Y110_D3 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X74Y110_D4 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X74Y110_D5 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X74Y110_D6 = 1'b1;
  assign CLBLM_R_X49Y110_SLICE_X74Y110_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_A1 = CLBLM_L_X56Y98_SLICE_X85Y98_DQ;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_A2 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_A3 = CLBLM_L_X62Y99_SLICE_X92Y99_AO5;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_A4 = CLBLM_L_X62Y99_SLICE_X93Y99_BO6;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_A5 = CLBLM_L_X60Y99_SLICE_X90Y99_AO6;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_A6 = CLBLM_L_X56Y98_SLICE_X85Y98_A5Q;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_AX = CLBLM_R_X63Y95_SLICE_X95Y95_AO6;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_B1 = CLBLM_L_X62Y103_SLICE_X92Y103_AQ;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_B2 = CLBLM_L_X62Y106_SLICE_X93Y106_AQ;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_B3 = CLBLM_L_X62Y110_SLICE_X92Y110_DO6;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_B4 = CLBLM_L_X62Y104_SLICE_X93Y104_AQ;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_B5 = CLBLM_R_X59Y102_SLICE_X89Y102_AQ;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_B6 = CLBLM_L_X60Y110_SLICE_X91Y110_AQ;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_C1 = CLBLM_L_X60Y99_SLICE_X91Y99_AO6;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_C2 = CLBLM_L_X62Y99_SLICE_X92Y99_AO5;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_C3 = CLBLM_L_X62Y100_SLICE_X93Y100_CO6;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_C4 = CLBLM_L_X56Y98_SLICE_X85Y98_A5Q;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_C5 = CLBLM_L_X56Y98_SLICE_X85Y98_DQ;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_C6 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_CE = CLBLM_L_X62Y100_SLICE_X92Y100_DO6;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_D1 = CLBLM_L_X60Y99_SLICE_X91Y99_AO6;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_D2 = CLBLM_L_X62Y99_SLICE_X92Y99_AO5;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_D3 = CLBLM_L_X56Y98_SLICE_X85Y98_DQ;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_D4 = CLBLM_L_X56Y98_SLICE_X85Y98_A5Q;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_D5 = CLBLM_L_X62Y99_SLICE_X93Y99_BO6;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_D6 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y99_SLICE_X93Y99_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_A1 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_A2 = CLBLM_R_X49Y119_SLICE_X74Y119_BQ;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_A3 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_A4 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_A5 = CLBLM_R_X49Y119_SLICE_X74Y119_AQ;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_A6 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_B1 = CLBLM_L_X62Y110_SLICE_X92Y110_DO6;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_B2 = CLBLM_L_X62Y99_SLICE_X92Y99_BQ;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_B3 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_B4 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_B5 = CLBLL_R_X57Y99_SLICE_X87Y99_AQ;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_B6 = CLBLM_L_X62Y99_SLICE_X92Y99_CO6;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_C1 = CLBLM_L_X62Y104_SLICE_X93Y104_AQ;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_C2 = CLBLM_L_X60Y110_SLICE_X91Y110_AQ;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_C3 = CLBLM_L_X62Y103_SLICE_X92Y103_AQ;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_C4 = CLBLM_R_X59Y102_SLICE_X88Y102_AQ;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_C5 = CLBLM_R_X59Y102_SLICE_X89Y102_AQ;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_C6 = CLBLM_L_X62Y106_SLICE_X93Y106_AQ;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_D1 = CLBLL_R_X57Y99_SLICE_X87Y99_AQ;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_D2 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_D3 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_D4 = CLBLM_L_X62Y99_SLICE_X92Y99_CO6;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_D5 = 1'b1;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_D6 = 1'b1;
  assign CLBLM_R_X53Y98_SLICE_X81Y98_C1 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLM_L_X62Y99_SLICE_X92Y99_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X49Y111_SLICE_X75Y111_A1 = 1'b1;
  assign CLBLM_R_X49Y111_SLICE_X75Y111_A2 = CLBLM_L_X62Y105_SLICE_X92Y105_CQ;
  assign CLBLM_R_X49Y111_SLICE_X75Y111_A3 = 1'b1;
  assign CLBLM_R_X49Y111_SLICE_X75Y111_A4 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X49Y111_SLICE_X75Y111_A5 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X49Y111_SLICE_X75Y111_A6 = 1'b1;
  assign CLBLM_R_X53Y98_SLICE_X81Y98_C5 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign CLBLM_R_X49Y111_SLICE_X75Y111_B1 = 1'b1;
  assign CLBLM_R_X49Y111_SLICE_X75Y111_B2 = CLBLM_R_X49Y119_SLICE_X74Y119_BQ;
  assign CLBLM_R_X49Y111_SLICE_X75Y111_B3 = 1'b1;
  assign CLBLM_R_X49Y111_SLICE_X75Y111_B4 = 1'b1;
  assign CLBLM_R_X49Y111_SLICE_X75Y111_B5 = CLBLM_R_X49Y119_SLICE_X74Y119_AQ;
  assign CLBLM_R_X49Y111_SLICE_X75Y111_B6 = 1'b1;
  assign CLBLM_R_X49Y111_SLICE_X75Y111_C1 = 1'b1;
  assign CLBLM_R_X49Y111_SLICE_X75Y111_C2 = 1'b1;
  assign CLBLM_R_X49Y111_SLICE_X75Y111_C3 = 1'b1;
  assign CLBLM_R_X49Y111_SLICE_X75Y111_C4 = 1'b1;
  assign CLBLM_R_X49Y111_SLICE_X75Y111_C5 = 1'b1;
  assign CLBLM_R_X49Y111_SLICE_X75Y111_C6 = 1'b1;
  assign CLBLM_R_X49Y111_SLICE_X75Y111_CE = CLBLM_R_X49Y111_SLICE_X75Y111_BO6;
  assign CLBLM_R_X49Y111_SLICE_X75Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X49Y111_SLICE_X75Y111_D1 = 1'b1;
  assign CLBLM_R_X49Y111_SLICE_X75Y111_D2 = 1'b1;
  assign CLBLM_R_X49Y111_SLICE_X75Y111_D3 = 1'b1;
  assign CLBLM_R_X49Y111_SLICE_X75Y111_D4 = 1'b1;
  assign CLBLM_R_X49Y111_SLICE_X75Y111_D5 = 1'b1;
  assign CLBLM_R_X49Y111_SLICE_X75Y111_D6 = 1'b1;
  assign CLBLM_R_X49Y111_SLICE_X75Y111_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X49Y111_SLICE_X74Y111_A1 = 1'b1;
  assign CLBLM_R_X49Y111_SLICE_X74Y111_A2 = CLBLL_R_X57Y102_SLICE_X86Y102_AQ;
  assign CLBLM_R_X49Y111_SLICE_X74Y111_A3 = 1'b1;
  assign CLBLM_R_X49Y111_SLICE_X74Y111_A4 = CLBLL_R_X57Y102_SLICE_X86Y102_BQ;
  assign CLBLM_R_X49Y111_SLICE_X74Y111_A5 = CLBLM_R_X49Y110_SLICE_X74Y110_AQ;
  assign CLBLM_R_X49Y111_SLICE_X74Y111_A6 = CLBLM_R_X49Y105_SLICE_X75Y105_CQ;
  assign CLBLM_R_X49Y111_SLICE_X74Y111_B1 = 1'b1;
  assign CLBLM_R_X49Y111_SLICE_X74Y111_B2 = CLBLM_R_X49Y106_SLICE_X74Y106_AQ;
  assign CLBLM_R_X49Y111_SLICE_X74Y111_B3 = CLBLM_R_X49Y110_SLICE_X74Y110_A5Q;
  assign CLBLM_R_X49Y111_SLICE_X74Y111_B4 = CLBLL_R_X57Y102_SLICE_X86Y102_BQ;
  assign CLBLM_R_X49Y111_SLICE_X74Y111_B5 = 1'b1;
  assign CLBLM_R_X49Y111_SLICE_X74Y111_B6 = CLBLL_R_X57Y102_SLICE_X86Y102_AQ;
  assign CLBLM_R_X49Y111_SLICE_X74Y111_C1 = CLBLM_L_X50Y107_SLICE_X76Y107_BQ;
  assign CLBLM_R_X49Y111_SLICE_X74Y111_C2 = CLBLM_R_X49Y108_SLICE_X74Y108_CQ;
  assign CLBLM_R_X49Y111_SLICE_X74Y111_C3 = CLBLL_R_X57Y102_SLICE_X86Y102_AQ;
  assign CLBLM_R_X49Y111_SLICE_X74Y111_C4 = CLBLL_R_X57Y102_SLICE_X86Y102_BQ;
  assign CLBLM_R_X49Y111_SLICE_X74Y111_C5 = 1'b1;
  assign CLBLM_R_X49Y111_SLICE_X74Y111_C6 = 1'b1;
  assign CLBLM_R_X49Y111_SLICE_X74Y111_CE = CLBLM_L_X62Y109_SLICE_X92Y109_BO6;
  assign CLBLM_R_X53Y98_SLICE_X81Y98_D4 = 1'b1;
  assign CLBLM_R_X53Y98_SLICE_X81Y98_D5 = 1'b1;
  assign CLBLM_R_X49Y111_SLICE_X74Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X53Y98_SLICE_X81Y98_D6 = 1'b1;
  assign CLBLM_R_X49Y111_SLICE_X74Y111_D1 = 1'b1;
  assign CLBLM_R_X49Y111_SLICE_X74Y111_D2 = 1'b1;
  assign CLBLM_R_X49Y111_SLICE_X74Y111_D3 = 1'b1;
  assign CLBLM_R_X49Y111_SLICE_X74Y111_D4 = 1'b1;
  assign CLBLM_R_X49Y111_SLICE_X74Y111_D5 = 1'b1;
  assign CLBLM_R_X49Y111_SLICE_X74Y111_D6 = 1'b1;
  assign CLBLM_R_X49Y111_SLICE_X74Y111_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X53Y98_SLICE_X80Y98_B4 = 1'b1;
  assign CLBLM_R_X53Y98_SLICE_X80Y98_B5 = 1'b1;
  assign CLBLM_R_X53Y98_SLICE_X80Y98_B6 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_A1 = CLBLM_R_X49Y105_SLICE_X75Y105_CQ;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_A2 = CLBLM_R_X63Y100_SLICE_X95Y100_AQ;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_A3 = CLBLM_L_X62Y100_SLICE_X92Y100_AO6;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_A4 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_A5 = CLBLM_L_X62Y101_SLICE_X93Y101_AQ;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_A6 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_B1 = CLBLM_R_X63Y100_SLICE_X95Y100_A5Q;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_B2 = CLBLM_L_X62Y100_SLICE_X92Y100_CQ;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_B3 = CLBLM_L_X62Y100_SLICE_X92Y100_AO6;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_B4 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_B5 = CLBLM_R_X49Y106_SLICE_X74Y106_AQ;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_B6 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_C1 = CLBLM_L_X62Y103_SLICE_X92Y103_AQ;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_C2 = CLBLM_L_X62Y104_SLICE_X93Y104_AQ;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_C3 = CLBLM_R_X59Y102_SLICE_X89Y102_AQ;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_C4 = CLBLM_L_X60Y110_SLICE_X91Y110_AQ;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_C5 = CLBLM_L_X62Y110_SLICE_X92Y110_DO6;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_C6 = CLBLM_L_X62Y106_SLICE_X93Y106_AQ;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_CE = CLBLM_L_X62Y100_SLICE_X92Y100_BO6;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_D1 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_D2 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_D3 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_D4 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_D5 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_D6 = 1'b1;
  assign CLBLM_L_X56Y103_SLICE_X85Y103_B1 = CLBLL_L_X54Y105_SLICE_X82Y105_B_XOR;
  assign CLBLM_L_X62Y100_SLICE_X93Y100_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_A1 = CLBLM_R_X59Y102_SLICE_X89Y102_AQ;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_A2 = CLBLM_L_X62Y102_SLICE_X93Y102_AO5;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_A3 = CLBLM_L_X62Y104_SLICE_X93Y104_AQ;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_A4 = CLBLM_R_X59Y102_SLICE_X88Y102_AQ;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_A5 = CLBLM_L_X60Y98_SLICE_X90Y98_BQ;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_A6 = 1'b1;
  assign CLBLM_R_X53Y98_SLICE_X80Y98_C6 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_AX = CLBLM_R_X49Y104_SLICE_X74Y104_AQ;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_B1 = CLBLM_L_X56Y103_SLICE_X85Y103_CO6;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_B2 = CLBLM_L_X62Y102_SLICE_X93Y102_AO5;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_B3 = CLBLM_R_X59Y102_SLICE_X89Y102_AQ;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_B4 = CLBLM_R_X59Y102_SLICE_X88Y102_AQ;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_B5 = CLBLM_L_X60Y98_SLICE_X90Y98_BQ;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_B6 = CLBLM_L_X62Y104_SLICE_X93Y104_AQ;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_BX = CLBLM_R_X49Y104_SLICE_X75Y104_AQ;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_C1 = CLBLM_L_X60Y99_SLICE_X90Y99_AO6;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_C2 = CLBLM_L_X60Y99_SLICE_X91Y99_BO6;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_C3 = CLBLM_R_X59Y102_SLICE_X89Y102_AQ;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_C4 = CLBLM_L_X62Y104_SLICE_X93Y104_AQ;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_C5 = CLBLM_L_X62Y99_SLICE_X92Y99_AO6;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_C6 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_CE = CLBLM_L_X62Y101_SLICE_X93Y101_AO6;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_CX = CLBLM_R_X49Y104_SLICE_X75Y104_CQ;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_D1 = CLBLM_L_X60Y99_SLICE_X90Y99_AO6;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_D2 = CLBLM_L_X62Y104_SLICE_X93Y104_AQ;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_D3 = CLBLM_R_X59Y102_SLICE_X89Y102_AQ;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_D4 = CLBLM_L_X62Y102_SLICE_X93Y102_AO5;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_D5 = CLBLM_L_X62Y99_SLICE_X92Y99_AO6;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_D6 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X56Y103_SLICE_X85Y103_C1 = 1'b1;
  assign CLBLM_L_X62Y100_SLICE_X92Y100_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X56Y103_SLICE_X85Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X56Y103_SLICE_X85Y103_D1 = 1'b1;
  assign CLBLM_L_X56Y103_SLICE_X85Y103_D2 = 1'b1;
  assign CLBLM_L_X56Y103_SLICE_X85Y103_D4 = 1'b1;
  assign CLBLL_R_X57Y110_SLICE_X86Y110_C2 = 1'b1;
  assign CLBLL_R_X57Y110_SLICE_X86Y110_C4 = 1'b1;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_A1 = 1'b1;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_A2 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_A3 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_A4 = CLBLM_R_X49Y119_SLICE_X74Y119_BQ;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_A5 = CLBLM_R_X49Y119_SLICE_X74Y119_AQ;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_A6 = 1'b1;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_AX = CLBLM_R_X49Y104_SLICE_X75Y104_BQ;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_B1 = 1'b1;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_B2 = 1'b1;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_B3 = 1'b1;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_B4 = 1'b1;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_B5 = 1'b1;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_B6 = 1'b1;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_BX = CLBLM_R_X49Y106_SLICE_X75Y106_DQ;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_C1 = 1'b1;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_C2 = 1'b1;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_C3 = 1'b1;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_C4 = 1'b1;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_C5 = 1'b1;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_C6 = 1'b1;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_CE = CLBLM_L_X62Y101_SLICE_X93Y101_AO6;
  assign CLBLM_L_X64Y108_SLICE_X97Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_CX = CLBLM_R_X49Y107_SLICE_X75Y107_CQ;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_D1 = 1'b1;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_D2 = 1'b1;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_D3 = 1'b1;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_D4 = 1'b1;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_D5 = 1'b1;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_D6 = 1'b1;
  assign CLBLM_L_X62Y101_SLICE_X93Y101_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_A1 = CLBLM_L_X60Y103_SLICE_X90Y103_F8MUX_O;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_A2 = CLBLM_R_X63Y97_SLICE_X94Y97_F7AMUX_O;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_A3 = CLBLM_R_X59Y102_SLICE_X89Y102_AQ;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_A4 = CLBLM_L_X62Y106_SLICE_X93Y106_AQ;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_A5 = 1'b1;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_A6 = CLBLM_L_X60Y110_SLICE_X91Y110_AQ;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_B1 = CLBLM_L_X60Y99_SLICE_X90Y99_BO5;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_B2 = CLBLM_L_X62Y104_SLICE_X92Y104_DO6;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_B3 = CLBLM_L_X62Y96_SLICE_X92Y96_F7AMUX_O;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_B4 = CLBLM_R_X59Y105_SLICE_X88Y105_F7AMUX_O;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_B5 = 1'b1;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_B6 = CLBLM_L_X62Y103_SLICE_X93Y103_BO6;
  assign CLBLM_L_X64Y108_SLICE_X97Y108_D2 = 1'b1;
  assign CLBLM_L_X64Y108_SLICE_X97Y108_D3 = 1'b1;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_C1 = 1'b1;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_C2 = CLBLM_L_X62Y96_SLICE_X93Y96_F7AMUX_O;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_C3 = CLBLM_L_X60Y99_SLICE_X90Y99_BO5;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_C4 = CLBLM_R_X59Y104_SLICE_X89Y104_F7AMUX_O;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_C5 = CLBLM_L_X62Y106_SLICE_X93Y106_DO6;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_C6 = CLBLM_L_X62Y103_SLICE_X93Y103_BO6;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_CE = CLBLM_L_X62Y99_SLICE_X92Y99_DO6;
  assign CLBLM_L_X64Y108_SLICE_X97Y108_D4 = 1'b1;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X64Y108_SLICE_X97Y108_D5 = 1'b1;
  assign CLBLM_L_X64Y108_SLICE_X97Y108_D6 = 1'b1;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_D1 = CLBLM_L_X62Y101_SLICE_X92Y101_BQ;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_D2 = CLBLM_L_X62Y99_SLICE_X92Y99_BQ;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_D3 = CLBLM_L_X62Y101_SLICE_X92Y101_AQ;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_D5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_D6 = 1'b1;
  assign CLBLM_L_X62Y101_SLICE_X92Y101_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X56Y103_SLICE_X84Y103_D2 = 1'b1;
  assign CLBLM_L_X56Y103_SLICE_X84Y103_D3 = CLBLM_L_X56Y103_SLICE_X84Y103_DQ;
  assign CLBLM_L_X56Y103_SLICE_X84Y103_D4 = 1'b1;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_A1 = CLBLM_L_X62Y110_SLICE_X92Y110_DO6;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_A2 = CLBLM_R_X59Y102_SLICE_X89Y102_AQ;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_A3 = CLBLM_L_X62Y103_SLICE_X92Y103_AQ;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_A4 = CLBLM_L_X60Y110_SLICE_X91Y110_AQ;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_A5 = CLBLM_L_X62Y106_SLICE_X93Y106_AQ;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_A6 = 1'b1;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_B1 = 1'b1;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_B2 = 1'b1;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_B3 = 1'b1;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_B4 = 1'b1;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_B5 = 1'b1;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_B6 = 1'b1;
  assign CLBLM_L_X64Y108_SLICE_X96Y108_D3 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X64Y108_SLICE_X96Y108_D4 = CLBLM_L_X62Y105_SLICE_X92Y105_BO5;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_C1 = 1'b1;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_C2 = 1'b1;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_C3 = 1'b1;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_C4 = 1'b1;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_C5 = 1'b1;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_C6 = 1'b1;
  assign CLBLM_L_X64Y108_SLICE_X96Y108_D5 = CLBLM_L_X64Y108_SLICE_X96Y108_BQ;
  assign CLBLM_L_X64Y108_SLICE_X96Y108_D6 = CLBLM_R_X63Y108_SLICE_X95Y108_C_XOR;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_D1 = 1'b1;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_D2 = 1'b1;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_D3 = 1'b1;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_D4 = 1'b1;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_D5 = 1'b1;
  assign CLBLM_L_X62Y102_SLICE_X93Y102_D6 = 1'b1;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_A1 = CLBLM_L_X50Y106_SLICE_X76Y106_AQ;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_A2 = 1'b1;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_A3 = CLBLM_R_X49Y104_SLICE_X75Y104_DQ;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_A4 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_A5 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_A6 = 1'b1;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_B1 = 1'b1;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_B2 = CLBLM_L_X62Y102_SLICE_X92Y102_BQ;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_B3 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_B4 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_B5 = CLBLM_R_X49Y104_SLICE_X74Y104_AQ;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_B6 = CLBLM_L_X50Y104_SLICE_X76Y104_AQ;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_C1 = CLBLM_L_X60Y99_SLICE_X90Y99_AO6;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_C2 = CLBLM_L_X62Y102_SLICE_X93Y102_AO6;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_C3 = CLBLM_L_X62Y104_SLICE_X93Y104_AQ;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_C4 = CLBLL_R_X57Y101_SLICE_X86Y101_AO5;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_C5 = CLBLM_L_X62Y99_SLICE_X92Y99_AO6;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_C6 = CLBLM_L_X60Y101_SLICE_X90Y101_BO6;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_CE = CLBLM_L_X62Y102_SLICE_X92Y102_DO6;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_D1 = CLBLM_L_X60Y100_SLICE_X91Y100_AO6;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_D2 = CLBLM_L_X62Y102_SLICE_X93Y102_AO6;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_D3 = 1'b1;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_D4 = CLBLM_L_X62Y104_SLICE_X93Y104_AQ;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_D5 = CLBLM_L_X62Y99_SLICE_X92Y99_AO6;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_D6 = CLBLM_L_X60Y101_SLICE_X90Y101_BO6;
  assign CLBLM_L_X62Y102_SLICE_X92Y102_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_A1 = CLBLM_R_X63Y110_SLICE_X94Y110_CO6;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_A2 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_A3 = CLBLM_L_X50Y105_SLICE_X77Y105_AQ;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_A4 = CLBLM_R_X49Y104_SLICE_X75Y104_AQ;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_A5 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_A6 = 1'b1;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_B1 = CLBLM_L_X60Y110_SLICE_X91Y110_AQ;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_B2 = CLBLM_L_X62Y104_SLICE_X93Y104_AQ;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_B3 = CLBLM_R_X59Y102_SLICE_X88Y102_AQ;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_B4 = CLBLM_R_X59Y102_SLICE_X89Y102_AQ;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_B5 = CLBLM_L_X62Y103_SLICE_X92Y103_AQ;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_B6 = 1'b1;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_C1 = 1'b1;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_C2 = 1'b1;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_C3 = 1'b1;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_C4 = 1'b1;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_C5 = 1'b1;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_C6 = 1'b1;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_CE = CLBLM_L_X62Y100_SLICE_X92Y100_DO6;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_D1 = 1'b1;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_D2 = 1'b1;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_D3 = 1'b1;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_D4 = 1'b1;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_D5 = 1'b1;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_D6 = 1'b1;
  assign CLBLM_L_X62Y103_SLICE_X93Y103_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_A1 = 1'b1;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_A2 = CLBLM_R_X49Y104_SLICE_X75Y104_BQ;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_A3 = CLBLM_L_X60Y108_SLICE_X91Y108_BO6;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_A4 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_A5 = CLBLM_L_X62Y103_SLICE_X92Y103_CO6;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_A6 = CLBLM_R_X59Y103_SLICE_X89Y103_DQ;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_B1 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_B2 = CLBLM_R_X59Y103_SLICE_X89Y103_CQ;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_B3 = CLBLM_L_X60Y102_SLICE_X91Y102_BQ;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_B4 = CLBLM_R_X59Y103_SLICE_X89Y103_DQ;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_B5 = CLBLM_L_X60Y103_SLICE_X91Y103_AQ;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_B6 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_C1 = CLBLM_L_X62Y104_SLICE_X92Y104_AQ;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_C2 = CLBLM_R_X59Y103_SLICE_X89Y103_CQ;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_C3 = CLBLM_L_X60Y105_SLICE_X91Y105_B_XOR;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_C4 = CLBLM_L_X60Y101_SLICE_X90Y101_CO6;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_C5 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_C6 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_CE = CLBLM_R_X59Y99_SLICE_X89Y99_CO6;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_D1 = 1'b1;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_D2 = 1'b1;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_D3 = 1'b1;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_D4 = 1'b1;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_D5 = 1'b1;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_D6 = 1'b1;
  assign CLBLM_L_X62Y103_SLICE_X92Y103_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_D = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_D = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X62Y104_SLICE_X93Y104_A1 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y104_SLICE_X93Y104_A2 = CLBLM_R_X49Y104_SLICE_X75Y104_AQ;
  assign CLBLM_L_X62Y104_SLICE_X93Y104_A3 = CLBLM_R_X59Y107_SLICE_X88Y107_AO6;
  assign CLBLM_L_X62Y104_SLICE_X93Y104_A4 = CLBLM_L_X60Y104_SLICE_X90Y104_BO6;
  assign CLBLM_L_X62Y104_SLICE_X93Y104_A5 = CLBLM_R_X59Y103_SLICE_X89Y103_DQ;
  assign CLBLM_L_X62Y104_SLICE_X93Y104_A6 = 1'b1;
  assign CLBLM_L_X62Y104_SLICE_X93Y104_B1 = 1'b1;
  assign CLBLM_L_X62Y104_SLICE_X93Y104_B2 = 1'b1;
  assign CLBLM_L_X62Y104_SLICE_X93Y104_B3 = 1'b1;
  assign CLBLM_L_X62Y104_SLICE_X93Y104_B4 = 1'b1;
  assign CLBLM_L_X62Y104_SLICE_X93Y104_B5 = 1'b1;
  assign CLBLM_L_X62Y104_SLICE_X93Y104_B6 = 1'b1;
  assign CLBLM_L_X62Y104_SLICE_X93Y104_C1 = 1'b1;
  assign CLBLM_L_X62Y104_SLICE_X93Y104_C2 = 1'b1;
  assign CLBLM_L_X62Y104_SLICE_X93Y104_C3 = 1'b1;
  assign CLBLM_L_X62Y104_SLICE_X93Y104_C4 = 1'b1;
  assign CLBLM_L_X62Y104_SLICE_X93Y104_C5 = 1'b1;
  assign CLBLM_L_X62Y104_SLICE_X93Y104_C6 = 1'b1;
  assign CLBLM_L_X62Y104_SLICE_X93Y104_CE = CLBLM_R_X59Y99_SLICE_X89Y99_CO6;
  assign CLBLM_L_X62Y104_SLICE_X93Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X62Y104_SLICE_X93Y104_D1 = 1'b1;
  assign CLBLM_L_X62Y104_SLICE_X93Y104_D2 = 1'b1;
  assign CLBLM_L_X62Y104_SLICE_X93Y104_D3 = 1'b1;
  assign CLBLM_L_X62Y104_SLICE_X93Y104_D4 = 1'b1;
  assign CLBLM_L_X62Y104_SLICE_X93Y104_D5 = 1'b1;
  assign CLBLM_L_X62Y104_SLICE_X93Y104_D6 = 1'b1;
  assign CLBLM_L_X62Y104_SLICE_X93Y104_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X62Y104_SLICE_X92Y104_A1 = CLBLM_L_X60Y102_SLICE_X91Y102_B_XOR;
  assign CLBLM_L_X62Y104_SLICE_X92Y104_A2 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X62Y104_SLICE_X92Y104_A3 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X62Y104_SLICE_X92Y104_A4 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y104_SLICE_X92Y104_A5 = CLBLM_L_X62Y105_SLICE_X92Y105_AO6;
  assign CLBLM_L_X62Y104_SLICE_X92Y104_A6 = CLBLM_L_X60Y105_SLICE_X91Y105_B_XOR;
  assign CLBLM_L_X62Y104_SLICE_X92Y104_B1 = CLBLM_L_X62Y106_SLICE_X93Y106_BO5;
  assign CLBLM_L_X62Y104_SLICE_X92Y104_B2 = CLBLM_L_X60Y103_SLICE_X91Y103_A_XOR;
  assign CLBLM_L_X62Y104_SLICE_X92Y104_B3 = CLBLM_L_X60Y106_SLICE_X91Y106_A_XOR;
  assign CLBLM_L_X62Y104_SLICE_X92Y104_B4 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X62Y104_SLICE_X92Y104_B5 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X62Y104_SLICE_X92Y104_B6 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y104_SLICE_X92Y104_C1 = CLBLM_L_X60Y104_SLICE_X91Y104_AQ;
  assign CLBLM_L_X62Y104_SLICE_X92Y104_C2 = CLBLM_R_X59Y103_SLICE_X89Y103_DQ;
  assign CLBLM_L_X62Y104_SLICE_X92Y104_C3 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X62Y104_SLICE_X92Y104_C4 = CLBLM_R_X59Y103_SLICE_X89Y103_CQ;
  assign CLBLM_L_X62Y104_SLICE_X92Y104_C5 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_L_X62Y104_SLICE_X92Y104_C6 = CLBLM_R_X59Y99_SLICE_X88Y99_BQ;
  assign CLBLM_L_X62Y104_SLICE_X92Y104_CE = CLBLM_L_X62Y102_SLICE_X92Y102_DO6;
  assign CLBLM_L_X62Y104_SLICE_X92Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X62Y104_SLICE_X92Y104_D1 = CLBLM_L_X62Y104_SLICE_X92Y104_BQ;
  assign CLBLM_L_X62Y104_SLICE_X92Y104_D2 = CLBLM_L_X60Y104_SLICE_X90Y104_CO6;
  assign CLBLM_L_X62Y104_SLICE_X92Y104_D3 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_L_X62Y104_SLICE_X92Y104_D4 = CLBLM_L_X62Y106_SLICE_X93Y106_CO6;
  assign CLBLM_L_X62Y104_SLICE_X92Y104_D5 = CLBLM_L_X62Y107_SLICE_X92Y107_A5Q;
  assign CLBLM_L_X62Y104_SLICE_X92Y104_D6 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_L_X62Y104_SLICE_X92Y104_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_A1 = CLBLM_R_X63Y105_SLICE_X94Y105_A_XOR;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_A2 = CLBLM_L_X62Y105_SLICE_X92Y105_CQ;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_A3 = CLBLM_R_X59Y103_SLICE_X89Y103_A5Q;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_A4 = CLBLM_R_X59Y101_SLICE_X89Y101_AQ;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_A5 = CLBLL_R_X57Y102_SLICE_X86Y102_AQ;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_A6 = 1'b1;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_B1 = CLBLM_R_X63Y106_SLICE_X95Y106_A_XOR;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_B2 = CLBLM_L_X62Y105_SLICE_X93Y105_BQ;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_B3 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_B4 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_B5 = CLBLM_L_X62Y105_SLICE_X92Y105_BO5;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_B6 = CLBLM_L_X62Y105_SLICE_X93Y105_CO6;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_C1 = CLBLM_L_X62Y105_SLICE_X93Y105_AO6;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_C2 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_C3 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_C4 = CLBLM_R_X63Y106_SLICE_X95Y106_A_XOR;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_C5 = CLBLM_R_X63Y106_SLICE_X94Y106_B_XOR;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_C6 = CLBLM_L_X50Y106_SLICE_X76Y106_CQ;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_CE = CLBLM_L_X62Y100_SLICE_X92Y100_CO6;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_D1 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_D2 = CLBLM_R_X49Y119_SLICE_X74Y119_BQ;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_D3 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_D4 = CLBLM_L_X62Y105_SLICE_X92Y105_BO6;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_D5 = CLBLM_R_X49Y119_SLICE_X74Y119_AQ;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_D6 = 1'b1;
  assign CLBLM_L_X62Y105_SLICE_X93Y105_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_A1 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_A2 = CLBLM_R_X49Y105_SLICE_X75Y105_CQ;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_A3 = CLBLM_R_X49Y104_SLICE_X75Y104_BQ;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_A4 = CLBLM_L_X64Y109_SLICE_X96Y109_CO6;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_A5 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_A6 = 1'b1;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_B1 = CLBLM_R_X59Y101_SLICE_X89Y101_AQ;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_B2 = CLBLL_R_X57Y102_SLICE_X86Y102_BQ;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_B3 = CLBLL_R_X57Y102_SLICE_X86Y102_AQ;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_B4 = CLBLM_R_X59Y103_SLICE_X89Y103_A5Q;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_B5 = 1'b1;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_B6 = 1'b1;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_C1 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_C2 = CLBLM_L_X62Y105_SLICE_X93Y105_AO5;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_C3 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_C4 = CLBLM_L_X50Y104_SLICE_X76Y104_AQ;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_C5 = CLBLM_L_X62Y105_SLICE_X92Y105_BO5;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_C6 = CLBLM_L_X62Y105_SLICE_X92Y105_CQ;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_CE = CLBLM_L_X62Y100_SLICE_X92Y100_CO6;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_D1 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_D2 = CLBLM_L_X62Y106_SLICE_X93Y106_CO6;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_D3 = CLBLM_L_X60Y108_SLICE_X90Y108_BQ;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_D4 = CLBLM_R_X59Y105_SLICE_X89Y105_DO6;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_D5 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_D6 = CLBLM_L_X62Y106_SLICE_X92Y106_BQ;
  assign CLBLM_L_X62Y105_SLICE_X92Y105_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLL_R_X57Y111_SLICE_X86Y111_A3 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X86Y111_B3 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X86Y111_C5 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X86Y111_C6 = 1'b1;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_A1 = CLBLM_R_X59Y103_SLICE_X89Y103_DQ;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_A2 = CLBLM_R_X59Y110_SLICE_X89Y110_CO6;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_A3 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_A4 = CLBLM_L_X62Y106_SLICE_X92Y106_DO6;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_A5 = CLBLM_R_X49Y106_SLICE_X75Y106_CQ;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_A6 = 1'b1;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_B1 = 1'b1;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_B2 = CLBLM_L_X50Y106_SLICE_X76Y106_CQ;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_B3 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_B4 = CLBLM_R_X49Y106_SLICE_X75Y106_CQ;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_B5 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_B6 = 1'b1;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_D = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_C1 = CLBLM_L_X62Y104_SLICE_X93Y104_AQ;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_C2 = CLBLM_L_X60Y110_SLICE_X91Y110_AQ;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_C3 = CLBLM_R_X59Y102_SLICE_X88Y102_AQ;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_C4 = CLBLM_R_X59Y102_SLICE_X89Y102_AQ;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_C5 = CLBLM_L_X62Y106_SLICE_X93Y106_AQ;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_C6 = CLBLM_L_X62Y103_SLICE_X92Y103_AQ;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_CE = CLBLM_R_X59Y99_SLICE_X89Y99_CO6;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_D = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_D1 = CLBLM_L_X62Y106_SLICE_X93Y106_CO6;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_D2 = CLBLM_L_X62Y107_SLICE_X92Y107_DO6;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_D3 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_D4 = CLBLM_L_X62Y106_SLICE_X92Y106_CQ;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_D5 = CLBLM_L_X62Y107_SLICE_X92Y107_BQ;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_D6 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_L_X62Y106_SLICE_X93Y106_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_A1 = CLBLM_L_X60Y106_SLICE_X90Y106_B_XOR;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_A2 = CLBLM_R_X59Y112_SLICE_X89Y112_AQ;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_A3 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_A4 = CLBLM_R_X59Y103_SLICE_X89Y103_CQ;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_A5 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_A6 = 1'b1;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_B1 = CLBLM_L_X62Y108_SLICE_X92Y108_BO5;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_B2 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_B3 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_B4 = CLBLM_L_X60Y106_SLICE_X91Y106_B_XOR;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_B5 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_B6 = CLBLM_L_X60Y103_SLICE_X91Y103_B_XOR;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_C1 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_C2 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_C3 = CLBLM_L_X62Y107_SLICE_X92Y107_BO5;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_C4 = CLBLM_L_X60Y103_SLICE_X91Y103_C_XOR;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_C5 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_C6 = CLBLM_L_X60Y106_SLICE_X91Y106_C_XOR;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_CE = CLBLM_L_X62Y102_SLICE_X92Y102_DO6;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X64Y109_SLICE_X97Y109_D4 = 1'b1;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_D1 = CLBLM_L_X62Y106_SLICE_X92Y106_AO6;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_D2 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_D3 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X64Y109_SLICE_X97Y109_D5 = 1'b1;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_D4 = CLBLM_L_X60Y106_SLICE_X91Y106_A_XOR;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_D5 = CLBLM_L_X62Y104_SLICE_X92Y104_BQ;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_D6 = CLBLM_R_X59Y103_SLICE_X89Y103_CQ;
  assign CLBLM_L_X64Y109_SLICE_X97Y109_D6 = 1'b1;
  assign CLBLM_L_X62Y106_SLICE_X92Y106_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X56Y104_SLICE_X84Y104_CX = 1'b0;
  assign CLBLM_L_X56Y104_SLICE_X84Y104_D1 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X84Y104_D2 = 1'b1;
  assign CLBLM_L_X64Y109_SLICE_X96Y109_A6 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X84Y104_DX = 1'b0;
  assign CLBLM_L_X56Y104_SLICE_X84Y104_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X64Y109_SLICE_X96Y109_B5 = CLBLM_L_X62Y105_SLICE_X92Y105_BO5;
  assign CLBLM_L_X64Y109_SLICE_X96Y109_B6 = CLBLM_R_X63Y108_SLICE_X95Y108_D_XOR;
  assign CLBLM_L_X64Y109_SLICE_X96Y109_C5 = CLBLM_R_X63Y109_SLICE_X94Y109_C_XOR;
  assign CLBLM_L_X64Y109_SLICE_X96Y109_C6 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X64Y109_SLICE_X96Y109_CE = CLBLM_L_X62Y100_SLICE_X92Y100_DO6;
  assign CLBLM_L_X64Y109_SLICE_X96Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_A1 = CLBLM_L_X60Y110_SLICE_X91Y110_AQ;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_A2 = CLBLM_R_X59Y102_SLICE_X89Y102_AQ;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_A3 = CLBLM_L_X62Y106_SLICE_X93Y106_AQ;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_A4 = CLBLM_L_X62Y104_SLICE_X93Y104_AQ;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_A5 = CLBLM_L_X62Y103_SLICE_X92Y103_AQ;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_A6 = CLBLM_R_X59Y102_SLICE_X88Y102_AQ;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_B1 = CLBLM_L_X60Y110_SLICE_X91Y110_AQ;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_B2 = CLBLM_R_X59Y102_SLICE_X89Y102_AQ;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_B3 = CLBLM_L_X62Y106_SLICE_X93Y106_AQ;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_B4 = CLBLM_L_X62Y104_SLICE_X93Y104_AQ;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_B5 = CLBLM_L_X62Y103_SLICE_X92Y103_AQ;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_B6 = CLBLM_R_X59Y102_SLICE_X88Y102_AQ;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_C1 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_C2 = CLBLM_L_X64Y105_SLICE_X97Y105_AQ;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_C3 = 1'b1;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_C4 = CLBLM_R_X49Y111_SLICE_X74Y111_BQ;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_C5 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_C6 = CLBLM_L_X64Y107_SLICE_X97Y107_AQ;
  assign CLBLM_L_X64Y109_SLICE_X96Y109_D4 = CLBLM_L_X64Y109_SLICE_X96Y109_A5Q;
  assign CLBLM_L_X64Y109_SLICE_X96Y109_D5 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_D1 = 1'b1;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_D2 = 1'b1;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_D3 = 1'b1;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_D4 = 1'b1;
  assign CLBLM_L_X64Y109_SLICE_X96Y109_D6 = CLBLM_R_X63Y109_SLICE_X95Y109_C_XOR;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_D6 = 1'b1;
  assign CLBLM_L_X62Y107_SLICE_X93Y107_D5 = 1'b1;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_A1 = CLBLM_L_X60Y107_SLICE_X91Y107_B_XOR;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_A2 = CLBLM_L_X62Y100_SLICE_X93Y100_AO6;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_A3 = CLBLM_L_X60Y104_SLICE_X91Y104_B_XOR;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_A4 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_A5 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_A6 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_AX = CLBLM_L_X62Y106_SLICE_X93Y106_BO6;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_B1 = CLBLM_R_X49Y107_SLICE_X75Y107_CQ;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_B2 = CLBLM_L_X50Y107_SLICE_X77Y107_AQ;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_B3 = 1'b1;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_B4 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_B5 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_B6 = 1'b1;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_C1 = CLBLM_L_X60Y106_SLICE_X90Y106_AQ;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_C2 = CLBLM_R_X59Y103_SLICE_X89Y103_CQ;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_C3 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_C4 = CLBLM_L_X62Y107_SLICE_X92Y107_A5Q;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_C5 = CLBLM_R_X59Y103_SLICE_X89Y103_DQ;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_C6 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_CE = CLBLM_L_X62Y102_SLICE_X92Y102_CO6;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X57Y111_SLICE_X87Y111_D5 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X87Y111_D6 = CLBLL_R_X57Y109_SLICE_X86Y109_CQ;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_D1 = CLBLM_L_X60Y107_SLICE_X91Y107_AQ;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_D2 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_D3 = CLBLM_R_X59Y100_SLICE_X89Y100_DQ;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_D4 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_D5 = CLBLM_R_X59Y106_SLICE_X89Y106_BQ;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_D6 = CLBLM_R_X59Y96_SLICE_X89Y96_A5Q;
  assign CLBLM_L_X62Y107_SLICE_X92Y107_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X49Y119_SLICE_X75Y119_A1 = 1'b1;
  assign CLBLM_R_X49Y119_SLICE_X75Y119_A2 = 1'b1;
  assign CLBLM_R_X49Y119_SLICE_X75Y119_A3 = 1'b1;
  assign CLBLM_R_X49Y119_SLICE_X75Y119_A4 = 1'b1;
  assign CLBLM_R_X49Y119_SLICE_X75Y119_A5 = 1'b1;
  assign CLBLM_R_X49Y119_SLICE_X75Y119_A6 = 1'b1;
  assign CLBLM_R_X49Y119_SLICE_X75Y119_B1 = 1'b1;
  assign CLBLM_R_X49Y119_SLICE_X75Y119_B2 = 1'b1;
  assign CLBLM_R_X49Y119_SLICE_X75Y119_B3 = 1'b1;
  assign CLBLM_R_X49Y119_SLICE_X75Y119_B4 = 1'b1;
  assign CLBLM_R_X49Y119_SLICE_X75Y119_B5 = 1'b1;
  assign CLBLM_R_X49Y119_SLICE_X75Y119_B6 = 1'b1;
  assign CLBLM_R_X49Y119_SLICE_X75Y119_C1 = 1'b1;
  assign CLBLM_R_X49Y119_SLICE_X75Y119_C2 = 1'b1;
  assign CLBLM_R_X49Y119_SLICE_X75Y119_C3 = 1'b1;
  assign CLBLM_R_X49Y119_SLICE_X75Y119_C4 = 1'b1;
  assign CLBLM_R_X49Y119_SLICE_X75Y119_C5 = 1'b1;
  assign CLBLM_R_X49Y119_SLICE_X75Y119_C6 = 1'b1;
  assign CLBLM_R_X49Y119_SLICE_X75Y119_D1 = 1'b1;
  assign CLBLM_R_X49Y119_SLICE_X75Y119_D2 = 1'b1;
  assign CLBLM_R_X49Y119_SLICE_X75Y119_D3 = 1'b1;
  assign CLBLM_R_X49Y119_SLICE_X75Y119_D4 = 1'b1;
  assign CLBLM_R_X49Y119_SLICE_X75Y119_D5 = 1'b1;
  assign CLBLM_R_X49Y119_SLICE_X75Y119_D6 = 1'b1;
  assign CLBLM_R_X49Y119_SLICE_X74Y119_A1 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLM_R_X49Y119_SLICE_X74Y119_A2 = CLBLM_R_X49Y119_SLICE_X74Y119_BQ;
  assign CLBLM_R_X49Y119_SLICE_X74Y119_A3 = CLBLM_R_X49Y119_SLICE_X74Y119_AQ;
  assign CLBLM_R_X49Y119_SLICE_X74Y119_A4 = CLBLM_R_X47Y119_SLICE_X73Y119_BO6;
  assign CLBLM_R_X49Y119_SLICE_X74Y119_A5 = CLBLM_R_X47Y119_SLICE_X73Y119_AO6;
  assign CLBLM_R_X49Y119_SLICE_X74Y119_A6 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLM_R_X49Y119_SLICE_X74Y119_B1 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLM_R_X49Y119_SLICE_X74Y119_B2 = CLBLM_R_X49Y119_SLICE_X74Y119_BQ;
  assign CLBLM_R_X49Y119_SLICE_X74Y119_B3 = CLBLM_R_X49Y119_SLICE_X74Y119_AQ;
  assign CLBLM_R_X49Y119_SLICE_X74Y119_B4 = CLBLM_R_X47Y119_SLICE_X73Y119_BO6;
  assign CLBLM_R_X49Y119_SLICE_X74Y119_B5 = CLBLM_L_X56Y102_SLICE_X85Y102_A5Q;
  assign CLBLM_R_X49Y119_SLICE_X74Y119_B6 = CLBLM_R_X47Y119_SLICE_X73Y119_AO5;
  assign CLBLM_R_X49Y119_SLICE_X74Y119_C1 = 1'b1;
  assign CLBLM_R_X49Y119_SLICE_X74Y119_C2 = 1'b1;
  assign CLBLM_R_X49Y119_SLICE_X74Y119_C3 = 1'b1;
  assign CLBLM_R_X49Y119_SLICE_X74Y119_C4 = 1'b1;
  assign CLBLM_R_X49Y119_SLICE_X74Y119_C5 = 1'b1;
  assign CLBLM_R_X49Y119_SLICE_X74Y119_C6 = 1'b1;
  assign CLBLM_R_X49Y119_SLICE_X74Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X49Y119_SLICE_X74Y119_D1 = 1'b1;
  assign CLBLM_R_X49Y119_SLICE_X74Y119_D2 = 1'b1;
  assign CLBLM_R_X49Y119_SLICE_X74Y119_D3 = 1'b1;
  assign CLBLM_R_X49Y119_SLICE_X74Y119_D4 = 1'b1;
  assign CLBLM_R_X49Y119_SLICE_X74Y119_D5 = 1'b1;
  assign CLBLM_R_X49Y119_SLICE_X74Y119_D6 = 1'b1;
  assign CLBLM_R_X49Y119_SLICE_X74Y119_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_D1 = CLBLM_R_X63Y103_SLICE_X95Y103_BQ;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_D1 = CLBLM_R_X65Y106_SLICE_X98Y106_DQ;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_T1 = 1'b1;
  assign CLBLM_L_X62Y108_SLICE_X93Y108_A1 = CLBLM_R_X59Y107_SLICE_X88Y107_CO6;
  assign CLBLM_L_X62Y108_SLICE_X93Y108_A2 = CLBLM_R_X59Y103_SLICE_X89Y103_DQ;
  assign CLBLM_L_X62Y108_SLICE_X93Y108_A3 = CLBLM_R_X49Y107_SLICE_X75Y107_CQ;
  assign CLBLM_L_X62Y108_SLICE_X93Y108_A4 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y108_SLICE_X93Y108_A5 = 1'b1;
  assign CLBLM_L_X62Y108_SLICE_X93Y108_A6 = CLBLM_L_X62Y108_SLICE_X93Y108_CO6;
  assign CLBLM_L_X62Y108_SLICE_X93Y108_B1 = CLBLM_R_X59Y103_SLICE_X89Y103_DQ;
  assign CLBLM_L_X62Y108_SLICE_X93Y108_B2 = CLBLM_R_X59Y103_SLICE_X89Y103_CQ;
  assign CLBLM_L_X62Y108_SLICE_X93Y108_B3 = CLBLM_L_X62Y107_SLICE_X92Y107_BQ;
  assign CLBLM_L_X62Y108_SLICE_X93Y108_B4 = CLBLM_L_X60Y107_SLICE_X91Y107_AQ;
  assign CLBLM_L_X62Y108_SLICE_X93Y108_B5 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_L_X62Y108_SLICE_X93Y108_B6 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X62Y108_SLICE_X93Y108_C1 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_L_X62Y108_SLICE_X93Y108_C2 = CLBLM_L_X62Y106_SLICE_X92Y106_CQ;
  assign CLBLM_L_X62Y108_SLICE_X93Y108_C3 = CLBLM_R_X59Y103_SLICE_X89Y103_CQ;
  assign CLBLM_L_X62Y108_SLICE_X93Y108_C4 = CLBLM_L_X60Y106_SLICE_X91Y106_C_XOR;
  assign CLBLM_L_X62Y108_SLICE_X93Y108_C5 = CLBLM_L_X62Y108_SLICE_X93Y108_DO6;
  assign CLBLM_L_X62Y108_SLICE_X93Y108_C6 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X62Y108_SLICE_X93Y108_CE = CLBLM_R_X59Y99_SLICE_X89Y99_CO6;
  assign CLBLM_L_X62Y108_SLICE_X93Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X62Y108_SLICE_X93Y108_D1 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_L_X62Y108_SLICE_X93Y108_D2 = CLBLM_R_X59Y106_SLICE_X89Y106_BQ;
  assign CLBLM_L_X62Y108_SLICE_X93Y108_D3 = 1'b1;
  assign CLBLM_L_X62Y108_SLICE_X93Y108_D4 = CLBLM_L_X60Y106_SLICE_X90Y106_D_XOR;
  assign CLBLM_L_X62Y108_SLICE_X93Y108_D5 = 1'b1;
  assign CLBLM_L_X62Y108_SLICE_X93Y108_D6 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X62Y108_SLICE_X93Y108_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X62Y108_SLICE_X92Y108_A1 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y108_SLICE_X92Y108_A2 = CLBLM_R_X59Y105_SLICE_X88Y105_CO6;
  assign CLBLM_L_X62Y108_SLICE_X92Y108_A3 = CLBLM_L_X62Y107_SLICE_X92Y107_CO6;
  assign CLBLM_L_X62Y108_SLICE_X92Y108_A4 = CLBLM_L_X62Y103_SLICE_X92Y103_BO6;
  assign CLBLM_L_X62Y108_SLICE_X92Y108_A5 = CLBLM_L_X62Y104_SLICE_X92Y104_CO6;
  assign CLBLM_L_X62Y108_SLICE_X92Y108_A6 = 1'b1;
  assign CLBLM_L_X62Y108_SLICE_X92Y108_B1 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y108_SLICE_X92Y108_B2 = 1'b1;
  assign CLBLM_L_X62Y108_SLICE_X92Y108_B3 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X62Y108_SLICE_X92Y108_B4 = CLBLM_R_X49Y106_SLICE_X75Y106_DQ;
  assign CLBLM_L_X62Y108_SLICE_X92Y108_B5 = CLBLM_L_X50Y107_SLICE_X76Y107_BQ;
  assign CLBLM_L_X62Y108_SLICE_X92Y108_B6 = 1'b1;
  assign CLBLL_R_X57Y97_SLICE_X86Y97_A1 = CLBLL_R_X57Y97_SLICE_X86Y97_BO6;
  assign CLBLL_R_X57Y97_SLICE_X86Y97_A2 = CLBLM_L_X60Y99_SLICE_X91Y99_DO6;
  assign CLBLL_R_X57Y97_SLICE_X86Y97_A3 = CLBLL_R_X57Y97_SLICE_X86Y97_AQ;
  assign CLBLL_R_X57Y97_SLICE_X86Y97_A4 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLL_R_X57Y97_SLICE_X86Y97_A5 = CLBLM_L_X50Y104_SLICE_X76Y104_AQ;
  assign CLBLL_R_X57Y97_SLICE_X86Y97_A6 = CLBLL_R_X57Y98_SLICE_X86Y98_AO6;
  assign CLBLM_L_X62Y108_SLICE_X92Y108_C1 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_L_X62Y108_SLICE_X92Y108_C2 = CLBLM_L_X60Y108_SLICE_X90Y108_BQ;
  assign CLBLL_R_X57Y97_SLICE_X86Y97_B1 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLL_R_X57Y97_SLICE_X86Y97_B2 = CLBLL_R_X57Y97_SLICE_X86Y97_CO6;
  assign CLBLL_R_X57Y97_SLICE_X86Y97_B3 = CLBLL_R_X57Y97_SLICE_X86Y97_AQ;
  assign CLBLL_R_X57Y97_SLICE_X86Y97_B4 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLL_R_X57Y97_SLICE_X86Y97_B5 = CLBLL_R_X57Y97_SLICE_X87Y97_AQ;
  assign CLBLL_R_X57Y97_SLICE_X86Y97_B6 = CLBLM_L_X50Y105_SLICE_X76Y105_AQ;
  assign CLBLM_L_X62Y108_SLICE_X92Y108_C6 = CLBLM_R_X59Y103_SLICE_X89Y103_DQ;
  assign CLBLM_L_X62Y108_SLICE_X92Y108_CE = CLBLM_R_X59Y99_SLICE_X89Y99_CO6;
  assign CLBLM_L_X62Y108_SLICE_X92Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X57Y97_SLICE_X86Y97_C1 = 1'b1;
  assign CLBLL_R_X57Y97_SLICE_X86Y97_C2 = 1'b1;
  assign CLBLL_R_X57Y97_SLICE_X86Y97_C3 = 1'b1;
  assign CLBLL_R_X57Y97_SLICE_X86Y97_C4 = CLBLM_L_X56Y98_SLICE_X85Y98_CQ;
  assign CLBLL_R_X57Y97_SLICE_X86Y97_C5 = 1'b1;
  assign CLBLL_R_X57Y97_SLICE_X86Y97_C6 = CLBLM_L_X56Y98_SLICE_X85Y98_BQ;
  assign CLBLM_L_X62Y108_SLICE_X92Y108_D1 = 1'b1;
  assign CLBLM_L_X62Y108_SLICE_X92Y108_D2 = 1'b1;
  assign CLBLL_R_X57Y97_SLICE_X86Y97_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X62Y108_SLICE_X92Y108_D3 = 1'b1;
  assign CLBLM_L_X62Y108_SLICE_X92Y108_D4 = 1'b1;
  assign CLBLM_L_X62Y108_SLICE_X92Y108_D5 = 1'b1;
  assign CLBLM_L_X62Y108_SLICE_X92Y108_D6 = 1'b1;
  assign CLBLL_R_X57Y97_SLICE_X86Y97_D1 = 1'b1;
  assign CLBLL_R_X57Y97_SLICE_X86Y97_D2 = 1'b1;
  assign CLBLL_R_X57Y97_SLICE_X86Y97_D3 = 1'b1;
  assign CLBLL_R_X57Y97_SLICE_X86Y97_D4 = 1'b1;
  assign CLBLL_R_X57Y97_SLICE_X86Y97_D5 = 1'b1;
  assign CLBLL_R_X57Y97_SLICE_X86Y97_D6 = 1'b1;
  assign CLBLL_R_X57Y97_SLICE_X86Y97_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_D = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_D = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_R_X57Y97_SLICE_X87Y97_A1 = CLBLM_L_X60Y98_SLICE_X91Y98_DQ;
  assign CLBLL_R_X57Y97_SLICE_X87Y97_A2 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLL_R_X57Y97_SLICE_X87Y97_A3 = 1'b1;
  assign CLBLL_R_X57Y97_SLICE_X87Y97_A4 = CLBLM_L_X56Y98_SLICE_X85Y98_BQ;
  assign CLBLL_R_X57Y97_SLICE_X87Y97_A5 = 1'b1;
  assign CLBLL_R_X57Y97_SLICE_X87Y97_A6 = CLBLM_L_X56Y98_SLICE_X85Y98_CQ;
  assign CLBLL_R_X57Y97_SLICE_X87Y97_AX = CLBLL_R_X57Y97_SLICE_X86Y97_AQ;
  assign CLBLL_R_X57Y97_SLICE_X87Y97_B1 = 1'b1;
  assign CLBLL_R_X57Y97_SLICE_X87Y97_B2 = 1'b1;
  assign CLBLL_R_X57Y97_SLICE_X87Y97_B3 = 1'b1;
  assign CLBLL_R_X57Y97_SLICE_X87Y97_B4 = 1'b1;
  assign CLBLL_R_X57Y97_SLICE_X87Y97_B5 = 1'b1;
  assign CLBLL_R_X57Y97_SLICE_X87Y97_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_R_X57Y97_SLICE_X87Y97_C1 = 1'b1;
  assign CLBLL_R_X57Y97_SLICE_X87Y97_C2 = 1'b1;
  assign CLBLL_R_X57Y97_SLICE_X87Y97_C3 = 1'b1;
  assign CLBLL_R_X57Y97_SLICE_X87Y97_C4 = 1'b1;
  assign CLBLL_R_X57Y97_SLICE_X87Y97_C5 = 1'b1;
  assign CLBLL_R_X57Y97_SLICE_X87Y97_C6 = 1'b1;
  assign CLBLL_R_X57Y97_SLICE_X87Y97_CE = CLBLL_R_X57Y97_SLICE_X87Y97_AO6;
  assign CLBLL_R_X57Y97_SLICE_X87Y97_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLL_R_X57Y97_SLICE_X87Y97_D1 = 1'b1;
  assign CLBLL_R_X57Y97_SLICE_X87Y97_D2 = 1'b1;
  assign CLBLL_R_X57Y97_SLICE_X87Y97_D3 = 1'b1;
  assign CLBLL_R_X57Y97_SLICE_X87Y97_D4 = 1'b1;
  assign CLBLL_R_X57Y97_SLICE_X87Y97_D5 = 1'b1;
  assign CLBLL_R_X57Y97_SLICE_X87Y97_D6 = 1'b1;
  assign CLBLL_R_X57Y97_SLICE_X87Y97_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X62Y109_SLICE_X93Y109_A1 = 1'b1;
  assign CLBLM_L_X62Y109_SLICE_X93Y109_A2 = 1'b1;
  assign CLBLM_L_X62Y109_SLICE_X93Y109_A3 = 1'b1;
  assign CLBLM_L_X62Y109_SLICE_X93Y109_A4 = 1'b1;
  assign CLBLM_L_X62Y109_SLICE_X93Y109_A5 = 1'b1;
  assign CLBLM_L_X62Y109_SLICE_X93Y109_A6 = 1'b1;
  assign CLBLM_L_X62Y109_SLICE_X93Y109_B1 = 1'b1;
  assign CLBLM_L_X62Y109_SLICE_X93Y109_B2 = 1'b1;
  assign CLBLM_L_X62Y109_SLICE_X93Y109_B3 = 1'b1;
  assign CLBLM_L_X62Y109_SLICE_X93Y109_B4 = 1'b1;
  assign CLBLM_L_X62Y109_SLICE_X93Y109_B5 = 1'b1;
  assign CLBLM_L_X62Y109_SLICE_X93Y109_B6 = 1'b1;
  assign CLBLM_L_X62Y109_SLICE_X93Y109_C1 = 1'b1;
  assign CLBLM_L_X62Y109_SLICE_X93Y109_C2 = 1'b1;
  assign CLBLM_L_X62Y109_SLICE_X93Y109_C3 = 1'b1;
  assign CLBLM_L_X62Y109_SLICE_X93Y109_C4 = 1'b1;
  assign CLBLM_L_X56Y97_SLICE_X85Y97_A1 = CLBLM_L_X56Y97_SLICE_X85Y97_BO5;
  assign CLBLM_L_X56Y97_SLICE_X85Y97_A2 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLM_L_X56Y97_SLICE_X85Y97_A3 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLM_L_X56Y97_SLICE_X85Y97_A4 = CLBLM_L_X56Y97_SLICE_X85Y97_BO6;
  assign CLBLM_L_X56Y97_SLICE_X85Y97_A5 = CLBLM_R_X49Y108_SLICE_X75Y108_DQ;
  assign CLBLM_L_X56Y97_SLICE_X85Y97_A6 = CLBLM_R_X49Y107_SLICE_X75Y107_DQ;
  assign CLBLM_L_X62Y109_SLICE_X93Y109_C5 = 1'b1;
  assign CLBLM_L_X62Y109_SLICE_X93Y109_C6 = 1'b1;
  assign CLBLM_L_X56Y97_SLICE_X85Y97_B1 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLM_L_X56Y97_SLICE_X85Y97_B2 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign CLBLM_L_X56Y97_SLICE_X85Y97_B3 = 1'b1;
  assign CLBLM_L_X56Y97_SLICE_X85Y97_B4 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLM_L_X56Y97_SLICE_X85Y97_B5 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLM_L_X56Y97_SLICE_X85Y97_B6 = 1'b1;
  assign CLBLM_L_X62Y109_SLICE_X93Y109_D1 = 1'b1;
  assign CLBLM_L_X62Y109_SLICE_X93Y109_D2 = 1'b1;
  assign CLBLM_L_X62Y109_SLICE_X93Y109_D3 = 1'b1;
  assign CLBLM_L_X56Y97_SLICE_X85Y97_C1 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign CLBLM_L_X56Y97_SLICE_X85Y97_C2 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLM_L_X56Y97_SLICE_X85Y97_C3 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLM_L_X56Y97_SLICE_X85Y97_C4 = CLBLM_R_X49Y107_SLICE_X75Y107_DQ;
  assign CLBLM_L_X56Y97_SLICE_X85Y97_C5 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLM_L_X56Y97_SLICE_X85Y97_C6 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLM_L_X56Y97_SLICE_X85Y97_CE = CLBLM_L_X60Y98_SLICE_X91Y98_DQ;
  assign CLBLM_L_X62Y109_SLICE_X92Y109_A1 = CLBLM_L_X60Y107_SLICE_X91Y107_B_XOR;
  assign CLBLM_L_X62Y109_SLICE_X92Y109_A2 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X62Y109_SLICE_X92Y109_A3 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_L_X62Y109_SLICE_X92Y109_A4 = CLBLM_R_X59Y103_SLICE_X89Y103_CQ;
  assign CLBLM_L_X62Y109_SLICE_X92Y109_A5 = CLBLM_L_X62Y107_SLICE_X92Y107_AQ;
  assign CLBLM_L_X62Y109_SLICE_X92Y109_A6 = CLBLM_L_X60Y110_SLICE_X91Y110_CO6;
  assign CLBLM_L_X56Y97_SLICE_X85Y97_D1 = CLBLM_L_X50Y105_SLICE_X76Y105_AQ;
  assign CLBLM_L_X56Y97_SLICE_X85Y97_D2 = CLBLM_L_X56Y97_SLICE_X85Y97_CQ;
  assign CLBLM_L_X56Y97_SLICE_X85Y97_D3 = CLBLM_L_X60Y98_SLICE_X90Y98_AQ;
  assign CLBLM_L_X56Y97_SLICE_X85Y97_D4 = CLBLM_L_X60Y97_SLICE_X90Y97_BO6;
  assign CLBLL_R_X57Y98_SLICE_X86Y98_A1 = CLBLL_L_X54Y99_SLICE_X83Y99_A5Q;
  assign CLBLL_R_X57Y98_SLICE_X86Y98_A2 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLL_R_X57Y98_SLICE_X86Y98_A3 = CLBLM_R_X53Y99_SLICE_X81Y99_AQ;
  assign CLBLL_R_X57Y98_SLICE_X86Y98_A4 = CLBLM_L_X62Y99_SLICE_X92Y99_AO6;
  assign CLBLL_R_X57Y98_SLICE_X86Y98_A5 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLL_R_X57Y98_SLICE_X86Y98_A6 = CLBLM_L_X56Y99_SLICE_X85Y99_A5Q;
  assign CLBLM_L_X56Y97_SLICE_X85Y97_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X56Y97_SLICE_X85Y97_D5 = CLBLM_L_X56Y97_SLICE_X84Y97_DQ;
  assign CLBLL_R_X57Y98_SLICE_X86Y98_B1 = CLBLL_L_X54Y99_SLICE_X83Y99_A5Q;
  assign CLBLL_R_X57Y98_SLICE_X86Y98_B2 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLL_R_X57Y98_SLICE_X86Y98_B3 = CLBLM_R_X53Y99_SLICE_X81Y99_AQ;
  assign CLBLL_R_X57Y98_SLICE_X86Y98_B4 = CLBLM_L_X62Y99_SLICE_X92Y99_AO6;
  assign CLBLL_R_X57Y98_SLICE_X86Y98_B5 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLL_R_X57Y98_SLICE_X86Y98_B6 = CLBLM_L_X56Y99_SLICE_X85Y99_A5Q;
  assign CLBLM_L_X56Y97_SLICE_X84Y97_A5 = CLBLM_R_X49Y107_SLICE_X75Y107_DQ;
  assign CLBLM_L_X56Y97_SLICE_X84Y97_A6 = 1'b1;
  assign CLBLL_R_X57Y98_SLICE_X86Y98_C1 = CLBLM_R_X53Y99_SLICE_X81Y99_AQ;
  assign CLBLL_R_X57Y98_SLICE_X86Y98_C2 = CLBLM_L_X56Y99_SLICE_X85Y99_A5Q;
  assign CLBLL_R_X57Y98_SLICE_X86Y98_C3 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLL_R_X57Y98_SLICE_X86Y98_C4 = CLBLL_L_X54Y99_SLICE_X83Y99_A5Q;
  assign CLBLL_R_X57Y98_SLICE_X86Y98_C5 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLL_R_X57Y98_SLICE_X86Y98_C6 = CLBLM_L_X62Y99_SLICE_X92Y99_AO6;
  assign CLBLM_L_X56Y97_SLICE_X84Y97_B1 = CLBLM_R_X49Y108_SLICE_X75Y108_DQ;
  assign CLBLM_L_X56Y97_SLICE_X84Y97_B2 = CLBLM_L_X56Y97_SLICE_X85Y97_BO5;
  assign CLBLM_L_X56Y97_SLICE_X84Y97_B3 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLM_L_X56Y97_SLICE_X84Y97_B4 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLM_L_X56Y97_SLICE_X84Y97_C1 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign CLBLM_L_X56Y97_SLICE_X84Y97_B5 = CLBLM_L_X56Y98_SLICE_X84Y98_CO6;
  assign CLBLM_L_X56Y97_SLICE_X84Y97_C4 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLL_R_X57Y98_SLICE_X86Y98_D1 = CLBLM_R_X53Y99_SLICE_X81Y99_AQ;
  assign CLBLL_R_X57Y98_SLICE_X86Y98_D2 = CLBLM_L_X56Y99_SLICE_X85Y99_A5Q;
  assign CLBLL_R_X57Y98_SLICE_X86Y98_D3 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLL_R_X57Y98_SLICE_X86Y98_D4 = CLBLL_L_X54Y99_SLICE_X83Y99_A5Q;
  assign CLBLL_R_X57Y98_SLICE_X86Y98_D5 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X56Y97_SLICE_X84Y97_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLL_R_X57Y98_SLICE_X86Y98_D6 = CLBLM_L_X62Y99_SLICE_X92Y99_AO6;
  assign CLBLM_L_X56Y97_SLICE_X84Y97_C3 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLM_L_X56Y97_SLICE_X84Y97_C5 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLM_L_X56Y97_SLICE_X84Y97_CE = CLBLM_L_X60Y98_SLICE_X91Y98_DQ;
  assign CLBLM_L_X56Y97_SLICE_X84Y97_D1 = CLBLM_L_X56Y98_SLICE_X84Y98_CO6;
  assign CLBLM_L_X56Y97_SLICE_X84Y97_D2 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLM_L_X56Y97_SLICE_X84Y97_D3 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLM_L_X56Y97_SLICE_X84Y97_D4 = CLBLM_L_X56Y97_SLICE_X84Y97_AO5;
  assign CLBLM_L_X56Y97_SLICE_X84Y97_D5 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLM_L_X56Y97_SLICE_X84Y97_D6 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign CLBLM_L_X56Y97_SLICE_X84Y97_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLL_R_X57Y98_SLICE_X87Y98_A1 = 1'b1;
  assign CLBLL_R_X57Y98_SLICE_X87Y98_A2 = 1'b1;
  assign CLBLL_R_X57Y98_SLICE_X87Y98_A3 = 1'b1;
  assign CLBLL_R_X57Y98_SLICE_X87Y98_A4 = 1'b1;
  assign CLBLL_R_X57Y98_SLICE_X87Y98_A5 = 1'b1;
  assign CLBLL_R_X57Y98_SLICE_X87Y98_A6 = 1'b1;
  assign CLBLL_R_X57Y98_SLICE_X87Y98_AX = CLBLM_R_X59Y98_SLICE_X89Y98_AQ;
  assign CLBLL_R_X57Y98_SLICE_X87Y98_B1 = 1'b1;
  assign CLBLL_R_X57Y98_SLICE_X87Y98_B2 = 1'b1;
  assign CLBLL_R_X57Y98_SLICE_X87Y98_B3 = 1'b1;
  assign CLBLL_R_X57Y98_SLICE_X87Y98_B4 = 1'b1;
  assign CLBLL_R_X57Y98_SLICE_X87Y98_B5 = 1'b1;
  assign CLBLL_R_X57Y98_SLICE_X87Y98_B6 = 1'b1;
  assign CLBLL_R_X57Y98_SLICE_X87Y98_BX = CLBLM_R_X59Y98_SLICE_X89Y98_A5Q;
  assign CLBLL_R_X57Y98_SLICE_X87Y98_C1 = 1'b1;
  assign CLBLL_R_X57Y98_SLICE_X87Y98_C2 = 1'b1;
  assign CLBLL_R_X57Y98_SLICE_X87Y98_C3 = 1'b1;
  assign CLBLL_R_X57Y98_SLICE_X87Y98_C4 = 1'b1;
  assign CLBLL_R_X57Y98_SLICE_X87Y98_C5 = 1'b1;
  assign CLBLL_R_X57Y98_SLICE_X87Y98_C6 = 1'b1;
  assign CLBLL_R_X57Y98_SLICE_X87Y98_CE = CLBLL_R_X57Y97_SLICE_X87Y97_AO6;
  assign CLBLL_R_X57Y98_SLICE_X87Y98_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLL_R_X57Y98_SLICE_X87Y98_CX = CLBLM_R_X59Y98_SLICE_X89Y98_CQ;
  assign CLBLL_R_X57Y98_SLICE_X87Y98_D1 = 1'b1;
  assign CLBLL_R_X57Y98_SLICE_X87Y98_D2 = 1'b1;
  assign CLBLL_R_X57Y98_SLICE_X87Y98_D3 = 1'b1;
  assign CLBLL_R_X57Y98_SLICE_X87Y98_D4 = 1'b1;
  assign CLBLL_R_X57Y98_SLICE_X87Y98_D5 = 1'b1;
  assign CLBLL_R_X57Y98_SLICE_X87Y98_D6 = 1'b1;
  assign CLBLL_R_X57Y98_SLICE_X87Y98_DX = CLBLM_R_X59Y98_SLICE_X89Y98_C5Q;
  assign CLBLL_R_X57Y98_SLICE_X87Y98_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLK_HROW_BOT_R_X139Y78_BUFHCE_X0Y20_CE = 1'b1;
  assign CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_CE = 1'b1;
  assign CLBLM_L_X62Y110_SLICE_X93Y110_A1 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_L_X62Y110_SLICE_X93Y110_A2 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y110_SLICE_X93Y110_A3 = CLBLM_L_X62Y110_SLICE_X93Y110_AQ;
  assign CLBLM_L_X62Y110_SLICE_X93Y110_A4 = CLBLM_L_X62Y105_SLICE_X92Y105_BO6;
  assign CLBLM_L_X62Y110_SLICE_X93Y110_A5 = CLBLM_L_X62Y110_SLICE_X93Y110_CO6;
  assign CLBLM_L_X62Y110_SLICE_X93Y110_A6 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X62Y110_SLICE_X93Y110_B1 = CLBLL_R_X57Y99_SLICE_X87Y99_AQ;
  assign CLBLM_L_X62Y110_SLICE_X93Y110_B2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_L_X62Y110_SLICE_X93Y110_B3 = CLBLM_L_X62Y110_SLICE_X93Y110_AQ;
  assign CLBLM_L_X62Y110_SLICE_X93Y110_B4 = CLBLM_R_X49Y119_SLICE_X74Y119_BQ;
  assign CLBLM_L_X62Y110_SLICE_X93Y110_B5 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLM_L_X62Y110_SLICE_X93Y110_B6 = CLBLM_R_X49Y119_SLICE_X74Y119_AQ;
  assign CLBLM_L_X62Y110_SLICE_X93Y110_C1 = CLBLM_R_X49Y119_SLICE_X74Y119_BQ;
  assign CLBLM_L_X62Y110_SLICE_X93Y110_C2 = 1'b1;
  assign CLBLM_L_X62Y110_SLICE_X93Y110_C3 = 1'b1;
  assign CLBLM_L_X62Y110_SLICE_X93Y110_C4 = 1'b1;
  assign CLBLM_L_X62Y110_SLICE_X93Y110_C5 = 1'b1;
  assign CLBLM_L_X62Y110_SLICE_X93Y110_C6 = CLBLM_R_X49Y119_SLICE_X74Y119_AQ;
  assign CLBLM_L_X56Y98_SLICE_X85Y98_A1 = CLBLM_R_X49Y104_SLICE_X75Y104_AQ;
  assign CLBLM_L_X56Y98_SLICE_X85Y98_A2 = CLBLM_L_X56Y100_SLICE_X85Y100_BO6;
  assign CLBLM_L_X62Y110_SLICE_X93Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X56Y98_SLICE_X85Y98_A3 = CLBLM_L_X56Y98_SLICE_X84Y98_CO6;
  assign CLBLM_L_X56Y98_SLICE_X85Y98_A4 = CLBLM_R_X49Y104_SLICE_X74Y104_AQ;
  assign CLBLM_L_X56Y98_SLICE_X85Y98_A5 = CLBLL_R_X57Y102_SLICE_X86Y102_CO6;
  assign CLBLM_L_X56Y98_SLICE_X85Y98_A6 = 1'b1;
  assign CLBLM_L_X62Y110_SLICE_X93Y110_D1 = 1'b1;
  assign CLBLM_L_X62Y110_SLICE_X93Y110_D2 = 1'b1;
  assign CLBLM_L_X62Y110_SLICE_X93Y110_D3 = 1'b1;
  assign CLBLM_L_X62Y110_SLICE_X93Y110_D4 = 1'b1;
  assign CLBLM_L_X62Y110_SLICE_X93Y110_D5 = 1'b1;
  assign CLBLM_L_X62Y110_SLICE_X93Y110_D6 = 1'b1;
  assign CLBLM_L_X56Y98_SLICE_X85Y98_B1 = CLBLL_L_X54Y98_SLICE_X83Y98_DO6;
  assign CLBLM_L_X56Y98_SLICE_X85Y98_B2 = CLBLL_L_X54Y102_SLICE_X82Y102_BO6;
  assign CLBLM_L_X62Y110_SLICE_X93Y110_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X56Y98_SLICE_X85Y98_B3 = CLBLL_R_X57Y103_SLICE_X86Y103_AQ;
  assign CLBLM_L_X56Y98_SLICE_X85Y98_B4 = CLBLM_R_X49Y104_SLICE_X74Y104_AQ;
  assign CLBLM_L_X56Y98_SLICE_X85Y98_B5 = CLBLL_R_X57Y103_SLICE_X86Y103_A5Q;
  assign CLBLM_L_X62Y110_SLICE_X92Y110_A1 = CLBLM_R_X59Y112_SLICE_X89Y112_CO6;
  assign CLBLM_L_X62Y110_SLICE_X92Y110_A2 = CLBLM_R_X49Y106_SLICE_X75Y106_DQ;
  assign CLBLM_L_X62Y110_SLICE_X92Y110_A3 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y110_SLICE_X92Y110_A4 = CLBLM_R_X59Y103_SLICE_X89Y103_DQ;
  assign CLBLM_L_X62Y110_SLICE_X92Y110_A5 = 1'b1;
  assign CLBLM_L_X62Y110_SLICE_X92Y110_A6 = CLBLM_L_X62Y110_SLICE_X92Y110_CO6;
  assign CLBLM_L_X56Y98_SLICE_X85Y98_C2 = CLBLL_R_X57Y103_SLICE_X86Y103_A5Q;
  assign CLBLM_L_X56Y98_SLICE_X85Y98_C3 = CLBLL_L_X54Y98_SLICE_X83Y98_DO6;
  assign CLBLM_L_X56Y98_SLICE_X85Y98_C4 = CLBLM_R_X49Y108_SLICE_X75Y108_DQ;
  assign CLBLM_L_X56Y98_SLICE_X85Y98_C6 = 1'b1;
  assign CLBLM_L_X62Y110_SLICE_X92Y110_B1 = CLBLM_L_X62Y109_SLICE_X92Y109_AO6;
  assign CLBLM_L_X62Y110_SLICE_X92Y110_B2 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLM_L_X62Y110_SLICE_X92Y110_B3 = 1'b1;
  assign CLBLM_L_X62Y110_SLICE_X92Y110_B4 = CLBLM_R_X59Y103_SLICE_X89Y103_DQ;
  assign CLBLM_L_X62Y110_SLICE_X92Y110_B5 = CLBLM_R_X59Y110_SLICE_X89Y110_BO6;
  assign CLBLM_L_X62Y110_SLICE_X92Y110_B6 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLL_R_X57Y99_SLICE_X86Y99_A1 = CLBLL_R_X57Y101_SLICE_X87Y101_BO5;
  assign CLBLL_R_X57Y99_SLICE_X86Y99_A2 = CLBLM_L_X56Y98_SLICE_X84Y98_BQ;
  assign CLBLL_R_X57Y99_SLICE_X86Y99_A3 = CLBLM_R_X59Y96_SLICE_X89Y96_A5Q;
  assign CLBLM_L_X62Y110_SLICE_X92Y110_C1 = CLBLM_L_X60Y106_SLICE_X91Y106_B_XOR;
  assign CLBLM_L_X62Y110_SLICE_X92Y110_C2 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLM_L_X62Y110_SLICE_X92Y110_C3 = CLBLM_L_X62Y106_SLICE_X92Y106_BQ;
  assign CLBLM_L_X62Y110_SLICE_X92Y110_C4 = CLBLM_R_X59Y103_SLICE_X89Y103_CQ;
  assign CLBLM_L_X62Y110_SLICE_X92Y110_C5 = CLBLM_L_X60Y110_SLICE_X91Y110_DO6;
  assign CLBLM_L_X62Y110_SLICE_X92Y110_C6 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_L_X62Y110_SLICE_X92Y110_CE = CLBLM_R_X59Y99_SLICE_X89Y99_CO6;
  assign CLBLL_R_X57Y99_SLICE_X86Y99_B1 = CLBLL_R_X57Y101_SLICE_X87Y101_BO5;
  assign CLBLL_R_X57Y99_SLICE_X86Y99_B2 = CLBLM_L_X56Y98_SLICE_X84Y98_BQ;
  assign CLBLM_L_X62Y110_SLICE_X92Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X57Y99_SLICE_X86Y99_B4 = CLBLL_L_X54Y99_SLICE_X82Y99_CQ;
  assign CLBLL_R_X57Y99_SLICE_X86Y99_B5 = CLBLM_R_X59Y96_SLICE_X89Y96_A5Q;
  assign CLBLL_R_X57Y99_SLICE_X86Y99_B6 = CLBLM_L_X62Y101_SLICE_X93Y101_CQ;
  assign CLBLL_R_X57Y99_SLICE_X86Y99_C1 = 1'b1;
  assign CLBLM_L_X62Y110_SLICE_X92Y110_D1 = CLBLM_L_X62Y108_SLICE_X92Y108_AQ;
  assign CLBLM_L_X62Y110_SLICE_X92Y110_D2 = 1'b1;
  assign CLBLM_L_X62Y110_SLICE_X92Y110_D3 = CLBLM_L_X62Y110_SLICE_X92Y110_BQ;
  assign CLBLM_L_X62Y110_SLICE_X92Y110_D4 = CLBLM_L_X62Y111_SLICE_X92Y111_CO6;
  assign CLBLM_L_X62Y110_SLICE_X92Y110_D5 = CLBLM_L_X62Y108_SLICE_X93Y108_AQ;
  assign CLBLM_L_X62Y110_SLICE_X92Y110_D6 = CLBLM_L_X60Y111_SLICE_X91Y111_AQ;
  assign CLBLL_R_X57Y99_SLICE_X86Y99_C6 = 1'b1;
  assign CLBLL_R_X57Y99_SLICE_X86Y99_CE = CLBLL_R_X57Y100_SLICE_X87Y100_DO6;
  assign CLBLL_R_X57Y99_SLICE_X86Y99_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X62Y110_SLICE_X92Y110_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X56Y98_SLICE_X84Y98_BX = CLBLM_L_X56Y98_SLICE_X84Y98_AO5;
  assign CLBLL_R_X57Y99_SLICE_X86Y99_D1 = 1'b1;
  assign CLBLL_R_X57Y99_SLICE_X86Y99_D2 = 1'b1;
  assign CLBLL_R_X57Y99_SLICE_X86Y99_D3 = 1'b1;
  assign CLBLL_R_X57Y99_SLICE_X86Y99_D4 = 1'b1;
  assign CLBLL_R_X57Y99_SLICE_X86Y99_D5 = 1'b1;
  assign CLBLL_R_X57Y99_SLICE_X86Y99_D6 = 1'b1;
  assign CLBLL_R_X57Y99_SLICE_X86Y99_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X56Y98_SLICE_X84Y98_C5 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLM_L_X56Y98_SLICE_X84Y98_C6 = CLBLL_L_X54Y102_SLICE_X82Y102_BO6;
  assign CLBLM_L_X56Y98_SLICE_X84Y98_CE = CLBLM_L_X56Y98_SLICE_X84Y98_DO6;
  assign CLBLM_L_X56Y98_SLICE_X84Y98_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_L_X56Y98_SLICE_X84Y98_D1 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLM_L_X56Y98_SLICE_X84Y98_D2 = CLBLM_L_X60Y98_SLICE_X91Y98_CQ;
  assign CLBLM_L_X56Y98_SLICE_X84Y98_D3 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLM_L_X56Y98_SLICE_X84Y98_D4 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_L_X56Y98_SLICE_X84Y98_D5 = 1'b1;
  assign CLBLM_L_X56Y98_SLICE_X84Y98_D6 = 1'b1;
  assign CLBLM_L_X56Y105_SLICE_X85Y105_C1 = CLBLM_L_X62Y100_SLICE_X92Y100_AO5;
  assign CLBLM_L_X56Y98_SLICE_X84Y98_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X56Y105_SLICE_X85Y105_C2 = CLBLM_L_X56Y105_SLICE_X85Y105_CQ;
  assign CLBLL_R_X57Y99_SLICE_X87Y99_A1 = CLBLL_R_X57Y99_SLICE_X87Y99_AQ;
  assign CLBLL_R_X57Y99_SLICE_X87Y99_A2 = CLBLL_R_X57Y100_SLICE_X86Y100_AO6;
  assign CLBLL_R_X57Y99_SLICE_X87Y99_A3 = CLBLM_R_X59Y100_SLICE_X88Y100_AO6;
  assign CLBLL_R_X57Y99_SLICE_X87Y99_A4 = CLBLM_L_X62Y99_SLICE_X92Y99_AO6;
  assign CLBLL_R_X57Y99_SLICE_X87Y99_A5 = CLBLM_L_X60Y98_SLICE_X90Y98_CO5;
  assign CLBLL_R_X57Y99_SLICE_X87Y99_A6 = CLBLL_R_X57Y99_SLICE_X87Y99_CO6;
  assign CLBLM_L_X56Y105_SLICE_X85Y105_C5 = CLBLM_L_X50Y107_SLICE_X76Y107_BQ;
  assign CLBLL_R_X57Y99_SLICE_X87Y99_B1 = CLBLM_L_X56Y99_SLICE_X84Y99_BQ;
  assign CLBLL_R_X57Y99_SLICE_X87Y99_B2 = CLBLM_L_X56Y99_SLICE_X84Y99_AQ;
  assign CLBLL_R_X57Y99_SLICE_X87Y99_B3 = CLBLM_L_X60Y98_SLICE_X91Y98_CQ;
  assign CLBLL_R_X57Y99_SLICE_X87Y99_B4 = 1'b1;
  assign CLBLL_R_X57Y99_SLICE_X87Y99_B5 = 1'b1;
  assign CLBLL_R_X57Y99_SLICE_X87Y99_B6 = 1'b1;
  assign CLBLL_R_X57Y99_SLICE_X87Y99_C1 = 1'b1;
  assign CLBLL_R_X57Y99_SLICE_X87Y99_C2 = CLBLM_L_X56Y99_SLICE_X85Y99_BQ;
  assign CLBLL_R_X57Y99_SLICE_X87Y99_C3 = CLBLL_L_X54Y99_SLICE_X82Y99_CQ;
  assign CLBLL_R_X57Y99_SLICE_X87Y99_C4 = 1'b1;
  assign CLBLL_R_X57Y99_SLICE_X87Y99_C5 = 1'b1;
  assign CLBLL_R_X57Y99_SLICE_X87Y99_C6 = 1'b1;
  assign CLBLL_R_X57Y99_SLICE_X87Y99_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLL_R_X57Y99_SLICE_X87Y99_D1 = 1'b1;
  assign CLBLL_R_X57Y99_SLICE_X87Y99_D2 = 1'b1;
  assign CLBLL_R_X57Y99_SLICE_X87Y99_D3 = 1'b1;
  assign CLBLL_R_X57Y99_SLICE_X87Y99_D4 = 1'b1;
  assign CLBLL_R_X57Y99_SLICE_X87Y99_D5 = 1'b1;
  assign CLBLL_R_X57Y99_SLICE_X87Y99_D6 = 1'b1;
  assign CLBLL_R_X57Y99_SLICE_X87Y99_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_D = LIOB33_X0Y119_IOB_X0Y120_I;
  assign LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y119_D = LIOB33_X0Y119_IOB_X0Y119_I;
  assign CLBLM_L_X56Y105_SLICE_X84Y105_B1 = CLBLL_L_X54Y107_SLICE_X82Y107_C_XOR;
  assign CLBLM_L_X56Y105_SLICE_X84Y105_B2 = CLBLM_L_X56Y105_SLICE_X84Y105_BQ;
  assign CLBLM_L_X62Y111_SLICE_X93Y111_A1 = 1'b1;
  assign CLBLM_L_X62Y111_SLICE_X93Y111_A2 = 1'b1;
  assign CLBLM_L_X62Y111_SLICE_X93Y111_A3 = 1'b1;
  assign CLBLM_L_X62Y111_SLICE_X93Y111_A4 = 1'b1;
  assign CLBLM_L_X62Y111_SLICE_X93Y111_A5 = 1'b1;
  assign CLBLM_L_X62Y111_SLICE_X93Y111_A6 = 1'b1;
  assign CLBLM_L_X62Y111_SLICE_X93Y111_B1 = 1'b1;
  assign CLBLM_L_X62Y111_SLICE_X93Y111_B2 = 1'b1;
  assign CLBLM_L_X62Y111_SLICE_X93Y111_B3 = 1'b1;
  assign CLBLM_L_X62Y111_SLICE_X93Y111_B4 = 1'b1;
  assign CLBLM_L_X62Y111_SLICE_X93Y111_B5 = 1'b1;
  assign CLBLM_L_X62Y111_SLICE_X93Y111_B6 = 1'b1;
  assign CLBLM_L_X56Y105_SLICE_X84Y105_B5 = CLBLL_L_X54Y101_SLICE_X83Y101_BO6;
  assign CLBLM_L_X62Y111_SLICE_X93Y111_C1 = 1'b1;
  assign CLBLM_L_X62Y111_SLICE_X93Y111_C2 = 1'b1;
  assign CLBLM_L_X62Y111_SLICE_X93Y111_C3 = 1'b1;
  assign CLBLM_L_X62Y111_SLICE_X93Y111_C4 = 1'b1;
  assign CLBLM_L_X62Y111_SLICE_X93Y111_C5 = 1'b1;
  assign CLBLM_L_X62Y111_SLICE_X93Y111_C6 = 1'b1;
  assign CLBLM_L_X56Y99_SLICE_X85Y99_A1 = 1'b1;
  assign CLBLM_L_X56Y99_SLICE_X85Y99_A2 = 1'b1;
  assign CLBLM_L_X56Y99_SLICE_X85Y99_A3 = 1'b1;
  assign CLBLM_L_X56Y99_SLICE_X85Y99_A4 = CLBLL_R_X57Y102_SLICE_X86Y102_AO6;
  assign CLBLM_L_X56Y99_SLICE_X85Y99_A5 = 1'b1;
  assign CLBLM_L_X56Y99_SLICE_X85Y99_A6 = CLBLL_L_X52Y99_SLICE_X79Y99_AO6;
  assign CLBLM_L_X56Y99_SLICE_X85Y99_AX = CLBLM_L_X56Y99_SLICE_X85Y99_AQ;
  assign CLBLM_L_X56Y99_SLICE_X85Y99_B1 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLM_L_X62Y111_SLICE_X93Y111_D1 = 1'b1;
  assign CLBLM_L_X62Y111_SLICE_X93Y111_D2 = 1'b1;
  assign CLBLM_L_X62Y111_SLICE_X93Y111_D3 = 1'b1;
  assign CLBLM_L_X62Y111_SLICE_X93Y111_D4 = 1'b1;
  assign CLBLM_L_X62Y111_SLICE_X93Y111_D5 = 1'b1;
  assign CLBLM_L_X62Y111_SLICE_X93Y111_D6 = 1'b1;
  assign CLBLM_L_X56Y99_SLICE_X85Y99_B2 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLM_L_X56Y99_SLICE_X85Y99_B3 = CLBLM_L_X56Y97_SLICE_X84Y97_CO5;
  assign CLBLM_L_X56Y99_SLICE_X85Y99_B4 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign CLBLM_L_X56Y99_SLICE_X85Y99_B5 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLM_L_X56Y99_SLICE_X85Y99_B6 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLM_L_X62Y111_SLICE_X92Y111_A1 = CLBLM_L_X60Y112_SLICE_X90Y112_BO6;
  assign CLBLM_L_X62Y111_SLICE_X92Y111_A2 = CLBLM_L_X62Y108_SLICE_X92Y108_CO6;
  assign CLBLM_L_X62Y111_SLICE_X92Y111_A3 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y111_SLICE_X92Y111_A4 = CLBLM_L_X60Y112_SLICE_X90Y112_AO6;
  assign CLBLM_L_X62Y111_SLICE_X92Y111_A5 = CLBLM_L_X62Y108_SLICE_X93Y108_BO6;
  assign CLBLM_L_X62Y111_SLICE_X92Y111_A6 = 1'b1;
  assign CLBLM_L_X56Y99_SLICE_X85Y99_C2 = CLBLL_L_X54Y102_SLICE_X82Y102_AO5;
  assign CLBLM_L_X56Y99_SLICE_X85Y99_C3 = CLBLM_R_X49Y104_SLICE_X75Y104_DQ;
  assign CLBLM_L_X56Y99_SLICE_X85Y99_C4 = 1'b1;
  assign CLBLM_L_X56Y99_SLICE_X85Y99_C6 = CLBLM_L_X56Y102_SLICE_X85Y102_BO6;
  assign CLBLM_L_X62Y111_SLICE_X92Y111_B1 = CLBLM_L_X62Y111_SLICE_X92Y111_DO6;
  assign CLBLM_L_X62Y111_SLICE_X92Y111_B2 = CLBLM_L_X60Y111_SLICE_X91Y111_AQ;
  assign CLBLM_L_X62Y111_SLICE_X92Y111_B3 = CLBLM_L_X62Y111_SLICE_X92Y111_AQ;
  assign CLBLM_L_X62Y111_SLICE_X92Y111_B4 = CLBLM_L_X62Y108_SLICE_X92Y108_A5Q;
  assign CLBLM_L_X62Y111_SLICE_X92Y111_B5 = CLBLM_L_X62Y108_SLICE_X92Y108_AQ;
  assign CLBLM_L_X62Y111_SLICE_X92Y111_B6 = CLBLM_L_X62Y111_SLICE_X92Y111_A5Q;
  assign CLBLL_R_X57Y100_SLICE_X86Y100_A4 = CLBLM_L_X56Y98_SLICE_X84Y98_AQ;
  assign CLBLL_R_X57Y100_SLICE_X86Y100_A5 = CLBLL_L_X54Y98_SLICE_X83Y98_BQ;
  assign CLBLL_R_X57Y100_SLICE_X86Y100_A6 = 1'b1;
  assign CLBLM_L_X62Y111_SLICE_X92Y111_C1 = CLBLM_L_X60Y111_SLICE_X91Y111_BQ;
  assign CLBLM_L_X62Y111_SLICE_X92Y111_C2 = CLBLM_L_X62Y111_SLICE_X92Y111_AQ;
  assign CLBLM_L_X62Y111_SLICE_X92Y111_C3 = CLBLM_L_X60Y111_SLICE_X90Y111_AQ;
  assign CLBLM_L_X62Y111_SLICE_X92Y111_C4 = CLBLM_L_X62Y111_SLICE_X92Y111_A5Q;
  assign CLBLM_L_X62Y111_SLICE_X92Y111_C5 = CLBLM_L_X62Y110_SLICE_X92Y110_AQ;
  assign CLBLM_L_X62Y111_SLICE_X92Y111_C6 = CLBLM_L_X62Y108_SLICE_X92Y108_A5Q;
  assign CLBLM_L_X62Y111_SLICE_X92Y111_CE = CLBLM_R_X59Y99_SLICE_X89Y99_CO6;
  assign CLBLL_R_X57Y100_SLICE_X86Y100_B6 = CLBLM_L_X56Y100_SLICE_X85Y100_AQ;
  assign CLBLM_L_X62Y111_SLICE_X92Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X56Y99_SLICE_X84Y99_A1 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLL_R_X57Y100_SLICE_X86Y100_C1 = CLBLM_L_X56Y99_SLICE_X85Y99_BQ;
  assign CLBLL_R_X57Y100_SLICE_X86Y100_C2 = CLBLM_L_X60Y100_SLICE_X90Y100_AO5;
  assign CLBLL_R_X57Y100_SLICE_X86Y100_C3 = CLBLM_L_X62Y100_SLICE_X92Y100_BQ;
  assign CLBLL_R_X57Y100_SLICE_X86Y100_C4 = CLBLM_R_X59Y98_SLICE_X89Y98_A5Q;
  assign CLBLM_L_X62Y111_SLICE_X92Y111_D1 = CLBLM_L_X62Y110_SLICE_X92Y110_BQ;
  assign CLBLM_L_X62Y111_SLICE_X92Y111_D2 = CLBLM_L_X60Y111_SLICE_X90Y111_AQ;
  assign CLBLM_L_X62Y111_SLICE_X92Y111_D3 = CLBLM_L_X62Y108_SLICE_X93Y108_AQ;
  assign CLBLM_L_X62Y111_SLICE_X92Y111_D4 = 1'b1;
  assign CLBLM_L_X62Y111_SLICE_X92Y111_D5 = CLBLM_L_X62Y110_SLICE_X92Y110_AQ;
  assign CLBLM_L_X62Y111_SLICE_X92Y111_D6 = CLBLM_L_X60Y111_SLICE_X91Y111_BQ;
  assign CLBLL_R_X57Y100_SLICE_X86Y100_D1 = CLBLM_L_X60Y100_SLICE_X90Y100_AO6;
  assign CLBLL_R_X57Y100_SLICE_X86Y100_D2 = CLBLM_R_X59Y98_SLICE_X89Y98_AQ;
  assign CLBLM_L_X62Y111_SLICE_X92Y111_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLL_R_X57Y100_SLICE_X86Y100_D3 = CLBLM_L_X56Y98_SLICE_X84Y98_AQ;
  assign CLBLL_R_X57Y100_SLICE_X86Y100_D4 = CLBLM_L_X62Y100_SLICE_X92Y100_AQ;
  assign CLBLL_R_X57Y100_SLICE_X86Y100_D5 = CLBLM_L_X56Y99_SLICE_X85Y99_BQ;
  assign CLBLL_R_X57Y100_SLICE_X86Y100_D6 = CLBLL_L_X54Y99_SLICE_X82Y99_CQ;
  assign CLBLL_R_X57Y100_SLICE_X86Y100_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X56Y99_SLICE_X84Y99_C1 = CLBLM_L_X56Y97_SLICE_X84Y97_CO5;
  assign CLBLM_L_X56Y99_SLICE_X84Y99_C2 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLM_L_X56Y99_SLICE_X84Y99_C3 = CLBLM_L_X56Y97_SLICE_X85Y97_BO5;
  assign CLBLM_L_X56Y99_SLICE_X84Y99_C4 = CLBLM_R_X49Y107_SLICE_X75Y107_DQ;
  assign CLBLM_L_X56Y99_SLICE_X84Y99_C5 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLM_L_X56Y99_SLICE_X84Y99_CE = CLBLM_L_X60Y98_SLICE_X91Y98_BQ;
  assign CLBLM_L_X56Y99_SLICE_X84Y99_D1 = 1'b1;
  assign CLBLM_L_X56Y99_SLICE_X84Y99_D2 = 1'b1;
  assign CLBLM_L_X56Y99_SLICE_X84Y99_D3 = 1'b1;
  assign CLBLM_L_X56Y99_SLICE_X84Y99_D4 = 1'b1;
  assign CLBLM_L_X56Y99_SLICE_X84Y99_D5 = 1'b1;
  assign CLBLM_L_X56Y99_SLICE_X84Y99_D6 = 1'b1;
  assign CLBLM_L_X56Y99_SLICE_X84Y99_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLL_R_X57Y100_SLICE_X87Y100_A1 = 1'b1;
  assign CLBLL_R_X57Y100_SLICE_X87Y100_A2 = CLBLM_R_X59Y98_SLICE_X89Y98_B5Q;
  assign CLBLL_R_X57Y100_SLICE_X87Y100_A3 = CLBLL_L_X54Y98_SLICE_X83Y98_BQ;
  assign CLBLL_R_X57Y100_SLICE_X87Y100_A4 = CLBLM_L_X60Y101_SLICE_X91Y101_CO5;
  assign CLBLL_R_X57Y100_SLICE_X87Y100_A5 = CLBLM_L_X56Y100_SLICE_X85Y100_BQ;
  assign CLBLL_R_X57Y100_SLICE_X87Y100_A6 = CLBLL_L_X54Y99_SLICE_X82Y99_AQ;
  assign CLBLM_L_X56Y105_SLICE_X84Y105_D1 = 1'b1;
  assign CLBLM_L_X56Y105_SLICE_X84Y105_D2 = 1'b1;
  assign CLBLL_R_X57Y100_SLICE_X87Y100_B1 = CLBLM_R_X59Y96_SLICE_X89Y96_AQ;
  assign CLBLL_R_X57Y100_SLICE_X87Y100_B2 = CLBLL_R_X57Y101_SLICE_X87Y101_BO6;
  assign CLBLL_R_X57Y100_SLICE_X87Y100_B3 = CLBLL_L_X54Y98_SLICE_X83Y98_BQ;
  assign CLBLL_R_X57Y100_SLICE_X87Y100_B4 = 1'b1;
  assign CLBLL_R_X57Y100_SLICE_X87Y100_B5 = CLBLM_L_X56Y100_SLICE_X85Y100_DQ;
  assign CLBLL_R_X57Y100_SLICE_X87Y100_B6 = CLBLL_L_X54Y99_SLICE_X82Y99_AQ;
  assign CLBLM_L_X56Y105_SLICE_X84Y105_D3 = 1'b1;
  assign CLBLM_L_X56Y105_SLICE_X84Y105_D4 = 1'b1;
  assign CLBLL_R_X57Y100_SLICE_X87Y100_C1 = CLBLM_R_X59Y98_SLICE_X89Y98_B5Q;
  assign CLBLL_R_X57Y100_SLICE_X87Y100_C2 = CLBLL_L_X54Y99_SLICE_X82Y99_CQ;
  assign CLBLL_R_X57Y100_SLICE_X87Y100_C3 = CLBLM_L_X60Y101_SLICE_X91Y101_CO5;
  assign CLBLL_R_X57Y100_SLICE_X87Y100_C4 = CLBLM_L_X62Y100_SLICE_X92Y100_CQ;
  assign CLBLL_R_X57Y100_SLICE_X87Y100_C5 = CLBLM_L_X56Y100_SLICE_X85Y100_BQ;
  assign CLBLL_R_X57Y100_SLICE_X87Y100_C6 = CLBLM_L_X56Y99_SLICE_X85Y99_BQ;
  assign CLBLL_R_X57Y100_SLICE_X87Y100_CE = CLBLL_R_X57Y100_SLICE_X87Y100_DO6;
  assign CLBLM_L_X56Y105_SLICE_X84Y105_D5 = 1'b1;
  assign CLBLL_R_X57Y100_SLICE_X87Y100_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X56Y105_SLICE_X84Y105_D6 = 1'b1;
  assign CLBLL_R_X57Y100_SLICE_X87Y100_D1 = 1'b1;
  assign CLBLL_R_X57Y100_SLICE_X87Y100_D2 = CLBLM_L_X60Y98_SLICE_X91Y98_BQ;
  assign CLBLL_R_X57Y100_SLICE_X87Y100_D3 = 1'b1;
  assign CLBLL_R_X57Y100_SLICE_X87Y100_D4 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLL_R_X57Y100_SLICE_X87Y100_D5 = 1'b1;
  assign CLBLL_R_X57Y100_SLICE_X87Y100_D6 = 1'b1;
  assign CLBLL_R_X57Y100_SLICE_X87Y100_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X56Y105_SLICE_X84Y105_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X62Y112_SLICE_X93Y112_A1 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X93Y112_A2 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X93Y112_A3 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X93Y112_A4 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X93Y112_A5 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X93Y112_A6 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X93Y112_B1 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X93Y112_B2 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X93Y112_B3 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X93Y112_B4 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X93Y112_B5 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X93Y112_B6 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X93Y112_C1 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X93Y112_C2 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X93Y112_C3 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X93Y112_C4 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X93Y112_C5 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X93Y112_C6 = 1'b1;
  assign CLBLM_L_X56Y100_SLICE_X85Y100_A1 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLM_L_X56Y100_SLICE_X85Y100_A2 = 1'b1;
  assign CLBLM_L_X56Y100_SLICE_X85Y100_A3 = 1'b1;
  assign CLBLM_L_X56Y100_SLICE_X85Y100_A4 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLM_L_X56Y100_SLICE_X85Y100_A5 = CLBLM_R_X49Y107_SLICE_X75Y107_DQ;
  assign CLBLM_L_X56Y100_SLICE_X85Y100_A6 = 1'b1;
  assign CLBLM_L_X56Y100_SLICE_X85Y100_AX = CLBLM_L_X56Y100_SLICE_X85Y100_BO5;
  assign CLBLM_L_X56Y100_SLICE_X85Y100_B1 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLM_L_X62Y112_SLICE_X93Y112_D1 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X93Y112_D2 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X93Y112_D3 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X93Y112_D4 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X93Y112_D5 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X93Y112_D6 = 1'b1;
  assign CLBLM_L_X56Y100_SLICE_X85Y100_B2 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLM_L_X56Y100_SLICE_X85Y100_B3 = CLBLM_R_X49Y108_SLICE_X75Y108_DQ;
  assign CLBLM_L_X56Y100_SLICE_X85Y100_B4 = CLBLM_L_X56Y97_SLICE_X84Y97_CO5;
  assign CLBLM_L_X56Y100_SLICE_X85Y100_B5 = CLBLM_R_X49Y107_SLICE_X75Y107_DQ;
  assign CLBLM_L_X56Y100_SLICE_X85Y100_B6 = 1'b1;
  assign CLBLM_L_X56Y100_SLICE_X85Y100_BX = CLBLM_L_X56Y100_SLICE_X85Y100_AO6;
  assign CLBLM_L_X56Y100_SLICE_X85Y100_C1 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X92Y112_A2 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X92Y112_A3 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X62Y112_SLICE_X92Y112_A4 = 1'b1;
  assign CLBLM_L_X56Y100_SLICE_X85Y100_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X62Y112_SLICE_X92Y112_A5 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X92Y112_A6 = 1'b1;
  assign CLBLM_L_X56Y100_SLICE_X85Y100_C3 = 1'b1;
  assign CLBLM_L_X56Y100_SLICE_X85Y100_C4 = 1'b1;
  assign CLBLM_L_X56Y100_SLICE_X85Y100_CX = CLBLM_L_X56Y100_SLICE_X85Y100_AO5;
  assign CLBLM_L_X56Y100_SLICE_X85Y100_D1 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X92Y112_B2 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X92Y112_B3 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X92Y112_B4 = 1'b1;
  assign CLBLM_L_X56Y100_SLICE_X85Y100_D5 = 1'b1;
  assign CLBLM_L_X56Y100_SLICE_X85Y100_D6 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X92Y112_B5 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X92Y112_B6 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X92Y112_B1 = 1'b1;
  assign CLBLL_R_X57Y101_SLICE_X86Y101_B3 = CLBLM_L_X60Y99_SLICE_X91Y99_AO5;
  assign CLBLM_L_X62Y112_SLICE_X92Y112_C1 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X92Y112_C2 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X92Y112_C3 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X92Y112_C4 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X92Y112_C5 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X92Y112_C6 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X92Y112_CE = CLBLM_L_X62Y110_SLICE_X93Y110_BO6;
  assign CLBLM_L_X56Y100_SLICE_X85Y100_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLL_R_X57Y101_SLICE_X86Y101_C2 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X92Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X57Y101_SLICE_X86Y101_C4 = 1'b1;
  assign CLBLL_R_X57Y101_SLICE_X86Y101_C5 = 1'b1;
  assign CLBLL_R_X57Y101_SLICE_X86Y101_C6 = 1'b1;
  assign CLBLL_R_X57Y101_SLICE_X86Y101_CE = CLBLM_L_X60Y100_SLICE_X90Y100_BO6;
  assign CLBLM_L_X56Y100_SLICE_X84Y100_B3 = CLBLM_L_X56Y102_SLICE_X85Y102_AQ;
  assign CLBLM_L_X62Y112_SLICE_X92Y112_D1 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X92Y112_D2 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X92Y112_D3 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X92Y112_D4 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X92Y112_D5 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X92Y112_D6 = 1'b1;
  assign CLBLL_R_X57Y101_SLICE_X86Y101_D1 = 1'b1;
  assign CLBLL_R_X57Y101_SLICE_X86Y101_D2 = 1'b1;
  assign CLBLL_R_X57Y101_SLICE_X86Y101_D3 = 1'b1;
  assign CLBLM_L_X62Y112_SLICE_X92Y112_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLL_R_X57Y101_SLICE_X86Y101_D6 = 1'b1;
  assign CLBLL_R_X57Y101_SLICE_X86Y101_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X56Y100_SLICE_X84Y100_BX = 1'b0;
  assign CLBLM_L_X56Y100_SLICE_X84Y100_C1 = CLBLM_L_X56Y102_SLICE_X85Y102_AQ;
  assign CLBLM_L_X56Y100_SLICE_X84Y100_C2 = CLBLM_L_X56Y100_SLICE_X84Y100_CQ;
  assign CLBLM_L_X56Y100_SLICE_X84Y100_C3 = CLBLM_L_X56Y102_SLICE_X85Y102_A5Q;
  assign CLBLM_L_X56Y100_SLICE_X84Y100_C4 = 1'b1;
  assign CLBLM_L_X56Y100_SLICE_X84Y100_C5 = 1'b1;
  assign CLBLM_L_X56Y100_SLICE_X84Y100_C6 = 1'b1;
  assign CLBLM_L_X56Y100_SLICE_X84Y100_CE = CLBLM_L_X56Y102_SLICE_X85Y102_CO6;
  assign CLBLM_L_X56Y100_SLICE_X84Y100_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X56Y100_SLICE_X84Y100_CX = 1'b0;
  assign CLBLM_L_X56Y100_SLICE_X84Y100_D1 = CLBLM_L_X56Y102_SLICE_X85Y102_AQ;
  assign CLBLM_L_X56Y100_SLICE_X84Y100_D2 = 1'b1;
  assign CLBLM_L_X56Y100_SLICE_X84Y100_D3 = CLBLM_L_X56Y100_SLICE_X84Y100_DQ;
  assign CLBLM_L_X56Y100_SLICE_X84Y100_D4 = 1'b1;
  assign CLBLM_L_X56Y100_SLICE_X84Y100_D5 = CLBLM_L_X56Y102_SLICE_X85Y102_A5Q;
  assign CLBLM_L_X56Y100_SLICE_X84Y100_D6 = 1'b1;
  assign CLBLL_R_X57Y101_SLICE_X87Y101_A1 = 1'b1;
  assign CLBLL_R_X57Y101_SLICE_X87Y101_A2 = CLBLM_L_X62Y101_SLICE_X92Y101_DO6;
  assign CLBLL_R_X57Y101_SLICE_X87Y101_A3 = CLBLL_L_X54Y98_SLICE_X83Y98_BQ;
  assign CLBLL_R_X57Y101_SLICE_X87Y101_A4 = CLBLL_L_X54Y99_SLICE_X82Y99_AQ;
  assign CLBLL_R_X57Y101_SLICE_X87Y101_A5 = CLBLL_L_X54Y101_SLICE_X82Y101_BQ;
  assign CLBLL_R_X57Y101_SLICE_X87Y101_A6 = CLBLM_R_X59Y98_SLICE_X89Y98_CQ;
  assign CLBLM_L_X56Y100_SLICE_X84Y100_DX = 1'b0;
  assign CLBLM_L_X56Y100_SLICE_X84Y100_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLL_R_X57Y101_SLICE_X87Y101_B1 = CLBLM_L_X62Y101_SLICE_X92Y101_CQ;
  assign CLBLL_R_X57Y101_SLICE_X87Y101_B2 = CLBLM_L_X62Y99_SLICE_X92Y99_BQ;
  assign CLBLL_R_X57Y101_SLICE_X87Y101_B3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_R_X57Y101_SLICE_X87Y101_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_R_X57Y101_SLICE_X87Y101_B5 = CLBLM_L_X60Y101_SLICE_X91Y101_BQ;
  assign CLBLL_R_X57Y101_SLICE_X87Y101_B6 = 1'b1;
  assign CLBLL_R_X57Y101_SLICE_X87Y101_C1 = CLBLL_L_X54Y101_SLICE_X82Y101_BQ;
  assign CLBLL_R_X57Y101_SLICE_X87Y101_C2 = CLBLM_R_X59Y98_SLICE_X89Y98_CQ;
  assign CLBLL_R_X57Y101_SLICE_X87Y101_C3 = CLBLL_L_X54Y99_SLICE_X82Y99_CQ;
  assign CLBLL_R_X57Y101_SLICE_X87Y101_C4 = CLBLM_L_X56Y99_SLICE_X85Y99_BQ;
  assign CLBLL_R_X57Y101_SLICE_X87Y101_C5 = CLBLM_L_X64Y100_SLICE_X97Y100_AQ;
  assign CLBLL_R_X57Y101_SLICE_X87Y101_C6 = CLBLM_L_X62Y101_SLICE_X92Y101_DO6;
  assign CLBLL_R_X57Y101_SLICE_X87Y101_CE = CLBLL_R_X57Y100_SLICE_X87Y100_DO6;
  assign CLBLL_R_X57Y101_SLICE_X87Y101_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X57Y101_SLICE_X87Y101_D1 = CLBLM_L_X56Y100_SLICE_X85Y100_DQ;
  assign CLBLL_R_X57Y101_SLICE_X87Y101_D2 = CLBLM_L_X56Y99_SLICE_X85Y99_BQ;
  assign CLBLL_R_X57Y101_SLICE_X87Y101_D3 = CLBLM_L_X62Y101_SLICE_X93Y101_BQ;
  assign CLBLL_R_X57Y101_SLICE_X87Y101_D4 = CLBLL_L_X54Y99_SLICE_X82Y99_CQ;
  assign CLBLL_R_X57Y101_SLICE_X87Y101_D5 = CLBLM_R_X59Y96_SLICE_X89Y96_AQ;
  assign CLBLL_R_X57Y101_SLICE_X87Y101_D6 = CLBLL_R_X57Y101_SLICE_X87Y101_BO6;
  assign RIOI3_X105Y111_OLOGIC_X1Y112_D1 = CLBLM_R_X65Y100_SLICE_X99Y100_BQ;
  assign CLBLL_R_X57Y101_SLICE_X87Y101_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign RIOI3_X105Y111_OLOGIC_X1Y112_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1 = CLBLM_R_X49Y109_SLICE_X74Y109_DQ;
  assign RIOI3_X105Y111_OLOGIC_X1Y111_D1 = CLBLM_L_X64Y106_SLICE_X97Y106_DQ;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1 = 1'b1;
  assign RIOI3_X105Y111_OLOGIC_X1Y111_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1 = CLBLM_R_X49Y109_SLICE_X74Y109_CQ;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1 = 1'b1;
  assign CLBLM_L_X56Y101_SLICE_X85Y101_A1 = CLBLM_L_X60Y101_SLICE_X91Y101_CO6;
  assign CLBLM_L_X56Y101_SLICE_X85Y101_A2 = CLBLM_R_X59Y98_SLICE_X89Y98_BQ;
  assign CLBLM_L_X56Y101_SLICE_X85Y101_A3 = CLBLL_L_X54Y98_SLICE_X83Y98_BQ;
  assign CLBLM_L_X56Y101_SLICE_X85Y101_A4 = 1'b1;
  assign CLBLM_L_X56Y101_SLICE_X85Y101_A5 = CLBLL_L_X54Y101_SLICE_X82Y101_AQ;
  assign CLBLM_L_X56Y101_SLICE_X85Y101_A6 = CLBLL_L_X54Y99_SLICE_X82Y99_AQ;
  assign CLBLM_L_X56Y101_SLICE_X85Y101_B1 = 1'b1;
  assign CLBLM_L_X56Y101_SLICE_X85Y101_B2 = CLBLM_R_X59Y98_SLICE_X89Y98_C5Q;
  assign CLBLM_L_X56Y101_SLICE_X85Y101_B3 = CLBLL_L_X54Y98_SLICE_X83Y98_BQ;
  assign CLBLM_L_X56Y101_SLICE_X85Y101_B4 = CLBLM_L_X56Y100_SLICE_X85Y100_CQ;
  assign CLBLM_L_X56Y101_SLICE_X85Y101_B5 = CLBLM_L_X62Y101_SLICE_X92Y101_DO5;
  assign CLBLM_L_X56Y101_SLICE_X85Y101_B6 = CLBLL_L_X54Y99_SLICE_X82Y99_AQ;
  assign CLBLL_R_X57Y102_SLICE_X86Y102_A1 = CLBLM_R_X49Y104_SLICE_X75Y104_AQ;
  assign CLBLL_R_X57Y102_SLICE_X86Y102_A2 = CLBLL_R_X57Y102_SLICE_X86Y102_DO6;
  assign CLBLL_R_X57Y102_SLICE_X86Y102_A3 = CLBLM_L_X56Y102_SLICE_X85Y102_BO6;
  assign CLBLL_R_X57Y102_SLICE_X86Y102_A4 = 1'b1;
  assign CLBLM_L_X56Y101_SLICE_X85Y101_C4 = CLBLM_L_X56Y99_SLICE_X85Y99_BQ;
  assign CLBLM_L_X56Y101_SLICE_X85Y101_C5 = CLBLM_L_X60Y101_SLICE_X91Y101_CO6;
  assign CLBLM_L_X56Y101_SLICE_X85Y101_C6 = CLBLM_R_X59Y98_SLICE_X89Y98_BQ;
  assign CLBLL_R_X57Y102_SLICE_X86Y102_A5 = CLBLL_R_X57Y102_SLICE_X86Y102_CO6;
  assign CLBLL_R_X57Y102_SLICE_X86Y102_A6 = 1'b1;
  assign CLBLM_L_X56Y101_SLICE_X85Y101_C1 = CLBLL_L_X54Y101_SLICE_X82Y101_AQ;
  assign CLBLM_L_X56Y101_SLICE_X85Y101_C2 = CLBLL_L_X54Y99_SLICE_X82Y99_CQ;
  assign CLBLL_R_X57Y102_SLICE_X86Y102_AX = CLBLL_R_X57Y102_SLICE_X86Y102_DO6;
  assign CLBLM_L_X56Y101_SLICE_X85Y101_C3 = CLBLM_L_X62Y101_SLICE_X93Y101_AQ;
  assign CLBLL_R_X57Y102_SLICE_X86Y102_B1 = CLBLL_R_X57Y102_SLICE_X86Y102_DO6;
  assign CLBLL_R_X57Y102_SLICE_X86Y102_B2 = 1'b1;
  assign CLBLL_R_X57Y102_SLICE_X86Y102_B3 = 1'b1;
  assign CLBLM_L_X56Y101_SLICE_X85Y101_D1 = CLBLM_L_X62Y101_SLICE_X92Y101_DO5;
  assign CLBLM_L_X56Y101_SLICE_X85Y101_D2 = CLBLL_L_X54Y99_SLICE_X82Y99_CQ;
  assign CLBLL_R_X57Y102_SLICE_X86Y102_B4 = 1'b1;
  assign CLBLM_L_X56Y101_SLICE_X85Y101_D4 = CLBLM_L_X56Y100_SLICE_X85Y100_CQ;
  assign CLBLM_L_X56Y101_SLICE_X85Y101_D5 = CLBLM_L_X64Y100_SLICE_X97Y100_BQ;
  assign CLBLM_L_X56Y101_SLICE_X85Y101_D6 = CLBLM_R_X59Y98_SLICE_X89Y98_C5Q;
  assign CLBLL_R_X57Y102_SLICE_X86Y102_B5 = 1'b1;
  assign CLBLL_R_X57Y102_SLICE_X86Y102_B6 = CLBLM_R_X49Y104_SLICE_X75Y104_BQ;
  assign CLBLM_L_X56Y101_SLICE_X85Y101_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLL_R_X57Y102_SLICE_X86Y102_C1 = CLBLM_R_X49Y106_SLICE_X75Y106_CQ;
  assign CLBLL_R_X57Y102_SLICE_X86Y102_C2 = CLBLM_R_X49Y106_SLICE_X75Y106_DQ;
  assign CLBLL_R_X57Y102_SLICE_X86Y102_C3 = CLBLM_R_X49Y104_SLICE_X75Y104_CQ;
  assign CLBLL_R_X57Y102_SLICE_X86Y102_C4 = CLBLM_R_X49Y104_SLICE_X75Y104_BQ;
  assign CLBLL_R_X57Y102_SLICE_X86Y102_C5 = CLBLM_R_X49Y104_SLICE_X75Y104_DQ;
  assign CLBLL_R_X57Y102_SLICE_X86Y102_C6 = CLBLM_R_X49Y107_SLICE_X75Y107_CQ;
  assign CLBLL_R_X57Y102_SLICE_X86Y102_CE = CLBLM_L_X60Y98_SLICE_X91Y98_DQ;
  assign CLBLL_R_X57Y102_SLICE_X86Y102_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X56Y101_SLICE_X84Y101_A1 = CLBLM_L_X56Y102_SLICE_X85Y102_A5Q;
  assign CLBLM_L_X56Y101_SLICE_X84Y101_A2 = 1'b1;
  assign CLBLM_L_X56Y101_SLICE_X84Y101_A3 = CLBLM_L_X56Y101_SLICE_X84Y101_AQ;
  assign CLBLM_L_X56Y101_SLICE_X84Y101_A4 = 1'b1;
  assign CLBLM_L_X56Y101_SLICE_X84Y101_A5 = CLBLM_L_X56Y102_SLICE_X85Y102_AQ;
  assign CLBLL_R_X57Y102_SLICE_X86Y102_D1 = CLBLM_R_X49Y106_SLICE_X75Y106_CQ;
  assign CLBLL_R_X57Y102_SLICE_X86Y102_D2 = CLBLM_R_X49Y106_SLICE_X75Y106_DQ;
  assign CLBLL_R_X57Y102_SLICE_X86Y102_D3 = CLBLM_R_X49Y104_SLICE_X75Y104_DQ;
  assign CLBLL_R_X57Y102_SLICE_X86Y102_D4 = CLBLM_R_X49Y104_SLICE_X75Y104_CQ;
  assign CLBLL_R_X57Y102_SLICE_X86Y102_D5 = CLBLM_R_X49Y107_SLICE_X75Y107_CQ;
  assign CLBLL_R_X57Y102_SLICE_X86Y102_D6 = CLBLM_L_X56Y100_SLICE_X85Y100_BO6;
  assign CLBLM_L_X56Y101_SLICE_X84Y101_AX = 1'b0;
  assign CLBLL_R_X57Y102_SLICE_X86Y102_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X56Y101_SLICE_X84Y101_B2 = CLBLM_L_X56Y101_SLICE_X84Y101_BQ;
  assign CLBLM_L_X56Y101_SLICE_X84Y101_B3 = CLBLM_L_X56Y102_SLICE_X85Y102_AQ;
  assign CLBLM_L_X56Y101_SLICE_X84Y101_B4 = 1'b1;
  assign CLBLM_L_X56Y101_SLICE_X84Y101_B5 = 1'b1;
  assign CLBLM_L_X56Y101_SLICE_X84Y101_B6 = 1'b1;
  assign CLBLM_L_X56Y101_SLICE_X84Y101_BX = 1'b0;
  assign CLBLM_L_X56Y101_SLICE_X84Y101_C1 = CLBLM_L_X56Y102_SLICE_X85Y102_AQ;
  assign CLBLM_L_X56Y101_SLICE_X84Y101_C2 = CLBLM_L_X56Y101_SLICE_X84Y101_CQ;
  assign CLBLM_L_X56Y101_SLICE_X84Y101_C3 = 1'b1;
  assign CLBLM_L_X56Y101_SLICE_X84Y101_C4 = 1'b1;
  assign CLBLM_L_X56Y101_SLICE_X84Y101_C5 = CLBLM_L_X56Y102_SLICE_X85Y102_A5Q;
  assign CLBLM_L_X56Y101_SLICE_X84Y101_C6 = 1'b1;
  assign CLBLM_L_X56Y101_SLICE_X84Y101_CE = CLBLM_L_X56Y102_SLICE_X85Y102_CO6;
  assign CLBLM_L_X56Y101_SLICE_X84Y101_CIN = CLBLM_L_X56Y100_SLICE_X84Y100_COUT;
  assign CLBLM_L_X56Y101_SLICE_X84Y101_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X56Y101_SLICE_X84Y101_CX = 1'b0;
  assign CLBLM_L_X56Y101_SLICE_X84Y101_D1 = CLBLM_L_X56Y102_SLICE_X85Y102_AQ;
  assign CLBLM_L_X56Y101_SLICE_X84Y101_D2 = 1'b1;
  assign CLBLM_L_X56Y101_SLICE_X84Y101_D3 = CLBLM_L_X56Y101_SLICE_X84Y101_DQ;
  assign CLBLL_R_X57Y102_SLICE_X87Y102_A1 = 1'b1;
  assign CLBLL_R_X57Y102_SLICE_X87Y102_A2 = 1'b1;
  assign CLBLL_R_X57Y102_SLICE_X87Y102_A3 = 1'b1;
  assign CLBLL_R_X57Y102_SLICE_X87Y102_A4 = 1'b1;
  assign CLBLL_R_X57Y102_SLICE_X87Y102_A5 = 1'b1;
  assign CLBLL_R_X57Y102_SLICE_X87Y102_A6 = 1'b1;
  assign CLBLM_L_X56Y101_SLICE_X84Y101_DX = 1'b0;
  assign CLBLM_L_X56Y101_SLICE_X84Y101_D4 = 1'b1;
  assign CLBLM_L_X56Y101_SLICE_X84Y101_D5 = CLBLM_L_X56Y102_SLICE_X85Y102_A5Q;
  assign CLBLM_L_X56Y101_SLICE_X84Y101_D6 = 1'b1;
  assign CLBLL_R_X57Y102_SLICE_X87Y102_B1 = 1'b1;
  assign CLBLL_R_X57Y102_SLICE_X87Y102_B2 = 1'b1;
  assign CLBLL_R_X57Y102_SLICE_X87Y102_B3 = 1'b1;
  assign CLBLL_R_X57Y102_SLICE_X87Y102_B4 = 1'b1;
  assign CLBLL_R_X57Y102_SLICE_X87Y102_B5 = 1'b1;
  assign CLBLL_R_X57Y102_SLICE_X87Y102_B6 = 1'b1;
  assign CLBLL_R_X57Y102_SLICE_X87Y102_C1 = 1'b1;
  assign CLBLL_R_X57Y102_SLICE_X87Y102_C2 = 1'b1;
  assign CLBLL_R_X57Y102_SLICE_X87Y102_C3 = 1'b1;
  assign CLBLL_R_X57Y102_SLICE_X87Y102_C4 = 1'b1;
  assign CLBLL_R_X57Y102_SLICE_X87Y102_C5 = 1'b1;
  assign CLBLL_R_X57Y102_SLICE_X87Y102_C6 = 1'b1;
  assign CLBLL_R_X57Y102_SLICE_X87Y102_D1 = 1'b1;
  assign CLBLL_R_X57Y102_SLICE_X87Y102_D2 = 1'b1;
  assign CLBLL_R_X57Y102_SLICE_X87Y102_D3 = 1'b1;
  assign CLBLL_R_X57Y102_SLICE_X87Y102_D4 = 1'b1;
  assign CLBLL_R_X57Y102_SLICE_X87Y102_D5 = 1'b1;
  assign CLBLL_R_X57Y102_SLICE_X87Y102_D6 = 1'b1;
  assign RIOI3_X105Y117_OLOGIC_X1Y118_D1 = CLBLM_R_X65Y107_SLICE_X98Y107_AQ;
  assign CLBLM_L_X56Y102_SLICE_X85Y102_A1 = 1'b1;
  assign CLBLM_L_X56Y102_SLICE_X85Y102_A2 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_L_X56Y102_SLICE_X85Y102_A3 = CLBLM_L_X56Y98_SLICE_X85Y98_AQ;
  assign CLBLM_L_X56Y102_SLICE_X85Y102_A4 = CLBLM_L_X60Y98_SLICE_X91Y98_DQ;
  assign CLBLM_L_X56Y102_SLICE_X85Y102_A5 = CLBLM_L_X56Y99_SLICE_X85Y99_CQ;
  assign CLBLM_L_X56Y102_SLICE_X85Y102_A6 = 1'b1;
  assign CLBLM_L_X56Y102_SLICE_X85Y102_B1 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLM_L_X56Y102_SLICE_X85Y102_B2 = CLBLM_R_X49Y104_SLICE_X74Y104_AQ;
  assign CLBLM_L_X56Y102_SLICE_X85Y102_B3 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLM_L_X56Y102_SLICE_X85Y102_B4 = CLBLM_L_X56Y97_SLICE_X84Y97_CO5;
  assign CLBLL_R_X57Y103_SLICE_X86Y103_A1 = CLBLM_R_X49Y119_SLICE_X74Y119_BQ;
  assign CLBLL_R_X57Y103_SLICE_X86Y103_A2 = CLBLL_R_X57Y103_SLICE_X86Y103_A5Q;
  assign CLBLL_R_X57Y103_SLICE_X86Y103_A3 = CLBLL_R_X57Y103_SLICE_X86Y103_AQ;
  assign CLBLL_R_X57Y103_SLICE_X86Y103_A4 = CLBLM_L_X60Y98_SLICE_X91Y98_DQ;
  assign CLBLL_R_X57Y103_SLICE_X86Y103_A5 = CLBLM_R_X49Y119_SLICE_X74Y119_AQ;
  assign CLBLL_R_X57Y103_SLICE_X86Y103_A6 = 1'b1;
  assign CLBLM_L_X56Y102_SLICE_X85Y102_C1 = CLBLM_R_X63Y100_SLICE_X94Y100_AQ;
  assign CLBLM_L_X56Y102_SLICE_X85Y102_B5 = CLBLM_R_X49Y107_SLICE_X75Y107_DQ;
  assign CLBLM_L_X56Y102_SLICE_X85Y102_B6 = CLBLM_R_X49Y108_SLICE_X75Y108_DQ;
  assign CLBLM_L_X56Y102_SLICE_X85Y102_C4 = CLBLM_L_X56Y102_SLICE_X85Y102_A5Q;
  assign CLBLM_L_X56Y102_SLICE_X85Y102_C6 = 1'b1;
  assign CLBLL_R_X57Y103_SLICE_X86Y103_B1 = 1'b1;
  assign CLBLM_L_X56Y102_SLICE_X85Y102_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X57Y103_SLICE_X86Y103_B2 = 1'b1;
  assign CLBLL_R_X57Y103_SLICE_X86Y103_B3 = 1'b1;
  assign CLBLL_R_X57Y103_SLICE_X86Y103_B4 = 1'b1;
  assign CLBLL_R_X57Y103_SLICE_X86Y103_B5 = 1'b1;
  assign CLBLL_R_X57Y103_SLICE_X86Y103_B6 = 1'b1;
  assign CLBLL_R_X57Y103_SLICE_X86Y103_C1 = 1'b1;
  assign CLBLL_R_X57Y103_SLICE_X86Y103_C2 = 1'b1;
  assign CLBLL_R_X57Y103_SLICE_X86Y103_C3 = 1'b1;
  assign CLBLL_R_X57Y103_SLICE_X86Y103_C4 = 1'b1;
  assign CLBLL_R_X57Y103_SLICE_X86Y103_C5 = 1'b1;
  assign CLBLM_L_X56Y102_SLICE_X85Y102_D6 = 1'b1;
  assign CLBLL_R_X57Y103_SLICE_X86Y103_C6 = 1'b1;
  assign CLBLM_L_X56Y102_SLICE_X85Y102_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLL_R_X57Y103_SLICE_X86Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X56Y102_SLICE_X85Y102_D3 = 1'b1;
  assign CLBLM_L_X56Y102_SLICE_X85Y102_D4 = 1'b1;
  assign CLBLM_L_X56Y102_SLICE_X85Y102_D5 = 1'b1;
  assign CLBLM_L_X56Y102_SLICE_X84Y102_A1 = 1'b1;
  assign CLBLL_R_X57Y103_SLICE_X86Y103_D1 = 1'b1;
  assign CLBLL_R_X57Y103_SLICE_X86Y103_D2 = 1'b1;
  assign CLBLL_R_X57Y103_SLICE_X86Y103_D3 = 1'b1;
  assign CLBLL_R_X57Y103_SLICE_X86Y103_D4 = 1'b1;
  assign CLBLL_R_X57Y103_SLICE_X86Y103_D5 = 1'b1;
  assign CLBLL_R_X57Y103_SLICE_X86Y103_D6 = 1'b1;
  assign CLBLM_L_X56Y102_SLICE_X84Y102_A2 = 1'b1;
  assign CLBLM_L_X56Y102_SLICE_X84Y102_A3 = CLBLM_L_X56Y102_SLICE_X84Y102_AQ;
  assign CLBLL_R_X57Y103_SLICE_X86Y103_SR = CLBLM_R_X15Y122_SLICE_X20Y122_AO6;
  assign CLBLM_L_X56Y102_SLICE_X84Y102_A5 = CLBLM_L_X56Y102_SLICE_X85Y102_AQ;
  assign CLBLM_L_X56Y102_SLICE_X84Y102_A6 = 1'b1;
  assign CLBLM_L_X56Y102_SLICE_X84Y102_AX = 1'b0;
  assign CLBLM_L_X56Y102_SLICE_X84Y102_B1 = 1'b1;
  assign CLBLM_L_X56Y102_SLICE_X84Y102_B2 = CLBLM_L_X56Y102_SLICE_X84Y102_BQ;
  assign CLBLM_L_X56Y102_SLICE_X84Y102_B3 = CLBLM_L_X56Y102_SLICE_X85Y102_A5Q;
  assign CLBLM_L_X56Y102_SLICE_X84Y102_B4 = 1'b1;
  assign CLBLM_L_X56Y102_SLICE_X84Y102_B5 = CLBLM_L_X56Y102_SLICE_X85Y102_AQ;
  assign CLBLM_L_X56Y102_SLICE_X84Y102_B6 = 1'b1;
  assign CLBLM_L_X56Y102_SLICE_X84Y102_BX = 1'b0;
  assign CLBLM_L_X56Y102_SLICE_X84Y102_C1 = CLBLM_L_X56Y102_SLICE_X85Y102_AQ;
  assign CLBLM_L_X56Y102_SLICE_X84Y102_C2 = CLBLM_L_X56Y102_SLICE_X84Y102_CQ;
  assign CLBLM_L_X56Y102_SLICE_X84Y102_C3 = 1'b1;
  assign CLBLM_L_X56Y102_SLICE_X84Y102_C4 = 1'b1;
  assign CLBLM_L_X56Y102_SLICE_X84Y102_C5 = 1'b1;
  assign CLBLM_L_X56Y102_SLICE_X84Y102_C6 = CLBLM_L_X56Y102_SLICE_X85Y102_A5Q;
  assign CLBLM_L_X56Y102_SLICE_X84Y102_CE = CLBLM_L_X56Y102_SLICE_X85Y102_CO6;
  assign CLBLM_L_X56Y102_SLICE_X84Y102_CIN = CLBLM_L_X56Y101_SLICE_X84Y101_COUT;
  assign CLBLM_L_X56Y102_SLICE_X84Y102_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X57Y103_SLICE_X87Y103_A1 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLL_R_X57Y103_SLICE_X87Y103_A2 = CLBLL_R_X57Y105_SLICE_X87Y105_D_XOR;
  assign CLBLL_R_X57Y103_SLICE_X87Y103_A3 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLL_R_X57Y103_SLICE_X87Y103_A4 = CLBLL_R_X57Y106_SLICE_X86Y106_D_XOR;
  assign CLBLM_L_X56Y102_SLICE_X84Y102_D3 = CLBLM_L_X56Y102_SLICE_X84Y102_DQ;
  assign CLBLM_L_X56Y102_SLICE_X84Y102_D4 = 1'b1;
  assign CLBLM_L_X56Y102_SLICE_X84Y102_D5 = 1'b1;
  assign CLBLL_R_X57Y103_SLICE_X87Y103_A5 = CLBLM_L_X62Y102_SLICE_X92Y102_AO5;
  assign CLBLL_R_X57Y103_SLICE_X87Y103_A6 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_L_X56Y102_SLICE_X84Y102_CX = 1'b0;
  assign CLBLM_L_X56Y102_SLICE_X84Y102_D1 = CLBLM_L_X56Y102_SLICE_X85Y102_AQ;
  assign CLBLM_L_X56Y102_SLICE_X84Y102_D2 = CLBLM_L_X56Y102_SLICE_X85Y102_A5Q;
  assign CLBLL_R_X57Y103_SLICE_X87Y103_B1 = 1'b1;
  assign CLBLL_R_X57Y103_SLICE_X87Y103_B2 = 1'b1;
  assign CLBLL_R_X57Y103_SLICE_X87Y103_B3 = 1'b1;
  assign CLBLL_R_X57Y103_SLICE_X87Y103_B4 = 1'b1;
  assign CLBLL_R_X57Y103_SLICE_X87Y103_B5 = 1'b1;
  assign CLBLL_R_X57Y103_SLICE_X87Y103_B6 = 1'b1;
  assign CLBLM_L_X56Y102_SLICE_X84Y102_DX = 1'b0;
  assign CLBLM_L_X56Y102_SLICE_X84Y102_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLL_R_X57Y103_SLICE_X87Y103_C1 = 1'b1;
  assign CLBLL_R_X57Y103_SLICE_X87Y103_C2 = 1'b1;
  assign CLBLL_R_X57Y103_SLICE_X87Y103_C3 = 1'b1;
  assign CLBLL_R_X57Y103_SLICE_X87Y103_C4 = 1'b1;
  assign CLBLL_R_X57Y103_SLICE_X87Y103_C5 = 1'b1;
  assign CLBLL_R_X57Y103_SLICE_X87Y103_C6 = 1'b1;
  assign CLBLL_R_X57Y103_SLICE_X87Y103_CE = CLBLM_L_X60Y100_SLICE_X90Y100_BO6;
  assign CLBLL_R_X57Y103_SLICE_X87Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X57Y103_SLICE_X87Y103_D1 = 1'b1;
  assign CLBLL_R_X57Y103_SLICE_X87Y103_D2 = 1'b1;
  assign CLBLL_R_X57Y103_SLICE_X87Y103_D3 = 1'b1;
  assign CLBLL_R_X57Y103_SLICE_X87Y103_D4 = 1'b1;
  assign CLBLL_R_X57Y103_SLICE_X87Y103_D5 = 1'b1;
  assign CLBLL_R_X57Y103_SLICE_X87Y103_D6 = 1'b1;
  assign CLBLL_R_X57Y103_SLICE_X87Y103_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign RIOI3_X105Y117_OLOGIC_X1Y118_T1 = 1'b1;
  assign RIOI3_X105Y115_OLOGIC_X1Y116_D1 = CLBLM_R_X63Y103_SLICE_X95Y103_CQ;
  assign RIOI3_X105Y115_OLOGIC_X1Y116_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1 = CLBLM_L_X50Y106_SLICE_X76Y106_AQ;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_B3 = 1'b1;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_B4 = 1'b1;
  assign RIOI3_X105Y115_OLOGIC_X1Y115_D1 = CLBLM_R_X63Y101_SLICE_X95Y101_AQ;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_B5 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1 = 1'b1;
  assign RIOI3_X105Y115_OLOGIC_X1Y115_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1 = CLBLM_R_X49Y106_SLICE_X74Y106_AQ;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1 = 1'b1;
  assign CLBLM_L_X56Y103_SLICE_X85Y103_A1 = CLBLM_L_X50Y106_SLICE_X76Y106_AQ;
  assign CLBLM_L_X56Y103_SLICE_X85Y103_A2 = CLBLM_L_X60Y99_SLICE_X90Y99_AO5;
  assign CLBLM_L_X56Y103_SLICE_X85Y103_A3 = CLBLM_L_X56Y103_SLICE_X85Y103_AQ;
  assign CLBLM_L_X56Y103_SLICE_X85Y103_A4 = CLBLL_L_X54Y101_SLICE_X83Y101_BO6;
  assign CLBLM_L_X56Y103_SLICE_X85Y103_A5 = CLBLL_L_X54Y107_SLICE_X82Y107_B_XOR;
  assign CLBLM_L_X56Y103_SLICE_X85Y103_A6 = 1'b1;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_C3 = 1'b1;
  assign CLBLM_R_X65Y106_SLICE_X99Y106_C4 = 1'b1;
  assign CLBLL_R_X57Y104_SLICE_X86Y104_A1 = CLBLL_L_X54Y106_SLICE_X82Y106_B_XOR;
  assign CLBLL_R_X57Y104_SLICE_X86Y104_A2 = 1'b1;
  assign CLBLM_L_X56Y103_SLICE_X85Y103_B2 = CLBLM_L_X56Y103_SLICE_X85Y103_BQ;
  assign CLBLM_L_X56Y103_SLICE_X85Y103_B3 = CLBLM_L_X50Y106_SLICE_X76Y106_AQ;
  assign CLBLM_L_X56Y103_SLICE_X85Y103_B4 = CLBLL_L_X54Y101_SLICE_X83Y101_BO6;
  assign CLBLM_L_X56Y103_SLICE_X85Y103_B5 = CLBLM_L_X62Y100_SLICE_X92Y100_AO5;
  assign CLBLM_L_X56Y103_SLICE_X85Y103_B6 = 1'b1;
  assign CLBLL_R_X57Y104_SLICE_X86Y104_A3 = CLBLL_R_X57Y104_SLICE_X86Y104_AQ;
  assign CLBLL_R_X57Y104_SLICE_X86Y104_A4 = CLBLM_L_X50Y104_SLICE_X76Y104_AQ;
  assign CLBLL_R_X57Y104_SLICE_X86Y104_A5 = CLBLL_L_X54Y101_SLICE_X83Y101_BO6;
  assign CLBLL_R_X57Y104_SLICE_X86Y104_A6 = CLBLM_L_X60Y99_SLICE_X90Y99_AO5;
  assign CLBLM_L_X56Y103_SLICE_X85Y103_C2 = 1'b1;
  assign CLBLM_L_X56Y103_SLICE_X85Y103_C3 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_L_X56Y103_SLICE_X85Y103_C4 = 1'b1;
  assign CLBLM_L_X56Y103_SLICE_X85Y103_C5 = 1'b1;
  assign CLBLM_L_X56Y103_SLICE_X85Y103_C6 = CLBLM_L_X60Y98_SLICE_X91Y98_DQ;
  assign CLBLM_L_X56Y103_SLICE_X85Y103_CE = CLBLM_L_X56Y103_SLICE_X85Y103_CO6;
  assign CLBLL_R_X57Y104_SLICE_X86Y104_B1 = 1'b1;
  assign CLBLL_R_X57Y104_SLICE_X86Y104_B2 = CLBLL_R_X57Y104_SLICE_X86Y104_BQ;
  assign CLBLL_R_X57Y104_SLICE_X86Y104_B3 = CLBLM_L_X62Y100_SLICE_X92Y100_AO5;
  assign CLBLL_R_X57Y104_SLICE_X86Y104_B4 = CLBLM_L_X50Y104_SLICE_X76Y104_AQ;
  assign CLBLL_R_X57Y104_SLICE_X86Y104_B5 = CLBLL_L_X54Y101_SLICE_X83Y101_BO6;
  assign CLBLL_R_X57Y104_SLICE_X86Y104_B6 = CLBLM_R_X53Y103_SLICE_X81Y103_A_XOR;
  assign CLBLL_R_X57Y104_SLICE_X86Y104_C1 = CLBLL_L_X54Y101_SLICE_X83Y101_BO6;
  assign CLBLL_R_X57Y104_SLICE_X86Y104_C2 = CLBLL_R_X57Y104_SLICE_X86Y104_CQ;
  assign CLBLL_R_X57Y104_SLICE_X86Y104_C3 = CLBLM_R_X53Y103_SLICE_X81Y103_B_XOR;
  assign CLBLL_R_X57Y104_SLICE_X86Y104_C4 = 1'b1;
  assign CLBLL_R_X57Y104_SLICE_X86Y104_C5 = CLBLM_L_X50Y105_SLICE_X77Y105_AQ;
  assign CLBLM_L_X56Y103_SLICE_X85Y103_D5 = 1'b1;
  assign CLBLM_L_X56Y103_SLICE_X85Y103_D6 = 1'b1;
  assign CLBLL_R_X57Y104_SLICE_X86Y104_C6 = CLBLM_L_X62Y100_SLICE_X92Y100_AO5;
  assign CLBLL_R_X57Y104_SLICE_X86Y104_CE = CLBLM_L_X56Y103_SLICE_X85Y103_CO6;
  assign CLBLM_L_X56Y103_SLICE_X85Y103_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLL_R_X57Y104_SLICE_X86Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X56Y103_SLICE_X85Y103_D3 = 1'b1;
  assign CLBLL_R_X57Y104_SLICE_X86Y104_D1 = CLBLL_R_X57Y104_SLICE_X86Y104_BQ;
  assign CLBLL_R_X57Y104_SLICE_X86Y104_D2 = CLBLL_R_X57Y104_SLICE_X86Y104_AQ;
  assign CLBLL_R_X57Y104_SLICE_X86Y104_D3 = CLBLL_R_X57Y101_SLICE_X86Y101_AQ;
  assign CLBLL_R_X57Y104_SLICE_X86Y104_D4 = CLBLM_L_X60Y108_SLICE_X91Y108_AQ;
  assign CLBLL_R_X57Y104_SLICE_X86Y104_D5 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLL_R_X57Y104_SLICE_X86Y104_D6 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_L_X56Y103_SLICE_X84Y103_A1 = CLBLM_L_X56Y102_SLICE_X85Y102_AQ;
  assign CLBLM_L_X56Y103_SLICE_X84Y103_A2 = CLBLM_L_X56Y102_SLICE_X85Y102_A5Q;
  assign CLBLL_R_X57Y104_SLICE_X86Y104_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X56Y103_SLICE_X84Y103_A3 = CLBLM_L_X56Y103_SLICE_X84Y103_AQ;
  assign CLBLM_L_X56Y103_SLICE_X84Y103_A4 = 1'b1;
  assign CLBLM_L_X56Y103_SLICE_X84Y103_A5 = 1'b1;
  assign CLBLM_L_X56Y103_SLICE_X84Y103_A6 = 1'b1;
  assign CLBLM_L_X56Y103_SLICE_X84Y103_AX = 1'b0;
  assign CLBLM_L_X56Y103_SLICE_X84Y103_B1 = CLBLM_L_X56Y102_SLICE_X85Y102_AQ;
  assign CLBLM_L_X56Y103_SLICE_X84Y103_B2 = CLBLM_L_X56Y103_SLICE_X84Y103_BQ;
  assign CLBLM_L_X56Y103_SLICE_X84Y103_B3 = CLBLM_L_X56Y102_SLICE_X85Y102_A5Q;
  assign CLBLM_L_X56Y103_SLICE_X84Y103_B4 = 1'b1;
  assign CLBLM_L_X56Y103_SLICE_X84Y103_B5 = 1'b1;
  assign CLBLM_L_X56Y103_SLICE_X84Y103_B6 = 1'b1;
  assign CLBLM_L_X56Y103_SLICE_X84Y103_BX = 1'b0;
  assign CLBLM_L_X56Y103_SLICE_X84Y103_C1 = CLBLM_L_X56Y102_SLICE_X85Y102_A5Q;
  assign CLBLM_L_X56Y103_SLICE_X84Y103_C2 = CLBLM_L_X56Y103_SLICE_X84Y103_CQ;
  assign CLBLM_L_X56Y103_SLICE_X84Y103_C3 = 1'b1;
  assign CLBLM_L_X56Y103_SLICE_X84Y103_C4 = 1'b1;
  assign CLBLM_L_X56Y103_SLICE_X84Y103_C5 = CLBLM_L_X56Y102_SLICE_X85Y102_AQ;
  assign CLBLM_L_X56Y103_SLICE_X84Y103_C6 = 1'b1;
  assign CLBLM_L_X56Y103_SLICE_X84Y103_CE = CLBLM_L_X56Y102_SLICE_X85Y102_CO6;
  assign CLBLM_L_X56Y103_SLICE_X84Y103_CIN = CLBLM_L_X56Y102_SLICE_X84Y102_COUT;
  assign CLBLL_R_X57Y104_SLICE_X87Y104_A1 = 1'b1;
  assign CLBLL_R_X57Y104_SLICE_X87Y104_A2 = CLBLM_L_X60Y99_SLICE_X90Y99_AO5;
  assign CLBLL_R_X57Y104_SLICE_X87Y104_A3 = CLBLL_R_X57Y104_SLICE_X87Y104_AQ;
  assign CLBLL_R_X57Y104_SLICE_X87Y104_A4 = CLBLL_L_X54Y106_SLICE_X82Y106_D_XOR;
  assign CLBLL_R_X57Y104_SLICE_X87Y104_A5 = CLBLL_L_X54Y101_SLICE_X83Y101_BO6;
  assign CLBLL_R_X57Y104_SLICE_X87Y104_A6 = CLBLM_R_X49Y105_SLICE_X75Y105_CQ;
  assign CLBLM_L_X56Y103_SLICE_X84Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X56Y103_SLICE_X84Y103_CX = 1'b0;
  assign CLBLM_L_X56Y103_SLICE_X84Y103_D1 = CLBLM_L_X56Y102_SLICE_X85Y102_A5Q;
  assign CLBLL_R_X57Y104_SLICE_X87Y104_B1 = CLBLM_L_X60Y99_SLICE_X90Y99_AO5;
  assign CLBLM_L_X56Y103_SLICE_X84Y103_D5 = CLBLM_L_X56Y102_SLICE_X85Y102_AQ;
  assign CLBLM_L_X56Y103_SLICE_X84Y103_D6 = 1'b1;
  assign CLBLL_R_X57Y104_SLICE_X87Y104_B2 = CLBLL_R_X57Y104_SLICE_X87Y104_BQ;
  assign CLBLL_R_X57Y104_SLICE_X87Y104_B3 = CLBLL_L_X54Y101_SLICE_X83Y101_BO6;
  assign CLBLL_R_X57Y104_SLICE_X87Y104_B4 = 1'b1;
  assign CLBLM_L_X56Y103_SLICE_X84Y103_DX = 1'b0;
  assign CLBLM_L_X56Y103_SLICE_X84Y103_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLL_R_X57Y104_SLICE_X87Y104_B5 = CLBLL_L_X54Y108_SLICE_X82Y108_A_XOR;
  assign CLBLL_R_X57Y104_SLICE_X87Y104_B6 = CLBLM_L_X50Y107_SLICE_X77Y107_AQ;
  assign CLBLL_R_X57Y104_SLICE_X87Y104_C1 = CLBLL_L_X54Y101_SLICE_X83Y101_BO6;
  assign CLBLL_R_X57Y104_SLICE_X87Y104_C2 = CLBLL_R_X57Y104_SLICE_X87Y104_CQ;
  assign CLBLL_R_X57Y104_SLICE_X87Y104_C3 = CLBLM_R_X53Y103_SLICE_X81Y103_C_XOR;
  assign CLBLL_R_X57Y104_SLICE_X87Y104_C4 = CLBLM_R_X49Y105_SLICE_X75Y105_CQ;
  assign CLBLL_R_X57Y104_SLICE_X87Y104_C5 = 1'b1;
  assign CLBLL_R_X57Y104_SLICE_X87Y104_C6 = CLBLM_L_X62Y100_SLICE_X92Y100_AO5;
  assign CLBLL_R_X57Y104_SLICE_X87Y104_CE = CLBLM_L_X56Y103_SLICE_X85Y103_CO6;
  assign CLBLL_R_X57Y104_SLICE_X87Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X57Y104_SLICE_X87Y104_D1 = CLBLL_R_X57Y105_SLICE_X86Y105_AQ;
  assign CLBLL_R_X57Y104_SLICE_X87Y104_D2 = CLBLL_R_X57Y104_SLICE_X87Y104_CQ;
  assign CLBLL_R_X57Y104_SLICE_X87Y104_D3 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLL_R_X57Y104_SLICE_X87Y104_D4 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLL_R_X57Y104_SLICE_X87Y104_D5 = CLBLL_R_X57Y104_SLICE_X87Y104_AQ;
  assign CLBLL_R_X57Y104_SLICE_X87Y104_D6 = CLBLL_R_X57Y109_SLICE_X86Y109_BQ;
  assign CLBLL_R_X57Y104_SLICE_X87Y104_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X59Y96_SLICE_X89Y96_A5 = CLBLM_L_X60Y96_SLICE_X90Y96_BQ;
  assign CLBLM_R_X59Y96_SLICE_X89Y96_A6 = 1'b1;
  assign CLBLM_R_X59Y96_SLICE_X89Y96_B6 = CLBLM_R_X59Y97_SLICE_X89Y97_A5Q;
  assign CLBLM_R_X59Y96_SLICE_X89Y96_C1 = 1'b1;
  assign CLBLM_R_X59Y96_SLICE_X89Y96_C2 = 1'b1;
  assign CLBLM_R_X59Y96_SLICE_X89Y96_C3 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X85Y104_A1 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X85Y104_A2 = CLBLM_L_X62Y100_SLICE_X92Y100_AO5;
  assign CLBLM_L_X56Y104_SLICE_X85Y104_A3 = CLBLM_L_X56Y104_SLICE_X85Y104_AQ;
  assign CLBLM_L_X56Y104_SLICE_X85Y104_A4 = CLBLL_L_X54Y101_SLICE_X83Y101_BO6;
  assign CLBLM_L_X56Y104_SLICE_X85Y104_A5 = CLBLM_L_X50Y107_SLICE_X77Y107_AQ;
  assign CLBLM_L_X56Y104_SLICE_X85Y104_A6 = CLBLL_L_X54Y106_SLICE_X82Y106_A_XOR;
  assign CLBLL_R_X57Y105_SLICE_X86Y105_A1 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLL_R_X57Y105_SLICE_X86Y105_A2 = CLBLM_L_X62Y105_SLICE_X92Y105_AO6;
  assign CLBLL_R_X57Y105_SLICE_X86Y105_A3 = CLBLL_R_X57Y105_SLICE_X87Y105_B_XOR;
  assign CLBLM_L_X56Y104_SLICE_X85Y104_B1 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X85Y104_B2 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X85Y104_B3 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X85Y104_B4 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X85Y104_B5 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X85Y104_B6 = 1'b1;
  assign CLBLL_R_X57Y105_SLICE_X86Y105_A4 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLL_R_X57Y105_SLICE_X86Y105_A5 = CLBLL_R_X57Y106_SLICE_X86Y106_B_XOR;
  assign CLBLL_R_X57Y105_SLICE_X86Y105_B3 = CLBLL_R_X57Y105_SLICE_X87Y105_C_XOR;
  assign CLBLM_L_X56Y104_SLICE_X85Y104_C1 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X85Y104_C2 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X85Y104_C3 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X85Y104_C4 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X85Y104_C5 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X85Y104_C6 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X85Y104_CE = CLBLM_L_X56Y103_SLICE_X85Y103_CO6;
  assign CLBLM_L_X56Y104_SLICE_X85Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X57Y105_SLICE_X86Y105_C1 = CLBLM_L_X56Y105_SLICE_X85Y105_AQ;
  assign CLBLL_R_X57Y105_SLICE_X86Y105_C2 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLL_R_X57Y105_SLICE_X86Y105_C3 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLL_R_X57Y105_SLICE_X86Y105_C4 = CLBLL_R_X57Y104_SLICE_X86Y104_CQ;
  assign CLBLL_R_X57Y105_SLICE_X86Y105_C5 = CLBLM_R_X59Y106_SLICE_X88Y106_BQ;
  assign CLBLM_L_X56Y104_SLICE_X85Y104_D1 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X85Y104_D2 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X85Y104_D3 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X85Y104_D4 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X85Y104_D5 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X85Y104_D6 = 1'b1;
  assign CLBLL_R_X57Y105_SLICE_X86Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X56Y104_SLICE_X85Y104_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLL_R_X57Y105_SLICE_X86Y105_D1 = CLBLL_R_X57Y105_SLICE_X86Y105_BQ;
  assign CLBLL_R_X57Y105_SLICE_X86Y105_D2 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLL_R_X57Y105_SLICE_X86Y105_D3 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLL_R_X57Y105_SLICE_X86Y105_D6 = CLBLM_L_X56Y105_SLICE_X85Y105_DQ;
  assign CLBLL_R_X57Y105_SLICE_X86Y105_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X56Y104_SLICE_X84Y104_A1 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X84Y104_A2 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X84Y104_A6 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X84Y104_A3 = CLBLM_L_X56Y104_SLICE_X84Y104_AQ;
  assign CLBLM_L_X56Y104_SLICE_X84Y104_A4 = CLBLM_L_X56Y102_SLICE_X85Y102_AQ;
  assign CLBLM_L_X56Y104_SLICE_X84Y104_A5 = CLBLM_L_X56Y102_SLICE_X85Y102_A5Q;
  assign CLBLM_L_X56Y104_SLICE_X84Y104_AX = 1'b0;
  assign CLBLM_R_X63Y94_SLICE_X95Y94_A1 = CLBLM_L_X56Y98_SLICE_X85Y98_DQ;
  assign CLBLM_L_X56Y104_SLICE_X84Y104_B1 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X84Y104_B2 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X84Y104_B3 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X84Y104_B4 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X84Y104_B5 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X84Y104_B6 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X95Y94_A3 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X63Y94_SLICE_X95Y94_A4 = CLBLM_L_X50Y104_SLICE_X76Y104_AQ;
  assign CLBLM_R_X63Y94_SLICE_X95Y94_A5 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X84Y104_BX = 1'b0;
  assign CLBLM_L_X56Y104_SLICE_X84Y104_C1 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X84Y104_C2 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X84Y104_C3 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X84Y104_C4 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X84Y104_C5 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X84Y104_C6 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X84Y104_CE = CLBLM_L_X56Y102_SLICE_X85Y102_CO6;
  assign CLBLL_R_X57Y105_SLICE_X87Y105_A1 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X84Y104_CIN = CLBLM_L_X56Y103_SLICE_X84Y103_COUT;
  assign CLBLM_L_X56Y104_SLICE_X84Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X57Y105_SLICE_X87Y105_A2 = 1'b1;
  assign CLBLL_R_X57Y105_SLICE_X87Y105_A3 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X95Y94_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLL_R_X57Y105_SLICE_X87Y105_A4 = CLBLM_R_X59Y106_SLICE_X88Y106_BQ;
  assign CLBLL_R_X57Y105_SLICE_X87Y105_A5 = 1'b1;
  assign CLBLL_R_X57Y105_SLICE_X87Y105_A6 = 1'b1;
  assign CLBLL_R_X57Y105_SLICE_X87Y105_AX = CLBLL_R_X57Y101_SLICE_X86Y101_AQ;
  assign CLBLM_L_X56Y104_SLICE_X84Y104_D3 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X95Y94_D1 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X95Y94_D2 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X95Y94_D3 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X84Y104_D4 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X95Y94_D5 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X95Y94_D6 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X84Y104_D5 = 1'b1;
  assign CLBLM_L_X56Y104_SLICE_X84Y104_D6 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X95Y94_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLL_R_X57Y105_SLICE_X87Y105_BX = CLBLL_R_X57Y105_SLICE_X86Y105_AQ;
  assign CLBLL_R_X57Y105_SLICE_X87Y105_C1 = 1'b1;
  assign CLBLL_R_X57Y105_SLICE_X87Y105_C2 = 1'b1;
  assign CLBLL_R_X57Y105_SLICE_X87Y105_C3 = 1'b1;
  assign CLBLL_R_X57Y105_SLICE_X87Y105_C4 = 1'b1;
  assign CLBLL_R_X57Y105_SLICE_X87Y105_C5 = 1'b1;
  assign CLBLL_R_X57Y105_SLICE_X87Y105_C6 = CLBLL_R_X57Y105_SLICE_X86Y105_BQ;
  assign CLBLM_R_X63Y94_SLICE_X94Y94_A1 = CLBLM_L_X56Y98_SLICE_X85Y98_DQ;
  assign CLBLM_R_X63Y94_SLICE_X94Y94_A2 = CLBLM_L_X50Y107_SLICE_X77Y107_AQ;
  assign CLBLL_R_X57Y105_SLICE_X87Y105_CX = CLBLL_R_X57Y105_SLICE_X86Y105_BQ;
  assign CLBLM_R_X63Y94_SLICE_X94Y94_A3 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLL_R_X57Y105_SLICE_X87Y105_D1 = CLBLL_R_X57Y103_SLICE_X87Y103_AQ;
  assign CLBLL_R_X57Y105_SLICE_X87Y105_D2 = 1'b1;
  assign CLBLL_R_X57Y105_SLICE_X87Y105_D3 = 1'b1;
  assign CLBLL_R_X57Y105_SLICE_X87Y105_D4 = 1'b1;
  assign CLBLL_R_X57Y105_SLICE_X87Y105_D5 = 1'b1;
  assign CLBLL_R_X57Y105_SLICE_X87Y105_D6 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X94Y94_A6 = CLBLM_R_X63Y96_SLICE_X94Y96_BO6;
  assign CLBLL_R_X57Y105_SLICE_X87Y105_DX = CLBLL_R_X57Y103_SLICE_X87Y103_AQ;
  assign CLBLM_R_X63Y94_SLICE_X94Y94_B1 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X94Y94_B2 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X94Y94_B3 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X94Y94_B4 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X94Y94_B5 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X94Y94_B6 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X94Y94_C1 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X94Y94_C2 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X94Y94_C3 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X94Y94_C4 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X94Y94_C5 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X94Y94_C6 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X94Y94_CE = CLBLM_L_X62Y99_SLICE_X93Y99_AO6;
  assign CLBLM_R_X63Y94_SLICE_X94Y94_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X63Y94_SLICE_X94Y94_D1 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X94Y94_D2 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X94Y94_D3 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X94Y94_D4 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X94Y94_D5 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X94Y94_D6 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X94Y94_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE = 1'b1;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_CE = 1'b1;
  assign CLBLL_R_X57Y106_SLICE_X86Y106_A1 = 1'b1;
  assign CLBLM_L_X56Y105_SLICE_X85Y105_A1 = CLBLL_L_X54Y101_SLICE_X83Y101_BO6;
  assign CLBLM_L_X56Y105_SLICE_X85Y105_A2 = CLBLM_L_X60Y99_SLICE_X90Y99_AO5;
  assign CLBLM_L_X56Y105_SLICE_X85Y105_A3 = CLBLM_L_X56Y105_SLICE_X85Y105_AQ;
  assign CLBLM_L_X56Y105_SLICE_X85Y105_A4 = CLBLM_L_X50Y105_SLICE_X77Y105_AQ;
  assign CLBLM_L_X56Y105_SLICE_X85Y105_A5 = 1'b1;
  assign CLBLM_L_X56Y105_SLICE_X85Y105_A6 = CLBLL_L_X54Y106_SLICE_X82Y106_C_XOR;
  assign CLBLL_R_X57Y106_SLICE_X86Y106_A2 = 1'b1;
  assign CLBLL_R_X57Y106_SLICE_X86Y106_A3 = 1'b1;
  assign CLBLL_R_X57Y106_SLICE_X86Y106_A4 = CLBLM_R_X59Y106_SLICE_X88Y106_BQ;
  assign CLBLM_L_X56Y105_SLICE_X85Y105_B1 = 1'b1;
  assign CLBLM_L_X56Y105_SLICE_X85Y105_B2 = CLBLM_L_X56Y105_SLICE_X85Y105_BQ;
  assign CLBLM_L_X56Y105_SLICE_X85Y105_B3 = CLBLL_L_X54Y101_SLICE_X83Y101_BO6;
  assign CLBLM_L_X56Y105_SLICE_X85Y105_B4 = CLBLM_L_X50Y106_SLICE_X76Y106_CQ;
  assign CLBLM_L_X56Y105_SLICE_X85Y105_B5 = CLBLM_L_X62Y100_SLICE_X92Y100_AO5;
  assign CLBLM_L_X56Y105_SLICE_X85Y105_B6 = CLBLL_L_X54Y105_SLICE_X82Y105_C_XOR;
  assign CLBLL_R_X57Y106_SLICE_X86Y106_AX = CLBLL_R_X57Y101_SLICE_X86Y101_AQ;
  assign CLBLL_R_X57Y106_SLICE_X86Y106_B1 = 1'b1;
  assign CLBLL_R_X57Y106_SLICE_X86Y106_B2 = 1'b1;
  assign CLBLL_R_X57Y106_SLICE_X86Y106_B3 = 1'b1;
  assign CLBLL_R_X57Y106_SLICE_X86Y106_B4 = 1'b1;
  assign CLBLL_R_X57Y106_SLICE_X86Y106_B5 = 1'b1;
  assign CLBLM_L_X56Y105_SLICE_X85Y105_C3 = 1'b1;
  assign CLBLM_L_X56Y105_SLICE_X85Y105_C4 = CLBLL_L_X54Y101_SLICE_X83Y101_BO6;
  assign CLBLL_R_X57Y106_SLICE_X86Y106_BX = 1'b0;
  assign CLBLL_R_X57Y106_SLICE_X86Y106_C1 = 1'b1;
  assign CLBLM_L_X56Y105_SLICE_X85Y105_CE = CLBLM_L_X56Y103_SLICE_X85Y103_CO6;
  assign CLBLL_R_X57Y106_SLICE_X86Y106_C2 = 1'b1;
  assign CLBLL_R_X57Y106_SLICE_X86Y106_C3 = 1'b1;
  assign CLBLL_R_X57Y106_SLICE_X86Y106_C4 = 1'b1;
  assign CLBLL_R_X57Y106_SLICE_X86Y106_C5 = 1'b1;
  assign CLBLL_R_X57Y106_SLICE_X86Y106_C6 = CLBLL_R_X57Y105_SLICE_X86Y105_BQ;
  assign CLBLM_L_X56Y105_SLICE_X85Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X56Y105_SLICE_X85Y105_C6 = CLBLL_L_X54Y105_SLICE_X82Y105_D_XOR;
  assign CLBLM_L_X56Y105_SLICE_X85Y105_D1 = CLBLM_R_X53Y103_SLICE_X81Y103_D_XOR;
  assign CLBLM_L_X56Y105_SLICE_X85Y105_D2 = CLBLM_R_X53Y106_SLICE_X81Y106_A_XOR;
  assign CLBLM_L_X56Y105_SLICE_X85Y105_D3 = CLBLM_L_X56Y105_SLICE_X85Y105_DQ;
  assign CLBLM_L_X56Y105_SLICE_X85Y105_D4 = CLBLM_R_X49Y106_SLICE_X74Y106_AQ;
  assign CLBLM_L_X56Y105_SLICE_X85Y105_D5 = CLBLL_L_X54Y101_SLICE_X83Y101_BO6;
  assign CLBLM_L_X56Y105_SLICE_X85Y105_D6 = CLBLM_L_X62Y100_SLICE_X92Y100_AO5;
  assign CLBLL_R_X57Y106_SLICE_X86Y106_CX = 1'b0;
  assign CLBLL_R_X57Y106_SLICE_X86Y106_D1 = 1'b1;
  assign CLBLM_L_X56Y105_SLICE_X85Y105_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLL_R_X57Y106_SLICE_X86Y106_D3 = 1'b1;
  assign CLBLL_R_X57Y106_SLICE_X86Y106_D4 = 1'b1;
  assign CLBLL_R_X57Y106_SLICE_X86Y106_D5 = 1'b1;
  assign CLBLL_R_X57Y106_SLICE_X86Y106_D6 = CLBLL_R_X57Y103_SLICE_X87Y103_AQ;
  assign CLBLL_R_X57Y106_SLICE_X86Y106_DX = 1'b0;
  assign CLBLM_L_X56Y105_SLICE_X84Y105_A1 = CLBLM_R_X49Y106_SLICE_X74Y106_AQ;
  assign CLBLM_L_X56Y105_SLICE_X84Y105_A2 = 1'b1;
  assign CLBLM_L_X56Y105_SLICE_X84Y105_A3 = CLBLM_L_X56Y105_SLICE_X84Y105_AQ;
  assign CLBLM_L_X56Y105_SLICE_X84Y105_A4 = CLBLM_L_X60Y99_SLICE_X90Y99_AO5;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_A1 = CLBLM_L_X56Y98_SLICE_X85Y98_DQ;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_A2 = CLBLM_L_X64Y95_SLICE_X96Y95_CO6;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_A3 = CLBLM_L_X50Y106_SLICE_X76Y106_CQ;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_A4 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_A5 = CLBLM_R_X63Y98_SLICE_X95Y98_C5Q;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_A6 = 1'b1;
  assign CLBLM_L_X56Y105_SLICE_X84Y105_A5 = CLBLL_L_X54Y101_SLICE_X83Y101_BO6;
  assign CLBLM_L_X56Y105_SLICE_X84Y105_A6 = CLBLL_L_X54Y107_SLICE_X82Y107_A_XOR;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_AX = CLBLM_R_X63Y97_SLICE_X94Y97_CO5;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_B1 = CLBLM_L_X56Y98_SLICE_X85Y98_DQ;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_B2 = 1'b1;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_B3 = CLBLM_L_X64Y95_SLICE_X96Y95_BO5;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_B4 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_B5 = CLBLM_R_X63Y99_SLICE_X95Y99_CQ;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_B6 = CLBLM_R_X49Y105_SLICE_X75Y105_CQ;
  assign CLBLM_L_X56Y105_SLICE_X84Y105_B3 = 1'b1;
  assign CLBLM_L_X56Y105_SLICE_X84Y105_B4 = CLBLM_L_X50Y106_SLICE_X76Y106_CQ;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_BX = CLBLM_R_X63Y95_SLICE_X95Y95_AO5;
  assign CLBLM_L_X56Y105_SLICE_X84Y105_B6 = CLBLM_L_X60Y99_SLICE_X90Y99_AO5;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_C1 = CLBLM_L_X64Y95_SLICE_X96Y95_BO6;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_C2 = CLBLM_R_X49Y106_SLICE_X74Y106_AQ;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_C3 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_C4 = 1'b1;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_C5 = CLBLM_L_X56Y98_SLICE_X85Y98_DQ;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_C6 = CLBLM_R_X63Y99_SLICE_X95Y99_C5Q;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_CE = CLBLM_L_X62Y99_SLICE_X93Y99_CO6;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_A4 = CLBLM_R_X49Y106_SLICE_X75Y106_DQ;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_A6 = 1'b1;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_AX = CLBLL_R_X57Y108_SLICE_X87Y108_AQ;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_B1 = 1'b1;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_B2 = CLBLL_R_X57Y108_SLICE_X87Y108_BQ;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_B3 = 1'b1;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_B4 = 1'b1;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_B5 = 1'b1;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_B6 = 1'b1;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_D3 = 1'b1;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_D4 = CLBLM_L_X50Y105_SLICE_X77Y105_AQ;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_D5 = CLBLM_L_X56Y98_SLICE_X85Y98_DQ;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_D6 = CLBLM_L_X64Y95_SLICE_X96Y95_AO6;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_BX = CLBLL_R_X57Y108_SLICE_X87Y108_BQ;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_C1 = CLBLM_R_X59Y106_SLICE_X88Y106_AQ;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_C2 = 1'b1;
  assign CLBLM_R_X63Y95_SLICE_X95Y95_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_C3 = 1'b1;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_C4 = 1'b1;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_C5 = 1'b1;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_C6 = 1'b1;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_CE = CLBLL_R_X57Y99_SLICE_X87Y99_BO6;
  assign CLBLM_R_X63Y95_SLICE_X94Y95_A3 = CLBLM_L_X62Y98_SLICE_X92Y98_DQ;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_CIN = CLBLL_R_X57Y105_SLICE_X87Y105_COUT;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_CX = CLBLM_R_X59Y106_SLICE_X88Y106_AQ;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_D1 = 1'b1;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_D2 = CLBLM_L_X60Y108_SLICE_X91Y108_AQ;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_D3 = 1'b1;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_D4 = 1'b1;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_D5 = 1'b1;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_D6 = 1'b1;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_DX = CLBLM_L_X60Y108_SLICE_X91Y108_AQ;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X63Y95_SLICE_X94Y95_A6 = 1'b1;
  assign CLBLM_R_X63Y95_SLICE_X94Y95_AI = CLBLM_R_X63Y97_SLICE_X94Y97_DQ;
  assign CLBLM_R_X63Y95_SLICE_X94Y95_AX = CLBLM_L_X62Y96_SLICE_X93Y96_CQ;
  assign CLBLM_R_X63Y95_SLICE_X94Y95_B1 = CLBLM_L_X62Y95_SLICE_X92Y95_AQ;
  assign CLBLM_R_X63Y95_SLICE_X94Y95_B2 = CLBLM_L_X62Y98_SLICE_X92Y98_CQ;
  assign CLBLM_R_X63Y95_SLICE_X94Y95_B3 = CLBLM_L_X62Y98_SLICE_X92Y98_DQ;
  assign CLBLM_R_X63Y95_SLICE_X94Y95_B4 = CLBLM_L_X62Y98_SLICE_X92Y98_AQ;
  assign CLBLM_R_X63Y95_SLICE_X94Y95_B5 = CLBLM_L_X62Y95_SLICE_X92Y95_A5Q;
  assign CLBLM_R_X63Y95_SLICE_X94Y95_B6 = 1'b1;
  assign CLBLM_R_X63Y95_SLICE_X94Y95_C2 = CLBLM_L_X62Y98_SLICE_X92Y98_CQ;
  assign CLBLM_R_X63Y95_SLICE_X94Y95_C3 = CLBLM_L_X62Y98_SLICE_X92Y98_DQ;
  assign CLBLM_R_X63Y95_SLICE_X94Y95_C4 = CLBLM_L_X62Y98_SLICE_X92Y98_AQ;
  assign CLBLM_R_X63Y95_SLICE_X94Y95_C5 = CLBLM_L_X62Y95_SLICE_X92Y95_A5Q;
  assign CLBLM_R_X63Y95_SLICE_X94Y95_C6 = 1'b1;
  assign CLBLM_R_X63Y95_SLICE_X94Y95_CE = CLBLM_L_X60Y98_SLICE_X91Y98_BQ;
  assign CLBLM_R_X63Y95_SLICE_X94Y95_BX = 1'b0;
  assign CLBLM_R_X63Y95_SLICE_X94Y95_C1 = CLBLM_L_X62Y95_SLICE_X92Y95_AQ;
  assign CLBLM_R_X63Y95_SLICE_X94Y95_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X63Y95_SLICE_X94Y95_CX = 1'b0;
  assign CLBLM_R_X63Y95_SLICE_X94Y95_D1 = CLBLM_L_X62Y95_SLICE_X93Y95_DQ;
  assign CLBLM_R_X63Y95_SLICE_X94Y95_D2 = CLBLM_L_X62Y95_SLICE_X93Y95_D5Q;
  assign CLBLM_R_X63Y95_SLICE_X94Y95_D3 = CLBLM_L_X62Y95_SLICE_X93Y95_AQ;
  assign CLBLM_R_X63Y95_SLICE_X94Y95_D4 = CLBLM_L_X62Y95_SLICE_X93Y95_BQ;
  assign CLBLM_R_X63Y95_SLICE_X94Y95_D5 = CLBLM_L_X62Y95_SLICE_X93Y95_CQ;
  assign CLBLM_R_X63Y95_SLICE_X94Y95_D6 = 1'b1;
  assign CLBLM_R_X63Y95_SLICE_X94Y95_DI = 1'b0;
  assign CLBLM_R_X63Y95_SLICE_X94Y95_DX = 1'b0;
  assign RIOI3_X105Y117_OLOGIC_X1Y117_D1 = CLBLM_R_X65Y107_SLICE_X98Y107_DQ;
  assign RIOI3_X105Y117_OLOGIC_X1Y117_T1 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X86Y107_A1 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X86Y107_A2 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X86Y107_A3 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X86Y107_A4 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X86Y107_A5 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X86Y107_A6 = CLBLL_R_X57Y108_SLICE_X87Y108_AQ;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLL_R_X57Y107_SLICE_X86Y107_AX = 1'b0;
  assign CLBLL_R_X57Y107_SLICE_X86Y107_B1 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X86Y107_B2 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X86Y107_B3 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X86Y107_B4 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X86Y107_B5 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X86Y107_B6 = CLBLL_R_X57Y108_SLICE_X87Y108_BQ;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLL_R_X57Y107_SLICE_X86Y107_BX = 1'b0;
  assign CLBLL_R_X57Y107_SLICE_X86Y107_C1 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X86Y107_C2 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X86Y107_C3 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X86Y107_C4 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X86Y107_C5 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X86Y107_C6 = CLBLM_R_X59Y106_SLICE_X88Y106_AQ;
  assign CLBLL_R_X57Y107_SLICE_X86Y107_CIN = CLBLL_R_X57Y106_SLICE_X86Y106_COUT;
  assign CLBLL_R_X57Y107_SLICE_X86Y107_CX = 1'b0;
  assign CLBLL_R_X57Y107_SLICE_X86Y107_D1 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X86Y107_D2 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X86Y107_D3 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X86Y107_D4 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X86Y107_D5 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X86Y107_D6 = CLBLM_L_X60Y108_SLICE_X91Y108_AQ;
  assign CLBLL_R_X57Y107_SLICE_X86Y107_DX = 1'b0;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_A1 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_A2 = CLBLM_R_X63Y98_SLICE_X95Y98_D5Q;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_A3 = CLBLM_L_X50Y107_SLICE_X77Y107_AQ;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_A4 = CLBLM_L_X64Y96_SLICE_X96Y96_AO6;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_A5 = CLBLM_L_X56Y98_SLICE_X85Y98_DQ;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_A6 = 1'b1;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_AX = CLBLM_R_X63Y95_SLICE_X95Y95_AO6;
  assign CLBLL_R_X57Y107_SLICE_X87Y107_A1 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X87Y107_A2 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X87Y107_A3 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X87Y107_A4 = CLBLL_R_X57Y109_SLICE_X86Y109_AQ;
  assign CLBLL_R_X57Y107_SLICE_X87Y107_A5 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X87Y107_A6 = 1'b1;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_B3 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_B4 = CLBLM_L_X64Y97_SLICE_X96Y97_B5Q;
  assign CLBLL_R_X57Y107_SLICE_X87Y107_AX = CLBLL_R_X57Y109_SLICE_X86Y109_AQ;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_B1 = CLBLM_R_X63Y96_SLICE_X94Y96_CO6;
  assign CLBLL_R_X57Y107_SLICE_X87Y107_B1 = CLBLL_R_X57Y109_SLICE_X86Y109_BQ;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_C2 = CLBLM_L_X62Y98_SLICE_X92Y98_AQ;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_C3 = CLBLM_L_X62Y96_SLICE_X93Y96_CQ;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_C4 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_C5 = CLBLM_L_X64Y96_SLICE_X97Y96_CQ;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_C6 = CLBLM_R_X63Y95_SLICE_X95Y95_CQ;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_CE = CLBLM_L_X62Y99_SLICE_X93Y99_DO6;
  assign CLBLL_R_X57Y107_SLICE_X87Y107_B2 = 1'b1;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLL_R_X57Y107_SLICE_X87Y107_B3 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X87Y107_B4 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X87Y107_B5 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X87Y107_B6 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X87Y107_BX = CLBLL_R_X57Y109_SLICE_X86Y109_BQ;
  assign CLBLL_R_X57Y107_SLICE_X87Y107_C1 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X87Y107_C2 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X87Y107_C3 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X87Y107_C4 = CLBLL_R_X57Y109_SLICE_X86Y109_CQ;
  assign CLBLL_R_X57Y107_SLICE_X87Y107_C5 = 1'b1;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_D5 = 1'b1;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_D6 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X87Y107_C6 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X87Y107_CIN = CLBLL_R_X57Y106_SLICE_X87Y106_COUT;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_D2 = 1'b1;
  assign CLBLM_R_X63Y96_SLICE_X95Y96_D3 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X87Y107_CX = 1'b0;
  assign CLBLL_R_X57Y107_SLICE_X87Y107_D1 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X87Y107_D2 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X87Y107_D3 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X87Y107_D4 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X87Y107_D5 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X87Y107_D6 = 1'b1;
  assign CLBLL_R_X57Y107_SLICE_X87Y107_DX = 1'b0;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_A1 = CLBLM_L_X62Y95_SLICE_X92Y95_AQ;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_A2 = CLBLM_L_X62Y98_SLICE_X92Y98_CQ;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_A3 = CLBLM_L_X62Y98_SLICE_X92Y98_DQ;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_A4 = CLBLM_L_X62Y98_SLICE_X92Y98_AQ;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_A5 = CLBLM_L_X62Y95_SLICE_X92Y95_A5Q;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_A6 = 1'b1;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_AI = CLBLM_L_X64Y97_SLICE_X97Y97_AQ;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_AX = CLBLM_L_X62Y96_SLICE_X92Y96_CQ;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_B1 = CLBLM_L_X62Y95_SLICE_X92Y95_AQ;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_B2 = CLBLM_L_X62Y98_SLICE_X92Y98_CQ;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_B3 = CLBLM_L_X62Y98_SLICE_X92Y98_DQ;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_B4 = CLBLM_L_X62Y98_SLICE_X92Y98_AQ;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_B5 = CLBLM_L_X62Y95_SLICE_X92Y95_A5Q;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_B6 = 1'b1;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_BI = CLBLM_L_X64Y97_SLICE_X97Y97_BQ;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_BX = CLBLM_R_X63Y94_SLICE_X94Y94_AQ;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_C1 = CLBLM_L_X62Y95_SLICE_X92Y95_AQ;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_C2 = CLBLM_L_X62Y98_SLICE_X92Y98_CQ;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_C3 = CLBLM_L_X62Y98_SLICE_X92Y98_DQ;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_C4 = CLBLM_L_X62Y98_SLICE_X92Y98_AQ;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_C5 = CLBLM_L_X62Y95_SLICE_X92Y95_A5Q;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_C6 = 1'b1;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_CE = CLBLM_L_X60Y98_SLICE_X91Y98_BQ;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_CI = CLBLM_L_X62Y96_SLICE_X93Y96_DQ;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_CX = CLBLM_R_X63Y96_SLICE_X95Y96_BQ;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_D1 = CLBLM_L_X62Y95_SLICE_X93Y95_DQ;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_D2 = CLBLM_L_X62Y95_SLICE_X93Y95_D5Q;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_D3 = CLBLM_L_X62Y95_SLICE_X93Y95_AQ;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_D4 = CLBLM_L_X62Y95_SLICE_X93Y95_BQ;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_D5 = CLBLM_L_X62Y95_SLICE_X93Y95_CQ;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_D6 = 1'b1;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_DI = 1'b0;
  assign CLBLM_R_X63Y96_SLICE_X94Y96_DX = 1'b0;
  assign CLBLL_R_X57Y108_SLICE_X86Y108_A1 = 1'b1;
  assign CLBLL_R_X57Y108_SLICE_X86Y108_A2 = 1'b1;
  assign CLBLL_R_X57Y108_SLICE_X86Y108_A3 = 1'b1;
  assign CLBLL_R_X57Y108_SLICE_X86Y108_A4 = 1'b1;
  assign CLBLL_R_X57Y108_SLICE_X86Y108_A5 = 1'b1;
  assign CLBLL_R_X57Y108_SLICE_X86Y108_A6 = CLBLL_R_X57Y109_SLICE_X86Y109_AQ;
  assign CLBLL_R_X57Y108_SLICE_X86Y108_AX = 1'b0;
  assign CLBLL_R_X57Y108_SLICE_X86Y108_B1 = 1'b1;
  assign CLBLL_R_X57Y108_SLICE_X86Y108_B2 = 1'b1;
  assign CLBLL_R_X57Y108_SLICE_X86Y108_B3 = 1'b1;
  assign CLBLL_R_X57Y108_SLICE_X86Y108_B4 = 1'b1;
  assign CLBLL_R_X57Y108_SLICE_X86Y108_B5 = 1'b1;
  assign CLBLL_R_X57Y108_SLICE_X86Y108_B6 = CLBLL_R_X57Y109_SLICE_X86Y109_BQ;
  assign CLBLL_R_X57Y108_SLICE_X86Y108_BX = 1'b0;
  assign CLBLL_R_X57Y108_SLICE_X86Y108_C1 = 1'b1;
  assign CLBLL_R_X57Y108_SLICE_X86Y108_C2 = 1'b1;
  assign CLBLL_R_X57Y108_SLICE_X86Y108_C3 = 1'b1;
  assign CLBLL_R_X57Y108_SLICE_X86Y108_C4 = 1'b1;
  assign CLBLL_R_X57Y108_SLICE_X86Y108_C5 = 1'b1;
  assign CLBLL_R_X57Y108_SLICE_X86Y108_C6 = CLBLL_R_X57Y109_SLICE_X86Y109_CQ;
  assign CLBLL_R_X57Y108_SLICE_X86Y108_CIN = CLBLL_R_X57Y107_SLICE_X86Y107_COUT;
  assign CLBLL_R_X57Y108_SLICE_X86Y108_CX = 1'b0;
  assign CLBLL_R_X57Y108_SLICE_X86Y108_D1 = 1'b1;
  assign CLBLL_R_X57Y108_SLICE_X86Y108_D2 = 1'b1;
  assign CLBLL_R_X57Y108_SLICE_X86Y108_D3 = 1'b1;
  assign CLBLL_R_X57Y108_SLICE_X86Y108_D4 = 1'b1;
  assign CLBLL_R_X57Y108_SLICE_X86Y108_D5 = 1'b1;
  assign CLBLL_R_X57Y108_SLICE_X86Y108_D6 = 1'b1;
  assign CLBLL_R_X57Y108_SLICE_X86Y108_DX = 1'b0;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_A1 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_A2 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_A3 = CLBLM_L_X62Y103_SLICE_X93Y103_AQ;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_A4 = CLBLM_R_X63Y99_SLICE_X95Y99_B5Q;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_A5 = CLBLM_R_X63Y97_SLICE_X95Y97_C5Q;
  assign CLBLL_R_X57Y108_SLICE_X87Y108_A1 = CLBLM_L_X62Y106_SLICE_X93Y106_BO5;
  assign CLBLL_R_X57Y108_SLICE_X87Y108_A2 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLL_R_X57Y108_SLICE_X87Y108_A3 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLL_R_X57Y108_SLICE_X87Y108_A4 = CLBLL_R_X57Y106_SLICE_X87Y106_A_XOR;
  assign CLBLL_R_X57Y108_SLICE_X87Y108_A5 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLL_R_X57Y108_SLICE_X87Y108_A6 = CLBLL_R_X57Y107_SLICE_X86Y107_A_XOR;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_B2 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_A6 = CLBLM_L_X62Y97_SLICE_X92Y97_BQ;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_AX = CLBLM_L_X62Y106_SLICE_X93Y106_CO6;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_B5 = CLBLM_R_X63Y96_SLICE_X95Y96_BQ;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_B1 = CLBLM_R_X63Y95_SLICE_X95Y95_DQ;
  assign CLBLL_R_X57Y108_SLICE_X87Y108_B1 = CLBLL_R_X57Y107_SLICE_X86Y107_B_XOR;
  assign CLBLL_R_X57Y108_SLICE_X87Y108_B2 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_C1 = CLBLM_L_X50Y104_SLICE_X76Y104_AQ;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_C2 = CLBLM_R_X63Y98_SLICE_X95Y98_AQ;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_C3 = CLBLM_R_X63Y98_SLICE_X95Y98_A5Q;
  assign CLBLL_R_X57Y108_SLICE_X87Y108_B3 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_C5 = CLBLM_R_X63Y99_SLICE_X94Y99_DO6;
  assign CLBLL_R_X57Y108_SLICE_X87Y108_B4 = CLBLL_R_X57Y106_SLICE_X87Y106_B_XOR;
  assign CLBLL_R_X57Y108_SLICE_X87Y108_B5 = CLBLM_L_X62Y108_SLICE_X92Y108_BO5;
  assign CLBLL_R_X57Y108_SLICE_X87Y108_B6 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLL_R_X57Y108_SLICE_X87Y108_C1 = CLBLL_R_X57Y109_SLICE_X87Y109_C_XOR;
  assign CLBLL_R_X57Y108_SLICE_X87Y108_C2 = CLBLL_R_X57Y105_SLICE_X86Y105_AQ;
  assign CLBLL_R_X57Y108_SLICE_X87Y108_C3 = CLBLL_R_X57Y106_SLICE_X86Y106_B_XOR;
  assign CLBLL_R_X57Y108_SLICE_X87Y108_C4 = CLBLM_R_X59Y103_SLICE_X88Y103_DQ;
  assign CLBLL_R_X57Y108_SLICE_X87Y108_C5 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLL_R_X57Y108_SLICE_X87Y108_C6 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLL_R_X57Y108_SLICE_X87Y108_CE = CLBLM_L_X60Y100_SLICE_X90Y100_BO6;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_D2 = CLBLM_R_X49Y106_SLICE_X74Y106_AQ;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_D3 = CLBLM_R_X63Y99_SLICE_X94Y99_DO6;
  assign CLBLL_R_X57Y108_SLICE_X87Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_D5 = CLBLM_L_X64Y97_SLICE_X96Y97_A5Q;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_D6 = 1'b1;
  assign CLBLM_R_X63Y97_SLICE_X95Y97_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLL_R_X57Y108_SLICE_X87Y108_D1 = CLBLL_R_X57Y106_SLICE_X87Y106_AQ;
  assign CLBLL_R_X57Y108_SLICE_X87Y108_D2 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLL_R_X57Y108_SLICE_X87Y108_D3 = CLBLL_R_X57Y110_SLICE_X87Y110_C_XOR;
  assign CLBLL_R_X57Y108_SLICE_X87Y108_D4 = CLBLL_R_X57Y108_SLICE_X87Y108_BQ;
  assign CLBLL_R_X57Y108_SLICE_X87Y108_D5 = CLBLL_R_X57Y107_SLICE_X86Y107_B_XOR;
  assign CLBLL_R_X57Y108_SLICE_X87Y108_D6 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLL_R_X57Y108_SLICE_X87Y108_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_A1 = CLBLM_L_X62Y97_SLICE_X92Y97_CQ;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_A2 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_A3 = CLBLM_R_X63Y98_SLICE_X94Y98_CQ;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_A4 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_A5 = CLBLM_L_X62Y97_SLICE_X93Y97_BQ;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_A6 = CLBLM_R_X63Y98_SLICE_X95Y98_CQ;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_AX = CLBLM_L_X62Y106_SLICE_X93Y106_CO6;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_B1 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_B2 = CLBLM_R_X63Y97_SLICE_X94Y97_BQ;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_B3 = CLBLM_R_X63Y95_SLICE_X95Y95_AQ;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_B4 = CLBLM_L_X62Y95_SLICE_X92Y95_A5Q;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_B5 = CLBLM_L_X64Y97_SLICE_X97Y97_AQ;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_B6 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_BX = CLBLM_R_X63Y97_SLICE_X94Y97_CO6;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_C1 = CLBLM_L_X56Y98_SLICE_X85Y98_DQ;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_C2 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_C3 = CLBLM_L_X50Y106_SLICE_X76Y106_AQ;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_C4 = CLBLM_R_X63Y98_SLICE_X95Y98_CQ;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_C5 = CLBLM_L_X64Y95_SLICE_X96Y95_CO5;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_C6 = 1'b1;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_CE = CLBLM_L_X62Y99_SLICE_X93Y99_DO6;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_CX = CLBLM_L_X62Y97_SLICE_X93Y97_CO6;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_D1 = CLBLM_L_X56Y98_SLICE_X85Y98_DQ;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_D2 = CLBLM_R_X49Y105_SLICE_X75Y105_CQ;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_D3 = 1'b1;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_D4 = CLBLM_R_X63Y95_SLICE_X94Y95_AO5;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_D5 = CLBLM_R_X63Y100_SLICE_X95Y100_AQ;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_D6 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X63Y97_SLICE_X94Y97_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign RIOI3_X105Y121_OLOGIC_X1Y122_D1 = CLBLM_L_X64Y106_SLICE_X97Y106_AQ;
  assign RIOI3_X105Y121_OLOGIC_X1Y122_T1 = 1'b1;
  assign RIOI3_X105Y121_OLOGIC_X1Y121_D1 = CLBLM_R_X65Y106_SLICE_X98Y106_AQ;
  assign RIOI3_X105Y121_OLOGIC_X1Y121_T1 = 1'b1;
  assign CLBLM_R_X65Y107_SLICE_X99Y107_B3 = 1'b1;
  assign CLBLM_R_X65Y107_SLICE_X99Y107_B4 = 1'b1;
  assign CLBLM_R_X65Y107_SLICE_X99Y107_B5 = 1'b1;
  assign CLBLL_R_X57Y109_SLICE_X86Y109_A1 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLL_R_X57Y109_SLICE_X86Y109_A2 = CLBLL_R_X57Y108_SLICE_X86Y108_A_XOR;
  assign CLBLL_R_X57Y109_SLICE_X86Y109_A3 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLL_R_X57Y109_SLICE_X86Y109_A4 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLL_R_X57Y109_SLICE_X86Y109_A5 = CLBLM_L_X62Y97_SLICE_X92Y97_BO6;
  assign CLBLL_R_X57Y109_SLICE_X86Y109_A6 = CLBLL_R_X57Y107_SLICE_X87Y107_A_XOR;
  assign CLBLL_R_X57Y109_SLICE_X86Y109_B1 = CLBLL_R_X57Y107_SLICE_X87Y107_B_XOR;
  assign CLBLL_R_X57Y109_SLICE_X86Y109_B2 = CLBLL_R_X57Y108_SLICE_X86Y108_B_XOR;
  assign CLBLL_R_X57Y109_SLICE_X86Y109_B3 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLL_R_X57Y109_SLICE_X86Y109_B4 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLL_R_X57Y109_SLICE_X86Y109_B5 = CLBLM_L_X62Y100_SLICE_X93Y100_AO6;
  assign CLBLL_R_X57Y109_SLICE_X86Y109_B6 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLL_R_X57Y109_SLICE_X86Y109_C1 = CLBLL_R_X57Y108_SLICE_X86Y108_C_XOR;
  assign CLBLL_R_X57Y109_SLICE_X86Y109_C2 = CLBLM_L_X62Y100_SLICE_X93Y100_BO6;
  assign CLBLL_R_X57Y109_SLICE_X86Y109_C3 = CLBLL_R_X57Y107_SLICE_X87Y107_C_XOR;
  assign CLBLL_R_X57Y109_SLICE_X86Y109_C4 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLL_R_X57Y109_SLICE_X86Y109_C5 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLL_R_X57Y109_SLICE_X86Y109_C6 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLL_R_X57Y109_SLICE_X86Y109_CE = CLBLM_L_X60Y100_SLICE_X90Y100_CO6;
  assign CLBLM_R_X65Y107_SLICE_X99Y107_C3 = 1'b1;
  assign CLBLL_R_X57Y109_SLICE_X86Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X65Y107_SLICE_X99Y107_C4 = 1'b1;
  assign CLBLL_R_X57Y109_SLICE_X86Y109_D1 = CLBLL_R_X57Y111_SLICE_X87Y111_C_XOR;
  assign CLBLL_R_X57Y109_SLICE_X86Y109_D2 = CLBLM_R_X59Y103_SLICE_X89Y103_BQ;
  assign CLBLL_R_X57Y109_SLICE_X86Y109_D3 = CLBLL_R_X57Y109_SLICE_X86Y109_BQ;
  assign CLBLL_R_X57Y109_SLICE_X86Y109_D4 = CLBLL_R_X57Y108_SLICE_X86Y108_B_XOR;
  assign CLBLL_R_X57Y109_SLICE_X86Y109_D5 = CLBLM_R_X59Y99_SLICE_X89Y99_BQ;
  assign CLBLL_R_X57Y109_SLICE_X86Y109_D6 = CLBLM_R_X59Y103_SLICE_X89Y103_AQ;
  assign CLBLM_R_X65Y107_SLICE_X99Y107_C5 = 1'b1;
  assign CLBLM_R_X65Y107_SLICE_X99Y107_C6 = 1'b1;
  assign CLBLL_R_X57Y109_SLICE_X86Y109_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLL_R_X57Y109_SLICE_X87Y109_A1 = 1'b1;
  assign CLBLL_R_X57Y109_SLICE_X87Y109_A2 = 1'b1;
  assign CLBLL_R_X57Y109_SLICE_X87Y109_A3 = 1'b1;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_A4 = CLBLM_R_X63Y97_SLICE_X95Y97_CQ;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_A5 = CLBLM_R_X63Y97_SLICE_X95Y97_C5Q;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_A6 = 1'b1;
  assign CLBLL_R_X57Y109_SLICE_X87Y109_A4 = 1'b1;
  assign CLBLL_R_X57Y109_SLICE_X87Y109_A5 = CLBLL_R_X57Y101_SLICE_X86Y101_AQ;
  assign CLBLL_R_X57Y109_SLICE_X87Y109_A6 = CLBLM_R_X59Y98_SLICE_X89Y98_AQ;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_A1 = CLBLM_R_X63Y99_SLICE_X94Y99_DO5;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_A2 = CLBLM_L_X64Y98_SLICE_X96Y98_AQ;
  assign CLBLL_R_X57Y109_SLICE_X87Y109_AX = CLBLL_R_X57Y101_SLICE_X86Y101_AQ;
  assign CLBLL_R_X57Y109_SLICE_X87Y109_B1 = 1'b1;
  assign CLBLL_R_X57Y109_SLICE_X87Y109_B2 = CLBLM_R_X59Y106_SLICE_X88Y106_BQ;
  assign CLBLL_R_X57Y109_SLICE_X87Y109_B3 = CLBLM_R_X59Y98_SLICE_X89Y98_A5Q;
  assign CLBLL_R_X57Y109_SLICE_X87Y109_B4 = 1'b1;
  assign CLBLL_R_X57Y109_SLICE_X87Y109_B5 = 1'b1;
  assign CLBLL_R_X57Y109_SLICE_X87Y109_B6 = 1'b1;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_B1 = CLBLM_R_X63Y99_SLICE_X94Y99_DO5;
  assign CLBLL_R_X57Y109_SLICE_X87Y109_BX = CLBLM_R_X59Y106_SLICE_X88Y106_BQ;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_C1 = CLBLM_L_X50Y106_SLICE_X76Y106_CQ;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_C2 = CLBLM_L_X50Y106_SLICE_X76Y106_AQ;
  assign CLBLL_R_X57Y109_SLICE_X87Y109_C1 = CLBLM_R_X59Y98_SLICE_X89Y98_BQ;
  assign CLBLL_R_X57Y109_SLICE_X87Y109_C2 = 1'b1;
  assign CLBLL_R_X57Y109_SLICE_X87Y109_C3 = 1'b1;
  assign CLBLL_R_X57Y109_SLICE_X87Y109_C4 = 1'b1;
  assign CLBLL_R_X57Y109_SLICE_X87Y109_C5 = 1'b1;
  assign CLBLL_R_X57Y109_SLICE_X87Y109_C6 = CLBLL_R_X57Y105_SLICE_X86Y105_AQ;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_C3 = CLBLM_L_X64Y99_SLICE_X97Y99_AQ;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_C4 = CLBLM_R_X65Y98_SLICE_X99Y98_AQ;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_C5 = CLBLM_R_X63Y99_SLICE_X94Y99_DO5;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_C6 = 1'b1;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_CE = CLBLM_L_X60Y98_SLICE_X91Y98_DQ;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLL_R_X57Y109_SLICE_X87Y109_CX = CLBLL_R_X57Y105_SLICE_X86Y105_AQ;
  assign CLBLL_R_X57Y109_SLICE_X87Y109_D1 = CLBLM_R_X59Y98_SLICE_X89Y98_B5Q;
  assign CLBLL_R_X57Y109_SLICE_X87Y109_D2 = 1'b1;
  assign CLBLL_R_X57Y109_SLICE_X87Y109_D3 = 1'b1;
  assign CLBLL_R_X57Y109_SLICE_X87Y109_D4 = 1'b1;
  assign CLBLL_R_X57Y109_SLICE_X87Y109_D5 = 1'b1;
  assign CLBLL_R_X57Y109_SLICE_X87Y109_D6 = CLBLL_R_X57Y105_SLICE_X86Y105_BQ;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_D1 = CLBLM_L_X50Y107_SLICE_X76Y107_BQ;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_D2 = CLBLM_L_X64Y99_SLICE_X96Y99_BQ;
  assign CLBLL_R_X57Y109_SLICE_X87Y109_DX = CLBLL_R_X57Y105_SLICE_X86Y105_BQ;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_D4 = CLBLM_R_X63Y99_SLICE_X94Y99_DO5;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_D5 = CLBLM_L_X50Y107_SLICE_X77Y107_AQ;
  assign CLBLM_R_X63Y98_SLICE_X95Y98_D6 = 1'b1;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_A1 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_A2 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_A3 = CLBLM_R_X63Y97_SLICE_X95Y97_CQ;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_A4 = CLBLM_R_X63Y99_SLICE_X95Y99_BQ;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_A5 = CLBLM_L_X64Y109_SLICE_X96Y109_AQ;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_A6 = CLBLM_L_X62Y97_SLICE_X92Y97_AQ;
  assign CLBLM_R_X65Y107_SLICE_X99Y107_D6 = 1'b1;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_AX = CLBLM_L_X62Y106_SLICE_X93Y106_CO6;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_B1 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_B2 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_B3 = CLBLM_R_X63Y94_SLICE_X95Y94_AQ;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_B4 = CLBLM_L_X64Y96_SLICE_X97Y96_DQ;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_B5 = CLBLM_L_X62Y95_SLICE_X92Y95_AQ;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_B6 = CLBLM_L_X62Y96_SLICE_X93Y96_DQ;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_C1 = CLBLM_L_X50Y106_SLICE_X76Y106_CQ;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_C2 = CLBLM_R_X63Y98_SLICE_X95Y98_BQ;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_C3 = CLBLM_R_X63Y98_SLICE_X95Y98_B5Q;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_C4 = CLBLM_L_X50Y106_SLICE_X76Y106_AQ;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_C5 = CLBLM_R_X63Y99_SLICE_X94Y99_DO6;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_C6 = 1'b1;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_CE = CLBLM_R_X63Y100_SLICE_X94Y100_BO6;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_A5 = 1'b1;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_D1 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_D2 = CLBLM_L_X56Y97_SLICE_X85Y97_AQ;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_D3 = CLBLM_R_X63Y94_SLICE_X94Y94_AQ;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_D4 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_D5 = 1'b1;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_D6 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X63Y98_SLICE_X94Y98_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_B5 = 1'b1;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_B6 = CLBLM_R_X59Y98_SLICE_X88Y98_AQ;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_BX = CLBLM_R_X59Y96_SLICE_X88Y96_AQ;
  assign CLBLL_L_X54Y97_SLICE_X82Y97_A1 = 1'b1;
  assign CLBLL_L_X54Y97_SLICE_X82Y97_A2 = 1'b1;
  assign CLBLL_L_X54Y97_SLICE_X82Y97_A3 = 1'b1;
  assign CLBLL_L_X54Y97_SLICE_X82Y97_A4 = 1'b1;
  assign CLBLL_L_X54Y97_SLICE_X82Y97_A5 = 1'b1;
  assign CLBLL_L_X54Y97_SLICE_X82Y97_A6 = 1'b1;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_C1 = 1'b1;
  assign CLBLL_L_X54Y97_SLICE_X82Y97_B1 = 1'b1;
  assign CLBLL_L_X54Y97_SLICE_X82Y97_B2 = 1'b1;
  assign CLBLL_L_X54Y97_SLICE_X82Y97_B3 = 1'b1;
  assign CLBLL_L_X54Y97_SLICE_X82Y97_B4 = 1'b1;
  assign CLBLL_L_X54Y97_SLICE_X82Y97_B5 = 1'b1;
  assign CLBLL_L_X54Y97_SLICE_X82Y97_B6 = 1'b1;
  assign CLBLL_L_X54Y97_SLICE_X82Y97_C1 = 1'b1;
  assign CLBLL_L_X54Y97_SLICE_X82Y97_C2 = 1'b1;
  assign CLBLL_L_X54Y97_SLICE_X82Y97_C3 = 1'b1;
  assign CLBLL_L_X54Y97_SLICE_X82Y97_C4 = 1'b1;
  assign CLBLL_L_X54Y97_SLICE_X82Y97_C5 = 1'b1;
  assign CLBLL_L_X54Y97_SLICE_X82Y97_C6 = 1'b1;
  assign CLBLM_R_X59Y97_SLICE_X89Y97_C4 = 1'b1;
  assign CLBLL_L_X54Y97_SLICE_X82Y97_D1 = 1'b1;
  assign CLBLL_L_X54Y97_SLICE_X82Y97_D2 = 1'b1;
  assign CLBLL_L_X54Y97_SLICE_X82Y97_D3 = 1'b1;
  assign CLBLL_L_X54Y97_SLICE_X82Y97_D4 = 1'b1;
  assign CLBLL_L_X54Y97_SLICE_X82Y97_D5 = 1'b1;
  assign CLBLL_L_X54Y97_SLICE_X82Y97_D6 = 1'b1;
  assign CLBLL_L_X54Y97_SLICE_X83Y97_A1 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLL_L_X54Y97_SLICE_X83Y97_A2 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLL_L_X54Y97_SLICE_X83Y97_A3 = CLBLM_R_X49Y107_SLICE_X75Y107_DQ;
  assign CLBLL_L_X54Y97_SLICE_X83Y97_A4 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLL_L_X54Y97_SLICE_X83Y97_A5 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign CLBLL_L_X54Y97_SLICE_X83Y97_A6 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLL_L_X54Y97_SLICE_X83Y97_B1 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLL_L_X54Y97_SLICE_X83Y97_B2 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLL_L_X54Y97_SLICE_X83Y97_B3 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLL_R_X57Y110_SLICE_X86Y110_A1 = 1'b1;
  assign CLBLL_R_X57Y110_SLICE_X86Y110_A2 = 1'b1;
  assign CLBLL_R_X57Y110_SLICE_X86Y110_A3 = 1'b1;
  assign CLBLL_L_X54Y97_SLICE_X83Y97_B6 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLL_R_X57Y110_SLICE_X86Y110_A4 = 1'b1;
  assign CLBLL_R_X57Y110_SLICE_X86Y110_A5 = 1'b1;
  assign CLBLL_L_X54Y97_SLICE_X83Y97_C1 = 1'b1;
  assign CLBLL_R_X57Y110_SLICE_X86Y110_A6 = 1'b1;
  assign CLBLL_L_X54Y97_SLICE_X83Y97_C3 = 1'b1;
  assign CLBLL_L_X54Y97_SLICE_X83Y97_C2 = 1'b1;
  assign CLBLL_L_X54Y97_SLICE_X83Y97_C5 = 1'b1;
  assign CLBLL_L_X54Y97_SLICE_X83Y97_C4 = 1'b1;
  assign CLBLL_R_X57Y110_SLICE_X86Y110_B1 = 1'b1;
  assign CLBLL_R_X57Y110_SLICE_X86Y110_B2 = 1'b1;
  assign CLBLL_R_X57Y110_SLICE_X86Y110_B3 = 1'b1;
  assign CLBLL_R_X57Y110_SLICE_X86Y110_B4 = 1'b1;
  assign CLBLL_R_X57Y110_SLICE_X86Y110_B5 = 1'b1;
  assign CLBLL_R_X57Y110_SLICE_X86Y110_B6 = 1'b1;
  assign CLBLL_L_X54Y97_SLICE_X83Y97_C6 = 1'b1;
  assign CLBLL_R_X57Y110_SLICE_X86Y110_C1 = 1'b1;
  assign CLBLL_R_X57Y110_SLICE_X86Y110_C3 = 1'b1;
  assign CLBLL_L_X54Y97_SLICE_X83Y97_D1 = 1'b1;
  assign CLBLL_L_X54Y97_SLICE_X83Y97_D2 = 1'b1;
  assign CLBLL_L_X54Y97_SLICE_X83Y97_D3 = 1'b1;
  assign CLBLL_L_X54Y97_SLICE_X83Y97_D4 = 1'b1;
  assign CLBLL_L_X54Y97_SLICE_X83Y97_D5 = 1'b1;
  assign CLBLL_L_X54Y97_SLICE_X83Y97_D6 = 1'b1;
  assign CLBLL_R_X57Y110_SLICE_X86Y110_C5 = 1'b1;
  assign CLBLL_R_X57Y110_SLICE_X86Y110_C6 = 1'b1;
  assign CLBLL_R_X57Y110_SLICE_X86Y110_D1 = 1'b1;
  assign CLBLL_R_X57Y110_SLICE_X86Y110_D2 = 1'b1;
  assign CLBLL_R_X57Y110_SLICE_X86Y110_D4 = 1'b1;
  assign CLBLL_R_X57Y110_SLICE_X86Y110_D5 = 1'b1;
  assign CLBLL_R_X57Y110_SLICE_X86Y110_D6 = 1'b1;
  assign CLBLL_R_X57Y110_SLICE_X86Y110_D3 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_T1 = 1'b1;
  assign CLBLL_R_X57Y110_SLICE_X87Y110_A1 = 1'b1;
  assign CLBLL_R_X57Y110_SLICE_X87Y110_A2 = 1'b1;
  assign CLBLL_R_X57Y110_SLICE_X87Y110_A3 = CLBLM_R_X59Y98_SLICE_X89Y98_CQ;
  assign CLBLL_R_X57Y110_SLICE_X87Y110_A4 = 1'b1;
  assign CLBLL_R_X57Y110_SLICE_X87Y110_A5 = CLBLL_R_X57Y103_SLICE_X87Y103_AQ;
  assign CLBLL_R_X57Y110_SLICE_X87Y110_A6 = 1'b1;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_A1 = CLBLM_R_X65Y105_SLICE_X98Y105_AQ;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_A2 = CLBLM_R_X63Y99_SLICE_X94Y99_DO5;
  assign CLBLL_R_X57Y110_SLICE_X87Y110_AX = CLBLL_R_X57Y103_SLICE_X87Y103_AQ;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_A3 = CLBLM_R_X63Y99_SLICE_X94Y99_C5Q;
  assign CLBLL_R_X57Y110_SLICE_X87Y110_B1 = 1'b1;
  assign CLBLL_R_X57Y110_SLICE_X87Y110_B2 = CLBLM_R_X59Y98_SLICE_X89Y98_C5Q;
  assign CLBLL_R_X57Y110_SLICE_X87Y110_B3 = CLBLL_R_X57Y108_SLICE_X87Y108_AQ;
  assign CLBLL_R_X57Y110_SLICE_X87Y110_B4 = 1'b1;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_B1 = CLBLM_L_X50Y105_SLICE_X77Y105_AQ;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_B2 = CLBLM_R_X63Y99_SLICE_X94Y99_DO5;
  assign CLBLL_R_X57Y110_SLICE_X87Y110_B5 = 1'b1;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_B4 = 1'b1;
  assign CLBLL_R_X57Y110_SLICE_X87Y110_B6 = 1'b1;
  assign CLBLL_R_X57Y110_SLICE_X87Y110_BX = CLBLL_R_X57Y108_SLICE_X87Y108_AQ;
  assign CLBLL_R_X57Y110_SLICE_X87Y110_C1 = CLBLL_R_X57Y108_SLICE_X87Y108_BQ;
  assign CLBLL_R_X57Y110_SLICE_X87Y110_C2 = CLBLM_R_X59Y96_SLICE_X89Y96_AQ;
  assign CLBLL_R_X57Y110_SLICE_X87Y110_C3 = 1'b1;
  assign CLBLL_R_X57Y110_SLICE_X87Y110_C4 = 1'b1;
  assign CLBLL_R_X57Y110_SLICE_X87Y110_C5 = 1'b1;
  assign CLBLL_R_X57Y110_SLICE_X87Y110_C6 = 1'b1;
  assign CLBLL_R_X57Y110_SLICE_X87Y110_CIN = CLBLL_R_X57Y109_SLICE_X87Y109_COUT;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_C4 = CLBLM_R_X49Y105_SLICE_X75Y105_CQ;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_C5 = CLBLM_R_X65Y99_SLICE_X99Y99_AQ;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_C6 = 1'b1;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_CE = CLBLM_L_X60Y98_SLICE_X91Y98_DQ;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_C1 = CLBLM_R_X65Y99_SLICE_X98Y99_AQ;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_C2 = CLBLM_R_X49Y106_SLICE_X74Y106_AQ;
  assign CLBLL_R_X57Y110_SLICE_X87Y110_CX = CLBLL_R_X57Y108_SLICE_X87Y108_BQ;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_C3 = CLBLM_R_X63Y99_SLICE_X94Y99_DO5;
  assign CLBLL_R_X57Y110_SLICE_X87Y110_D1 = CLBLM_R_X59Y106_SLICE_X88Y106_AQ;
  assign CLBLL_R_X57Y110_SLICE_X87Y110_D2 = CLBLM_R_X59Y96_SLICE_X89Y96_A5Q;
  assign CLBLL_R_X57Y110_SLICE_X87Y110_D3 = 1'b1;
  assign CLBLL_R_X57Y110_SLICE_X87Y110_D4 = 1'b1;
  assign CLBLL_R_X57Y110_SLICE_X87Y110_D5 = 1'b1;
  assign CLBLL_R_X57Y110_SLICE_X87Y110_D6 = 1'b1;
  assign CLBLL_R_X57Y110_SLICE_X87Y110_DX = CLBLM_R_X59Y106_SLICE_X88Y106_AQ;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_D1 = 1'b1;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_D2 = 1'b1;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_D3 = 1'b1;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_D4 = 1'b1;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_D5 = 1'b1;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_D6 = 1'b1;
  assign CLBLM_R_X63Y99_SLICE_X95Y99_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_A1 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_A2 = CLBLM_R_X63Y105_SLICE_X94Y105_AQ;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_A3 = CLBLM_L_X62Y100_SLICE_X93Y100_AQ;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_A4 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_A5 = CLBLM_R_X63Y97_SLICE_X95Y97_DQ;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_A6 = CLBLM_R_X63Y99_SLICE_X95Y99_CQ;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_AX = CLBLM_L_X62Y106_SLICE_X93Y106_CO6;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_B1 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_B2 = CLBLM_R_X63Y95_SLICE_X95Y95_BQ;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_B3 = CLBLM_L_X62Y98_SLICE_X92Y98_DQ;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_B4 = CLBLM_L_X64Y96_SLICE_X97Y96_BQ;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_B5 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_B6 = CLBLM_R_X63Y97_SLICE_X94Y97_DQ;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_C1 = CLBLM_R_X63Y99_SLICE_X95Y99_AQ;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_C2 = CLBLM_R_X63Y99_SLICE_X95Y99_A5Q;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_C3 = CLBLM_L_X50Y107_SLICE_X76Y107_BQ;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_C4 = CLBLM_L_X50Y107_SLICE_X77Y107_AQ;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_C5 = CLBLM_R_X63Y99_SLICE_X94Y99_DO6;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_C6 = 1'b1;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_CE = CLBLM_R_X63Y100_SLICE_X94Y100_BO6;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_D1 = CLBLM_L_X62Y104_SLICE_X93Y104_AQ;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_D2 = CLBLM_L_X60Y98_SLICE_X90Y98_BQ;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_D3 = CLBLM_R_X59Y102_SLICE_X89Y102_AQ;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_D4 = CLBLM_L_X62Y102_SLICE_X93Y102_AO5;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_D5 = CLBLM_R_X59Y102_SLICE_X88Y102_AQ;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_D6 = 1'b1;
  assign CLBLM_R_X63Y99_SLICE_X94Y99_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLL_L_X54Y98_SLICE_X82Y98_A1 = CLBLL_L_X54Y98_SLICE_X82Y98_BO6;
  assign CLBLL_L_X54Y98_SLICE_X82Y98_A2 = CLBLM_R_X53Y100_SLICE_X81Y100_DO6;
  assign CLBLL_L_X54Y98_SLICE_X82Y98_A3 = CLBLM_R_X53Y99_SLICE_X80Y99_AO5;
  assign CLBLL_L_X54Y98_SLICE_X82Y98_A4 = CLBLM_R_X53Y98_SLICE_X81Y98_AO6;
  assign CLBLL_L_X54Y98_SLICE_X82Y98_A5 = CLBLM_R_X49Y107_SLICE_X75Y107_DQ;
  assign CLBLL_L_X54Y98_SLICE_X82Y98_A6 = CLBLM_R_X53Y100_SLICE_X81Y100_AO5;
  assign CLBLL_L_X54Y98_SLICE_X82Y98_B1 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLL_L_X54Y98_SLICE_X82Y98_B2 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign CLBLL_L_X54Y98_SLICE_X82Y98_B3 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLL_L_X54Y98_SLICE_X82Y98_B4 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLL_L_X54Y98_SLICE_X82Y98_B5 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLL_L_X54Y98_SLICE_X82Y98_B6 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLL_L_X54Y98_SLICE_X82Y98_C1 = CLBLM_R_X49Y107_SLICE_X75Y107_DQ;
  assign CLBLL_L_X54Y98_SLICE_X82Y98_C2 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLL_L_X54Y98_SLICE_X82Y98_C3 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLL_L_X54Y98_SLICE_X82Y98_C4 = CLBLM_R_X53Y100_SLICE_X81Y100_AO5;
  assign CLBLL_L_X54Y98_SLICE_X82Y98_C5 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLL_L_X54Y98_SLICE_X82Y98_C6 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign CLBLL_L_X54Y98_SLICE_X82Y98_D1 = CLBLM_R_X49Y107_SLICE_X75Y107_DQ;
  assign CLBLL_L_X54Y98_SLICE_X82Y98_D2 = CLBLL_L_X54Y99_SLICE_X83Y99_BO5;
  assign CLBLL_L_X54Y98_SLICE_X82Y98_D3 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLL_L_X54Y98_SLICE_X82Y98_D4 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLL_L_X54Y98_SLICE_X82Y98_D5 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLL_L_X54Y98_SLICE_X82Y98_D6 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign RIOI3_X105Y123_OLOGIC_X1Y124_D1 = CLBLM_R_X65Y106_SLICE_X98Y106_BQ;
  assign CLBLL_L_X54Y98_SLICE_X83Y98_A1 = CLBLM_R_X53Y99_SLICE_X81Y99_AO6;
  assign CLBLL_L_X54Y98_SLICE_X83Y98_A2 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign CLBLL_L_X54Y98_SLICE_X83Y98_A3 = CLBLL_L_X54Y97_SLICE_X83Y97_AO6;
  assign CLBLL_L_X54Y98_SLICE_X83Y98_A4 = CLBLL_L_X54Y98_SLICE_X82Y98_CO6;
  assign CLBLL_L_X54Y98_SLICE_X83Y98_A5 = CLBLL_L_X54Y98_SLICE_X83Y98_CO5;
  assign CLBLL_L_X54Y98_SLICE_X83Y98_A6 = CLBLL_L_X54Y99_SLICE_X83Y99_BO5;
  assign RIOI3_X105Y123_OLOGIC_X1Y124_T1 = 1'b1;
  assign CLBLL_L_X54Y98_SLICE_X83Y98_B1 = CLBLM_R_X53Y99_SLICE_X80Y99_AO5;
  assign CLBLL_L_X54Y98_SLICE_X83Y98_B2 = CLBLM_R_X53Y99_SLICE_X81Y99_CO6;
  assign CLBLL_L_X54Y98_SLICE_X83Y98_B3 = CLBLL_L_X54Y97_SLICE_X83Y97_BO6;
  assign CLBLL_L_X54Y98_SLICE_X83Y98_B4 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLL_L_X54Y98_SLICE_X83Y98_B5 = CLBLM_L_X56Y98_SLICE_X84Y98_AO6;
  assign CLBLL_R_X57Y111_SLICE_X86Y111_A4 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X86Y111_A5 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X86Y111_A6 = 1'b1;
  assign CLBLL_L_X54Y98_SLICE_X83Y98_B6 = CLBLL_L_X54Y98_SLICE_X83Y98_CO6;
  assign CLBLL_R_X57Y111_SLICE_X86Y111_A1 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X86Y111_A2 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X86Y111_B1 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X86Y111_B2 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X86Y111_B4 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X86Y111_B5 = 1'b1;
  assign CLBLL_L_X54Y98_SLICE_X83Y98_C1 = 1'b1;
  assign CLBLL_L_X54Y98_SLICE_X83Y98_C2 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLL_L_X54Y98_SLICE_X83Y98_C3 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLL_L_X54Y98_SLICE_X83Y98_C4 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X86Y111_B6 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X86Y111_C1 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X86Y111_C2 = 1'b1;
  assign CLBLL_L_X54Y98_SLICE_X83Y98_C6 = 1'b1;
  assign CLBLL_L_X54Y98_SLICE_X83Y98_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X0Y20_O;
  assign CLBLL_R_X57Y111_SLICE_X86Y111_C3 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X86Y111_C4 = 1'b1;
  assign CLBLL_L_X54Y98_SLICE_X83Y98_D1 = CLBLM_R_X49Y107_SLICE_X75Y107_DQ;
  assign CLBLL_L_X54Y98_SLICE_X83Y98_D2 = CLBLL_L_X54Y99_SLICE_X83Y99_BO5;
  assign CLBLL_L_X54Y98_SLICE_X83Y98_D3 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLL_L_X54Y98_SLICE_X83Y98_D4 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLL_L_X54Y98_SLICE_X83Y98_D5 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign CLBLL_L_X54Y98_SLICE_X83Y98_D6 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLL_L_X54Y98_SLICE_X83Y98_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLL_R_X57Y111_SLICE_X86Y111_D1 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X86Y111_D2 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X86Y111_D3 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X86Y111_D4 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X86Y111_D5 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X86Y111_D6 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X87Y111_A1 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X87Y111_A2 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X87Y111_A3 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X87Y111_A4 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X87Y111_A5 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X87Y111_A6 = CLBLM_L_X60Y108_SLICE_X91Y108_AQ;
  assign CLBLL_R_X57Y111_SLICE_X87Y111_AX = 1'b0;
  assign CLBLL_R_X57Y111_SLICE_X87Y111_B1 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X87Y111_B2 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X87Y111_B3 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X87Y111_B4 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X87Y111_B5 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X87Y111_B6 = CLBLL_R_X57Y109_SLICE_X86Y109_AQ;
  assign CLBLM_R_X63Y100_SLICE_X95Y100_A1 = CLBLM_L_X62Y100_SLICE_X93Y100_BQ;
  assign CLBLM_R_X63Y100_SLICE_X95Y100_A2 = CLBLM_L_X62Y100_SLICE_X93Y100_AQ;
  assign CLBLL_R_X57Y111_SLICE_X87Y111_BX = 1'b0;
  assign CLBLM_R_X63Y100_SLICE_X95Y100_A3 = CLBLM_R_X63Y99_SLICE_X94Y99_DO5;
  assign CLBLL_R_X57Y111_SLICE_X87Y111_C1 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X87Y111_C2 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X87Y111_C3 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X87Y111_C4 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X87Y111_C5 = 1'b1;
  assign CLBLM_R_X63Y100_SLICE_X95Y100_B6 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLL_R_X57Y111_SLICE_X87Y111_C6 = CLBLL_R_X57Y109_SLICE_X86Y109_BQ;
  assign CLBLL_R_X57Y111_SLICE_X87Y111_CIN = CLBLL_R_X57Y110_SLICE_X87Y110_COUT;
  assign CLBLM_R_X63Y100_SLICE_X95Y100_B1 = 1'b1;
  assign CLBLM_R_X63Y100_SLICE_X95Y100_C1 = 1'b1;
  assign CLBLM_R_X63Y100_SLICE_X95Y100_C2 = CLBLM_R_X63Y97_SLICE_X95Y97_D5Q;
  assign CLBLM_R_X63Y100_SLICE_X95Y100_C3 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_R_X63Y100_SLICE_X95Y100_C4 = CLBLM_L_X62Y100_SLICE_X93Y100_BQ;
  assign CLBLM_R_X63Y100_SLICE_X95Y100_C5 = 1'b1;
  assign CLBLM_R_X63Y100_SLICE_X95Y100_C6 = 1'b1;
  assign CLBLM_R_X63Y100_SLICE_X95Y100_CE = CLBLM_L_X60Y98_SLICE_X91Y98_DQ;
  assign CLBLL_R_X57Y111_SLICE_X87Y111_CX = 1'b0;
  assign CLBLM_R_X63Y100_SLICE_X95Y100_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X57Y111_SLICE_X87Y111_D1 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X87Y111_D2 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X87Y111_D3 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X87Y111_D4 = 1'b1;
  assign CLBLL_R_X57Y111_SLICE_X87Y111_DX = 1'b0;
  assign CLBLM_R_X63Y100_SLICE_X95Y100_D1 = 1'b1;
  assign CLBLM_R_X63Y100_SLICE_X95Y100_D2 = 1'b1;
  assign CLBLM_R_X63Y100_SLICE_X95Y100_D3 = 1'b1;
  assign CLBLM_R_X63Y100_SLICE_X95Y100_D4 = 1'b1;
  assign CLBLM_R_X63Y100_SLICE_X95Y100_D5 = 1'b1;
  assign CLBLM_R_X63Y100_SLICE_X95Y100_D6 = 1'b1;
  assign CLBLM_R_X63Y100_SLICE_X95Y100_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X63Y100_SLICE_X94Y100_A1 = CLBLM_R_X63Y100_SLICE_X94Y100_DO6;
  assign CLBLM_R_X63Y100_SLICE_X94Y100_A2 = CLBLM_L_X60Y100_SLICE_X91Y100_CO6;
  assign CLBLM_R_X63Y100_SLICE_X94Y100_A3 = CLBLM_R_X63Y100_SLICE_X94Y100_AQ;
  assign CLBLM_R_X63Y100_SLICE_X94Y100_A4 = CLBLM_L_X50Y104_SLICE_X76Y104_AQ;
  assign CLBLM_R_X63Y100_SLICE_X94Y100_A5 = CLBLM_L_X60Y99_SLICE_X91Y99_AO6;
  assign CLBLM_R_X63Y100_SLICE_X94Y100_A6 = CLBLM_L_X56Y103_SLICE_X85Y103_CO6;
  assign CLBLM_R_X63Y100_SLICE_X94Y100_B1 = CLBLM_L_X62Y102_SLICE_X93Y102_AO5;
  assign CLBLM_R_X63Y100_SLICE_X94Y100_B2 = CLBLM_R_X59Y102_SLICE_X89Y102_AQ;
  assign CLBLM_R_X63Y100_SLICE_X94Y100_B3 = CLBLM_R_X59Y102_SLICE_X88Y102_AQ;
  assign CLBLM_R_X63Y100_SLICE_X94Y100_B4 = CLBLM_L_X56Y103_SLICE_X85Y103_CO6;
  assign CLBLM_R_X63Y100_SLICE_X94Y100_B5 = CLBLM_L_X60Y98_SLICE_X90Y98_BQ;
  assign CLBLM_R_X63Y100_SLICE_X94Y100_B6 = CLBLM_L_X62Y104_SLICE_X93Y104_AQ;
  assign CLBLM_R_X63Y100_SLICE_X94Y100_C1 = CLBLM_L_X60Y99_SLICE_X91Y99_AO6;
  assign CLBLM_R_X63Y100_SLICE_X94Y100_C2 = CLBLM_L_X62Y99_SLICE_X92Y99_AO6;
  assign CLBLM_R_X63Y100_SLICE_X94Y100_C3 = CLBLM_R_X59Y102_SLICE_X89Y102_AQ;
  assign CLBLM_R_X63Y100_SLICE_X94Y100_C4 = CLBLM_L_X62Y104_SLICE_X93Y104_AQ;
  assign CLBLM_R_X63Y100_SLICE_X94Y100_C5 = CLBLM_L_X60Y99_SLICE_X91Y99_BO6;
  assign CLBLM_R_X63Y100_SLICE_X94Y100_C6 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X63Y100_SLICE_X94Y100_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X63Y100_SLICE_X94Y100_D1 = 1'b1;
  assign CLBLM_R_X63Y100_SLICE_X94Y100_D2 = 1'b1;
  assign CLBLM_R_X63Y100_SLICE_X94Y100_D3 = 1'b1;
  assign CLBLM_R_X63Y100_SLICE_X94Y100_D4 = CLBLM_L_X62Y104_SLICE_X93Y104_AQ;
  assign CLBLM_R_X63Y100_SLICE_X94Y100_D5 = CLBLM_R_X59Y102_SLICE_X89Y102_AQ;
  assign CLBLM_R_X63Y100_SLICE_X94Y100_D6 = 1'b1;
  assign CLBLM_R_X63Y100_SLICE_X94Y100_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLL_L_X54Y99_SLICE_X82Y99_A1 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLL_L_X54Y99_SLICE_X82Y99_A2 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLL_L_X54Y99_SLICE_X82Y99_A3 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLL_L_X54Y99_SLICE_X82Y99_A4 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign CLBLL_L_X54Y99_SLICE_X82Y99_A5 = 1'b1;
  assign CLBLL_L_X54Y99_SLICE_X82Y99_A6 = 1'b1;
  assign CLBLL_L_X54Y99_SLICE_X82Y99_AX = CLBLL_L_X54Y99_SLICE_X82Y99_BO5;
  assign CLBLL_L_X54Y99_SLICE_X82Y99_B1 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLL_L_X54Y99_SLICE_X82Y99_B2 = CLBLM_R_X53Y99_SLICE_X81Y99_CO6;
  assign CLBLL_L_X54Y99_SLICE_X82Y99_B3 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLL_L_X54Y99_SLICE_X82Y99_B4 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign CLBLL_L_X54Y99_SLICE_X82Y99_B5 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLL_L_X54Y99_SLICE_X82Y99_B6 = 1'b1;
  assign CLBLL_L_X54Y99_SLICE_X82Y99_C1 = CLBLM_L_X56Y97_SLICE_X84Y97_CO5;
  assign CLBLL_L_X54Y99_SLICE_X82Y99_C2 = CLBLM_R_X53Y99_SLICE_X80Y99_DO6;
  assign CLBLL_L_X54Y99_SLICE_X82Y99_C3 = CLBLL_L_X54Y99_SLICE_X82Y99_AO5;
  assign CLBLL_L_X54Y99_SLICE_X82Y99_C4 = CLBLL_L_X54Y98_SLICE_X82Y98_DO6;
  assign CLBLL_L_X54Y99_SLICE_X82Y99_C5 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLL_L_X54Y99_SLICE_X82Y99_C6 = CLBLM_R_X53Y98_SLICE_X81Y98_AO6;
  assign CLBLL_L_X54Y99_SLICE_X82Y99_CE = CLBLM_L_X60Y98_SLICE_X91Y98_DQ;
  assign CLBLL_L_X54Y99_SLICE_X82Y99_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X0Y20_O;
  assign CLBLL_L_X54Y99_SLICE_X82Y99_D1 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLL_L_X54Y99_SLICE_X82Y99_D2 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLL_L_X54Y99_SLICE_X82Y99_D3 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLL_L_X54Y99_SLICE_X82Y99_D4 = CLBLM_R_X53Y100_SLICE_X81Y100_AO5;
  assign CLBLL_L_X54Y99_SLICE_X82Y99_D5 = CLBLM_R_X53Y99_SLICE_X81Y99_AO6;
  assign CLBLL_L_X54Y99_SLICE_X82Y99_D6 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign CLBLL_L_X54Y99_SLICE_X82Y99_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLL_L_X54Y99_SLICE_X83Y99_A1 = CLBLL_L_X54Y99_SLICE_X83Y99_DO6;
  assign CLBLL_L_X54Y99_SLICE_X83Y99_A2 = CLBLM_R_X53Y99_SLICE_X80Y99_AO5;
  assign CLBLL_L_X54Y99_SLICE_X83Y99_A3 = CLBLL_L_X52Y99_SLICE_X79Y99_AO6;
  assign CLBLL_L_X54Y99_SLICE_X83Y99_A4 = CLBLL_L_X54Y99_SLICE_X83Y99_BO6;
  assign CLBLL_L_X54Y99_SLICE_X83Y99_A5 = CLBLM_R_X49Y107_SLICE_X75Y107_DQ;
  assign CLBLL_L_X54Y99_SLICE_X83Y99_A6 = CLBLL_L_X54Y100_SLICE_X83Y100_AO5;
  assign CLBLL_L_X54Y99_SLICE_X83Y99_AX = CLBLL_L_X54Y99_SLICE_X83Y99_AQ;
  assign CLBLL_L_X54Y99_SLICE_X83Y99_B1 = 1'b1;
  assign CLBLL_L_X54Y99_SLICE_X83Y99_B2 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLL_L_X54Y99_SLICE_X83Y99_B3 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLL_L_X54Y99_SLICE_X83Y99_B4 = 1'b1;
  assign CLBLL_L_X54Y99_SLICE_X83Y99_B5 = 1'b1;
  assign CLBLL_L_X54Y99_SLICE_X83Y99_B6 = 1'b1;
  assign CLBLL_L_X54Y99_SLICE_X83Y99_C1 = CLBLL_L_X54Y98_SLICE_X83Y98_CO5;
  assign CLBLL_L_X54Y99_SLICE_X83Y99_C2 = CLBLM_R_X49Y108_SLICE_X75Y108_DQ;
  assign CLBLL_L_X54Y99_SLICE_X83Y99_C3 = CLBLM_R_X49Y107_SLICE_X75Y107_DQ;
  assign CLBLL_L_X54Y99_SLICE_X83Y99_C4 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign CLBLL_L_X54Y99_SLICE_X83Y99_C5 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLL_L_X54Y99_SLICE_X83Y99_C6 = CLBLL_L_X54Y99_SLICE_X83Y99_BO6;
  assign CLBLL_L_X54Y99_SLICE_X83Y99_CE = CLBLM_L_X60Y98_SLICE_X91Y98_DQ;
  assign CLBLL_L_X54Y99_SLICE_X83Y99_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X0Y20_O;
  assign CLBLL_L_X54Y109_SLICE_X82Y109_AX = CLBLL_L_X54Y103_SLICE_X82Y103_AQ;
  assign CLBLL_L_X54Y99_SLICE_X83Y99_D1 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLL_L_X54Y99_SLICE_X83Y99_D2 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLL_L_X54Y99_SLICE_X83Y99_D3 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLL_L_X54Y99_SLICE_X83Y99_D4 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLL_L_X54Y99_SLICE_X83Y99_D5 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLL_L_X54Y99_SLICE_X83Y99_D6 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign CLBLL_L_X54Y99_SLICE_X83Y99_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X56Y111_SLICE_X85Y111_A1 = 1'b1;
  assign CLBLM_L_X56Y111_SLICE_X85Y111_A2 = 1'b1;
  assign CLBLM_L_X56Y111_SLICE_X85Y111_A3 = 1'b1;
  assign CLBLM_L_X56Y111_SLICE_X85Y111_A4 = 1'b1;
  assign CLBLM_L_X56Y111_SLICE_X85Y111_A5 = 1'b1;
  assign CLBLM_L_X56Y111_SLICE_X85Y111_A6 = 1'b1;
  assign CLBLM_L_X56Y111_SLICE_X85Y111_B1 = 1'b1;
  assign CLBLM_L_X56Y111_SLICE_X85Y111_B2 = 1'b1;
  assign CLBLM_L_X56Y111_SLICE_X85Y111_B3 = 1'b1;
  assign CLBLM_L_X56Y111_SLICE_X85Y111_B4 = 1'b1;
  assign CLBLM_L_X56Y111_SLICE_X85Y111_B5 = 1'b1;
  assign CLBLM_L_X56Y111_SLICE_X85Y111_B6 = 1'b1;
  assign CLBLM_L_X56Y111_SLICE_X85Y111_C1 = 1'b1;
  assign CLBLM_L_X56Y111_SLICE_X85Y111_C2 = 1'b1;
  assign CLBLM_L_X56Y111_SLICE_X85Y111_C3 = 1'b1;
  assign CLBLM_L_X56Y111_SLICE_X85Y111_C4 = 1'b1;
  assign CLBLM_L_X56Y111_SLICE_X85Y111_C5 = 1'b1;
  assign CLBLM_L_X56Y111_SLICE_X85Y111_C6 = 1'b1;
  assign CLBLM_L_X56Y111_SLICE_X85Y111_D1 = 1'b1;
  assign CLBLM_L_X56Y111_SLICE_X85Y111_D2 = 1'b1;
  assign CLBLM_L_X56Y111_SLICE_X85Y111_D3 = 1'b1;
  assign CLBLM_L_X56Y111_SLICE_X85Y111_D4 = 1'b1;
  assign CLBLM_L_X56Y111_SLICE_X85Y111_D5 = 1'b1;
  assign CLBLM_L_X56Y111_SLICE_X85Y111_D6 = 1'b1;
  assign CLBLM_L_X56Y111_SLICE_X84Y111_A1 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_L_X56Y111_SLICE_X84Y111_A2 = CLBLL_R_X57Y102_SLICE_X86Y102_BQ;
  assign CLBLM_L_X56Y111_SLICE_X84Y111_A3 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_L_X56Y111_SLICE_X84Y111_A4 = 1'b1;
  assign CLBLM_L_X56Y111_SLICE_X84Y111_A5 = CLBLL_R_X57Y102_SLICE_X86Y102_AQ;
  assign CLBLM_L_X56Y111_SLICE_X84Y111_A6 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_A1 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_A2 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_A3 = CLBLM_L_X64Y98_SLICE_X97Y98_AQ;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_A4 = CLBLL_R_X57Y103_SLICE_X86Y103_AQ;
  assign CLBLM_L_X56Y111_SLICE_X84Y111_B1 = 1'b1;
  assign CLBLM_L_X56Y111_SLICE_X84Y111_B2 = 1'b1;
  assign CLBLM_L_X56Y111_SLICE_X84Y111_B3 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_A5 = CLBLM_L_X64Y107_SLICE_X97Y107_BQ;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_A6 = CLBLL_R_X57Y103_SLICE_X86Y103_A5Q;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_B1 = CLBLM_L_X64Y109_SLICE_X96Y109_A5Q;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_B2 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_B3 = CLBLM_R_X63Y99_SLICE_X95Y99_C5Q;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_B4 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_B5 = CLBLM_R_X63Y100_SLICE_X95Y100_CO6;
  assign CLBLM_L_X56Y111_SLICE_X84Y111_C1 = 1'b1;
  assign CLBLM_L_X56Y111_SLICE_X84Y111_C2 = 1'b1;
  assign CLBLM_L_X56Y111_SLICE_X84Y111_C3 = 1'b1;
  assign CLBLM_L_X56Y111_SLICE_X84Y111_C4 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_B6 = CLBLM_L_X62Y106_SLICE_X93Y106_CO6;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_C1 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_C2 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_C3 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_C4 = CLBLM_R_X49Y104_SLICE_X75Y104_BQ;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_C5 = CLBLM_L_X64Y102_SLICE_X97Y102_C_XOR;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_C6 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_CE = CLBLM_L_X62Y105_SLICE_X93Y105_DO6;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X56Y111_SLICE_X84Y111_C6 = 1'b1;
  assign CLBLM_L_X56Y111_SLICE_X84Y111_CE = CLBLM_R_X49Y111_SLICE_X75Y111_BO6;
  assign CLBLM_L_X56Y111_SLICE_X84Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_D1 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_D2 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_D3 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_D4 = CLBLM_L_X64Y102_SLICE_X97Y102_A_XOR;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_D5 = CLBLM_R_X49Y104_SLICE_X74Y104_AQ;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_D6 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_L_X56Y111_SLICE_X84Y111_D2 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X95Y101_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_L_X56Y111_SLICE_X84Y111_D5 = 1'b1;
  assign CLBLM_L_X56Y111_SLICE_X84Y111_D6 = 1'b1;
  assign CLBLM_L_X56Y111_SLICE_X84Y111_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_A1 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_A2 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_A3 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_A4 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_A5 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_A6 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_B1 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_B2 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_B3 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_B4 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_B5 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_B6 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_C1 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_C2 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_C3 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_C4 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_C5 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_C6 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_D1 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_D2 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_D3 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_D4 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_D5 = 1'b1;
  assign CLBLM_R_X63Y101_SLICE_X94Y101_D6 = 1'b1;
  assign CLBLL_L_X54Y100_SLICE_X82Y100_A1 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLL_L_X54Y100_SLICE_X82Y100_A2 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign CLBLL_L_X54Y100_SLICE_X82Y100_A3 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLL_L_X54Y100_SLICE_X82Y100_A4 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLL_L_X54Y100_SLICE_X82Y100_A5 = 1'b1;
  assign CLBLL_L_X54Y100_SLICE_X82Y100_A6 = 1'b1;
  assign CLBLL_L_X54Y100_SLICE_X82Y100_B1 = CLBLL_L_X54Y100_SLICE_X82Y100_DO6;
  assign CLBLL_L_X54Y100_SLICE_X82Y100_B2 = CLBLL_L_X54Y100_SLICE_X83Y100_BO6;
  assign CLBLL_L_X54Y100_SLICE_X82Y100_B3 = CLBLL_L_X54Y100_SLICE_X83Y100_AO6;
  assign CLBLL_L_X54Y100_SLICE_X82Y100_B4 = CLBLM_L_X56Y99_SLICE_X84Y99_CO6;
  assign CLBLL_L_X54Y100_SLICE_X82Y100_B5 = 1'b1;
  assign CLBLL_L_X54Y100_SLICE_X82Y100_B6 = CLBLL_L_X54Y100_SLICE_X82Y100_CO6;
  assign CLBLL_L_X54Y100_SLICE_X82Y100_C1 = CLBLL_L_X54Y100_SLICE_X82Y100_AO6;
  assign CLBLL_L_X54Y100_SLICE_X82Y100_C2 = CLBLM_R_X49Y107_SLICE_X75Y107_DQ;
  assign CLBLL_L_X54Y100_SLICE_X82Y100_C3 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLL_L_X54Y100_SLICE_X82Y100_C4 = CLBLM_R_X53Y99_SLICE_X80Y99_AO5;
  assign CLBLL_L_X54Y100_SLICE_X82Y100_C5 = CLBLL_L_X54Y99_SLICE_X82Y99_DO6;
  assign CLBLL_L_X54Y100_SLICE_X82Y100_C6 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLL_L_X54Y100_SLICE_X82Y100_CE = CLBLM_L_X60Y98_SLICE_X91Y98_DQ;
  assign CLBLL_L_X54Y100_SLICE_X82Y100_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X54Y100_SLICE_X82Y100_D1 = CLBLL_L_X54Y99_SLICE_X82Y99_BO6;
  assign CLBLL_L_X54Y100_SLICE_X82Y100_D2 = CLBLL_L_X54Y100_SLICE_X83Y100_CO6;
  assign CLBLL_L_X54Y100_SLICE_X82Y100_D3 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLL_L_X54Y100_SLICE_X82Y100_D4 = CLBLL_L_X54Y100_SLICE_X82Y100_AO5;
  assign CLBLL_L_X54Y100_SLICE_X82Y100_D5 = CLBLL_L_X54Y99_SLICE_X82Y99_AO6;
  assign CLBLL_L_X54Y100_SLICE_X82Y100_D6 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLL_L_X54Y100_SLICE_X82Y100_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLL_L_X54Y100_SLICE_X83Y100_A1 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLL_L_X54Y100_SLICE_X83Y100_A2 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLL_L_X54Y100_SLICE_X83Y100_A3 = CLBLM_R_X49Y107_SLICE_X75Y107_DQ;
  assign CLBLL_L_X54Y100_SLICE_X83Y100_A4 = CLBLM_R_X49Y108_SLICE_X75Y108_DQ;
  assign CLBLL_L_X54Y100_SLICE_X83Y100_A5 = CLBLM_L_X56Y97_SLICE_X84Y97_CO5;
  assign CLBLL_L_X54Y100_SLICE_X83Y100_A6 = 1'b1;
  assign CLBLL_L_X54Y100_SLICE_X83Y100_B1 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLL_L_X54Y100_SLICE_X83Y100_B2 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLL_L_X54Y100_SLICE_X83Y100_B3 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLL_L_X54Y100_SLICE_X83Y100_B4 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign CLBLL_L_X54Y100_SLICE_X83Y100_B5 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLL_L_X54Y100_SLICE_X83Y100_B6 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLL_L_X54Y100_SLICE_X83Y100_C1 = CLBLL_L_X54Y99_SLICE_X82Y99_AO6;
  assign CLBLL_L_X54Y100_SLICE_X83Y100_C2 = CLBLM_R_X53Y99_SLICE_X80Y99_AO5;
  assign CLBLL_L_X54Y100_SLICE_X83Y100_C3 = CLBLL_L_X54Y99_SLICE_X83Y99_CO6;
  assign CLBLL_L_X54Y100_SLICE_X83Y100_C4 = CLBLM_R_X49Y107_SLICE_X75Y107_DQ;
  assign CLBLL_L_X54Y100_SLICE_X83Y100_C5 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLL_L_X54Y100_SLICE_X83Y100_C6 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLL_L_X54Y100_SLICE_X83Y100_D1 = 1'b1;
  assign CLBLL_L_X54Y100_SLICE_X83Y100_D2 = 1'b1;
  assign CLBLL_L_X54Y100_SLICE_X83Y100_D3 = 1'b1;
  assign CLBLL_L_X54Y100_SLICE_X83Y100_D4 = 1'b1;
  assign CLBLL_L_X54Y100_SLICE_X83Y100_D5 = 1'b1;
  assign CLBLL_L_X54Y100_SLICE_X83Y100_D6 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_A1 = CLBLM_R_X49Y104_SLICE_X75Y104_AQ;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_A2 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_A3 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_A4 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_A5 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_A6 = CLBLM_L_X64Y102_SLICE_X97Y102_B_XOR;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_B1 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_B2 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_B3 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_B4 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_B5 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_B6 = 1'b1;
  assign RIOI3_X105Y125_OLOGIC_X1Y126_D1 = CLBLM_L_X64Y106_SLICE_X97Y106_CQ;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_C1 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_C2 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_C3 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_C4 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_C5 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_C6 = 1'b1;
  assign RIOI3_X105Y125_OLOGIC_X1Y126_T1 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_D1 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_D2 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_D3 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_D4 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_D5 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X95Y102_D6 = 1'b1;
  assign RIOI3_X105Y125_OLOGIC_X1Y125_D1 = CLBLM_L_X64Y106_SLICE_X97Y106_BQ;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_A1 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_A2 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_A3 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_A4 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_A5 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_A6 = 1'b1;
  assign RIOI3_X105Y125_OLOGIC_X1Y125_T1 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_B1 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_B2 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_B3 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_B4 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_B6 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_B5 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_C1 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_C2 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_C3 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_C4 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_C5 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_C6 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_D1 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_D2 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_D3 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_D4 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_D5 = 1'b1;
  assign CLBLM_R_X63Y102_SLICE_X94Y102_D6 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_A1 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_A2 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_A3 = CLBLM_R_X49Y107_SLICE_X75Y107_DQ;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_A4 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_A5 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_A6 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_B1 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_B2 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_B3 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_B4 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_B5 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_B6 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_BX = CLBLL_L_X54Y101_SLICE_X82Y101_AO5;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_C1 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_C2 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_C3 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_C4 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_C5 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_C6 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_CE = CLBLM_L_X56Y98_SLICE_X84Y98_DO6;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_D1 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_D2 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_D3 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_D4 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_D5 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_D6 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X82Y101_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_A1 = CLBLM_R_X53Y100_SLICE_X80Y100_AQ;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_A2 = CLBLM_R_X53Y101_SLICE_X81Y101_AQ;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_A3 = CLBLM_R_X53Y101_SLICE_X80Y101_BQ;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_A4 = CLBLL_L_X54Y100_SLICE_X82Y100_BQ;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_A5 = CLBLM_R_X53Y100_SLICE_X81Y100_AQ;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_A6 = CLBLM_R_X53Y100_SLICE_X80Y100_A5Q;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_B1 = CLBLM_R_X53Y100_SLICE_X80Y100_AQ;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_B2 = CLBLM_R_X53Y101_SLICE_X81Y101_AQ;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_B3 = CLBLM_R_X53Y100_SLICE_X81Y100_AQ;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_B4 = CLBLL_L_X54Y100_SLICE_X82Y100_BQ;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_B5 = CLBLM_R_X53Y101_SLICE_X80Y101_BQ;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_B6 = CLBLM_R_X53Y100_SLICE_X80Y100_A5Q;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_C1 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_C2 = CLBLM_R_X53Y100_SLICE_X80Y100_A5Q;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_C3 = CLBLM_R_X53Y100_SLICE_X80Y100_AQ;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_C4 = CLBLM_R_X53Y101_SLICE_X80Y101_BQ;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_C5 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_C6 = CLBLM_R_X53Y101_SLICE_X81Y101_AQ;
  assign LIOB33_X0Y123_IOB_X0Y124_O = CLBLM_R_X49Y109_SLICE_X74Y109_DQ;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_D1 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_D2 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_D3 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_D4 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_D5 = 1'b1;
  assign CLBLL_L_X54Y101_SLICE_X83Y101_D6 = 1'b1;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_A1 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_A2 = CLBLM_R_X65Y103_SLICE_X99Y103_BQ;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_A3 = CLBLM_L_X64Y109_SLICE_X96Y109_AQ;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_A4 = 1'b1;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_A5 = CLBLL_R_X57Y103_SLICE_X86Y103_AQ;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_A6 = CLBLL_R_X57Y103_SLICE_X86Y103_A5Q;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_B1 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_B2 = 1'b1;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_B3 = CLBLM_L_X64Y99_SLICE_X96Y99_BQ;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_B4 = CLBLM_L_X64Y106_SLICE_X96Y106_BQ;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_B5 = CLBLL_R_X57Y103_SLICE_X86Y103_AQ;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_B6 = CLBLL_R_X57Y103_SLICE_X86Y103_A5Q;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_C1 = CLBLL_R_X57Y103_SLICE_X86Y103_AQ;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_C2 = CLBLL_R_X57Y103_SLICE_X86Y103_A5Q;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_C3 = CLBLM_L_X64Y98_SLICE_X96Y98_AQ;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_C4 = 1'b1;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_C5 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_C6 = CLBLM_L_X64Y107_SLICE_X96Y107_AQ;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_CE = CLBLM_L_X62Y105_SLICE_X93Y105_DO6;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_D1 = CLBLM_R_X49Y107_SLICE_X75Y107_CQ;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_D2 = CLBLM_L_X64Y103_SLICE_X97Y103_D_XOR;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_D3 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_D4 = 1'b1;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_D5 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_D6 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_R_X63Y103_SLICE_X95Y103_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_A1 = 1'b1;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_A2 = CLBLM_R_X49Y107_SLICE_X74Y107_AQ;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_A3 = CLBLM_L_X62Y107_SLICE_X93Y107_BO6;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_A4 = CLBLM_L_X64Y107_SLICE_X96Y107_AQ;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_A5 = CLBLM_R_X63Y104_SLICE_X94Y104_AQ;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_A6 = CLBLM_L_X62Y107_SLICE_X93Y107_AO6;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_B1 = 1'b1;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_B2 = 1'b1;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_B3 = 1'b1;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_B4 = 1'b1;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_B5 = 1'b1;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_B6 = 1'b1;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_C1 = 1'b1;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_C2 = 1'b1;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_C3 = 1'b1;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_C4 = 1'b1;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_C5 = 1'b1;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_C6 = 1'b1;
  assign CLBLM_R_X59Y98_SLICE_X89Y98_A3 = CLBLL_R_X57Y98_SLICE_X87Y98_AQ;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_D1 = 1'b1;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_D2 = 1'b1;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_D3 = 1'b1;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_D4 = 1'b1;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_D5 = 1'b1;
  assign CLBLM_R_X63Y103_SLICE_X94Y103_D6 = 1'b1;
  assign CLBLM_R_X59Y98_SLICE_X89Y98_A4 = CLBLL_R_X57Y98_SLICE_X87Y98_BQ;
  assign CLBLM_R_X59Y98_SLICE_X89Y98_A5 = CLBLM_L_X50Y105_SLICE_X77Y105_AQ;
  assign CLBLL_L_X54Y102_SLICE_X82Y102_A1 = CLBLM_R_X49Y106_SLICE_X75Y106_DQ;
  assign CLBLL_L_X54Y102_SLICE_X82Y102_A2 = CLBLM_R_X49Y104_SLICE_X75Y104_BQ;
  assign CLBLL_L_X54Y102_SLICE_X82Y102_A3 = CLBLM_R_X49Y107_SLICE_X75Y107_CQ;
  assign CLBLL_L_X54Y102_SLICE_X82Y102_A4 = CLBLM_R_X49Y106_SLICE_X75Y106_CQ;
  assign CLBLL_L_X54Y102_SLICE_X82Y102_A5 = CLBLM_R_X49Y104_SLICE_X75Y104_CQ;
  assign CLBLL_L_X54Y102_SLICE_X82Y102_A6 = 1'b1;
  assign CLBLL_L_X54Y102_SLICE_X82Y102_B1 = CLBLM_R_X49Y106_SLICE_X75Y106_DQ;
  assign CLBLL_L_X54Y102_SLICE_X82Y102_B2 = CLBLM_R_X49Y106_SLICE_X75Y106_CQ;
  assign CLBLL_L_X54Y102_SLICE_X82Y102_B3 = CLBLM_R_X49Y107_SLICE_X75Y107_CQ;
  assign CLBLL_L_X54Y102_SLICE_X82Y102_B4 = CLBLM_R_X49Y104_SLICE_X75Y104_CQ;
  assign CLBLL_L_X54Y102_SLICE_X82Y102_B5 = CLBLM_R_X49Y104_SLICE_X75Y104_BQ;
  assign CLBLL_L_X54Y102_SLICE_X82Y102_B6 = CLBLL_L_X54Y102_SLICE_X82Y102_CO6;
  assign CLBLM_R_X59Y98_SLICE_X89Y98_B5 = CLBLM_R_X49Y106_SLICE_X74Y106_AQ;
  assign CLBLM_R_X59Y98_SLICE_X89Y98_B6 = 1'b1;
  assign CLBLL_L_X54Y102_SLICE_X82Y102_C1 = CLBLM_R_X49Y107_SLICE_X75Y107_DQ;
  assign CLBLL_L_X54Y102_SLICE_X82Y102_C2 = CLBLM_L_X56Y97_SLICE_X84Y97_CO5;
  assign CLBLL_L_X54Y102_SLICE_X82Y102_C3 = CLBLM_R_X49Y104_SLICE_X75Y104_DQ;
  assign CLBLL_L_X54Y102_SLICE_X82Y102_C4 = CLBLM_R_X49Y108_SLICE_X75Y108_DQ;
  assign CLBLL_L_X54Y102_SLICE_X82Y102_C5 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLL_L_X54Y102_SLICE_X82Y102_C6 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLL_L_X54Y102_SLICE_X82Y102_D1 = 1'b1;
  assign CLBLL_L_X54Y102_SLICE_X82Y102_D2 = 1'b1;
  assign CLBLL_L_X54Y102_SLICE_X82Y102_D3 = 1'b1;
  assign CLBLL_L_X54Y102_SLICE_X82Y102_D4 = 1'b1;
  assign CLBLL_L_X54Y102_SLICE_X82Y102_D5 = 1'b1;
  assign CLBLL_L_X54Y102_SLICE_X82Y102_D6 = 1'b1;
  assign CLBLM_R_X59Y98_SLICE_X89Y98_C4 = CLBLM_L_X60Y98_SLICE_X90Y98_DO6;
  assign LIOB33_X0Y125_IOB_X0Y126_O = CLBLM_R_X49Y111_SLICE_X74Y111_AQ;
  assign LIOB33_X0Y125_IOB_X0Y125_O = CLBLM_R_X49Y107_SLICE_X74Y107_AQ;
  assign CLBLL_L_X54Y102_SLICE_X83Y102_A1 = 1'b1;
  assign CLBLL_L_X54Y102_SLICE_X83Y102_A2 = 1'b1;
  assign CLBLL_L_X54Y102_SLICE_X83Y102_A3 = 1'b1;
  assign CLBLL_L_X54Y102_SLICE_X83Y102_A4 = 1'b1;
  assign CLBLL_L_X54Y102_SLICE_X83Y102_A5 = 1'b1;
  assign CLBLL_L_X54Y102_SLICE_X83Y102_A6 = 1'b1;
  assign CLBLL_L_X54Y102_SLICE_X83Y102_B1 = 1'b1;
  assign CLBLL_L_X54Y102_SLICE_X83Y102_B2 = 1'b1;
  assign CLBLL_L_X54Y102_SLICE_X83Y102_B3 = 1'b1;
  assign CLBLL_L_X54Y102_SLICE_X83Y102_B4 = 1'b1;
  assign CLBLL_L_X54Y102_SLICE_X83Y102_B5 = 1'b1;
  assign CLBLL_L_X54Y102_SLICE_X83Y102_B6 = 1'b1;
  assign CLBLL_L_X54Y102_SLICE_X83Y102_C1 = 1'b1;
  assign CLBLL_L_X54Y102_SLICE_X83Y102_C2 = 1'b1;
  assign CLBLL_L_X54Y102_SLICE_X83Y102_C3 = 1'b1;
  assign CLBLL_L_X54Y102_SLICE_X83Y102_C4 = 1'b1;
  assign CLBLL_L_X54Y102_SLICE_X83Y102_C5 = 1'b1;
  assign CLBLL_L_X54Y102_SLICE_X83Y102_C6 = 1'b1;
  assign CLBLL_L_X54Y102_SLICE_X83Y102_D1 = 1'b1;
  assign CLBLL_L_X54Y102_SLICE_X83Y102_D2 = 1'b1;
  assign CLBLL_L_X54Y102_SLICE_X83Y102_D3 = 1'b1;
  assign CLBLL_L_X54Y102_SLICE_X83Y102_D4 = 1'b1;
  assign CLBLL_L_X54Y102_SLICE_X83Y102_D5 = 1'b1;
  assign CLBLL_L_X54Y102_SLICE_X83Y102_D6 = 1'b1;
  assign CLBLM_R_X59Y98_SLICE_X89Y98_D2 = 1'b1;
  assign CLBLM_R_X63Y104_SLICE_X95Y104_A1 = CLBLM_L_X64Y104_SLICE_X97Y104_A_XOR;
  assign CLBLM_R_X63Y104_SLICE_X95Y104_A2 = CLBLM_L_X56Y97_SLICE_X84Y97_BQ;
  assign CLBLM_R_X63Y104_SLICE_X95Y104_A3 = CLBLM_L_X60Y97_SLICE_X90Y97_AQ;
  assign CLBLM_R_X63Y104_SLICE_X95Y104_A4 = CLBLM_L_X60Y97_SLICE_X90Y97_CQ;
  assign CLBLM_R_X63Y104_SLICE_X95Y104_A5 = CLBLM_R_X49Y108_SLICE_X75Y108_DQ;
  assign CLBLM_R_X63Y104_SLICE_X95Y104_A6 = 1'b1;
  assign CLBLM_R_X63Y104_SLICE_X95Y104_B1 = 1'b1;
  assign CLBLM_R_X63Y104_SLICE_X95Y104_B2 = 1'b1;
  assign CLBLM_R_X63Y104_SLICE_X95Y104_B3 = 1'b1;
  assign CLBLM_R_X63Y104_SLICE_X95Y104_B4 = 1'b1;
  assign CLBLM_R_X63Y104_SLICE_X95Y104_B5 = 1'b1;
  assign CLBLM_R_X63Y104_SLICE_X95Y104_B6 = 1'b1;
  assign CLBLM_R_X63Y104_SLICE_X95Y104_C1 = 1'b1;
  assign CLBLM_R_X63Y104_SLICE_X95Y104_C2 = 1'b1;
  assign CLBLM_R_X63Y104_SLICE_X95Y104_C3 = 1'b1;
  assign CLBLM_R_X63Y104_SLICE_X95Y104_C4 = 1'b1;
  assign CLBLM_R_X63Y104_SLICE_X95Y104_C5 = 1'b1;
  assign CLBLM_R_X63Y104_SLICE_X95Y104_C6 = 1'b1;
  assign CLBLM_R_X63Y104_SLICE_X95Y104_D1 = 1'b1;
  assign CLBLM_R_X63Y104_SLICE_X95Y104_D2 = 1'b1;
  assign CLBLM_R_X63Y104_SLICE_X95Y104_D3 = 1'b1;
  assign CLBLM_R_X63Y104_SLICE_X95Y104_D4 = 1'b1;
  assign CLBLM_R_X63Y104_SLICE_X95Y104_D5 = 1'b1;
  assign CLBLM_R_X63Y104_SLICE_X95Y104_D6 = 1'b1;
  assign CLBLM_R_X63Y104_SLICE_X94Y104_A1 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X63Y104_SLICE_X94Y104_A2 = CLBLM_L_X62Y105_SLICE_X92Y105_BO5;
  assign CLBLM_R_X63Y104_SLICE_X94Y104_A3 = CLBLM_R_X63Y104_SLICE_X94Y104_AQ;
  assign CLBLM_R_X63Y104_SLICE_X94Y104_A4 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X63Y104_SLICE_X94Y104_A5 = CLBLM_R_X63Y104_SLICE_X94Y104_CO6;
  assign CLBLM_R_X63Y104_SLICE_X94Y104_A6 = CLBLM_R_X63Y105_SLICE_X95Y105_A_XOR;
  assign CLBLM_R_X63Y104_SLICE_X94Y104_B1 = CLBLM_R_X63Y104_SLICE_X94Y104_DO6;
  assign CLBLM_R_X63Y104_SLICE_X94Y104_B2 = CLBLM_R_X63Y104_SLICE_X94Y104_BQ;
  assign CLBLM_R_X63Y104_SLICE_X94Y104_B3 = CLBLM_R_X63Y105_SLICE_X95Y105_D_XOR;
  assign CLBLM_R_X63Y104_SLICE_X94Y104_B4 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X63Y104_SLICE_X94Y104_B5 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X63Y104_SLICE_X94Y104_B6 = CLBLM_L_X62Y105_SLICE_X92Y105_BO5;
  assign CLBLM_R_X63Y104_SLICE_X94Y104_C1 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X63Y104_SLICE_X94Y104_C2 = CLBLM_L_X62Y105_SLICE_X93Y105_AO6;
  assign CLBLM_R_X63Y104_SLICE_X94Y104_C3 = CLBLM_L_X50Y105_SLICE_X77Y105_AQ;
  assign CLBLM_R_X63Y104_SLICE_X94Y104_C4 = CLBLM_R_X63Y105_SLICE_X95Y105_A_XOR;
  assign CLBLM_R_X63Y104_SLICE_X94Y104_C5 = CLBLM_R_X63Y105_SLICE_X94Y105_B_XOR;
  assign CLBLM_R_X63Y104_SLICE_X94Y104_C6 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X63Y104_SLICE_X94Y104_CE = CLBLM_L_X62Y100_SLICE_X92Y100_CO6;
  assign CLBLM_R_X63Y104_SLICE_X94Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X63Y104_SLICE_X94Y104_D1 = CLBLM_R_X63Y105_SLICE_X95Y105_D_XOR;
  assign CLBLM_R_X63Y104_SLICE_X94Y104_D2 = CLBLM_L_X62Y105_SLICE_X93Y105_AO6;
  assign CLBLM_R_X63Y104_SLICE_X94Y104_D3 = CLBLM_L_X50Y106_SLICE_X76Y106_AQ;
  assign CLBLM_R_X63Y104_SLICE_X94Y104_D4 = CLBLM_R_X63Y106_SLICE_X94Y106_A_XOR;
  assign CLBLM_R_X63Y104_SLICE_X94Y104_D5 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X63Y104_SLICE_X94Y104_D6 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X63Y104_SLICE_X94Y104_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLL_L_X54Y103_SLICE_X82Y103_A1 = CLBLM_R_X49Y104_SLICE_X75Y104_AQ;
  assign CLBLL_L_X54Y103_SLICE_X82Y103_A2 = CLBLM_R_X49Y104_SLICE_X74Y104_AQ;
  assign CLBLL_L_X54Y103_SLICE_X82Y103_A3 = CLBLM_R_X49Y106_SLICE_X75Y106_DQ;
  assign CLBLL_L_X54Y103_SLICE_X82Y103_A4 = CLBLM_L_X56Y104_SLICE_X84Y104_AQ;
  assign CLBLL_L_X54Y103_SLICE_X82Y103_A5 = CLBLL_L_X54Y102_SLICE_X82Y102_AO6;
  assign CLBLL_L_X54Y103_SLICE_X82Y103_A6 = CLBLL_L_X54Y102_SLICE_X82Y102_CO6;
  assign CLBLL_L_X54Y103_SLICE_X82Y103_B1 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X82Y103_B2 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X82Y103_B3 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X82Y103_B4 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X82Y103_B5 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X82Y103_B6 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X82Y103_C1 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X82Y103_C2 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X82Y103_C3 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X82Y103_C4 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X82Y103_C5 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X82Y103_C6 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X82Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_D1 = CLBLM_R_X59Y102_SLICE_X88Y102_AQ;
  assign CLBLL_L_X54Y103_SLICE_X82Y103_D1 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X82Y103_D2 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X82Y103_D3 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X82Y103_D4 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X82Y103_D5 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X82Y103_D6 = 1'b1;
  assign LIOB33_X0Y127_IOB_X0Y127_O = CLBLM_R_X49Y111_SLICE_X74Y111_BQ;
  assign LIOB33_X0Y127_IOB_X0Y128_O = CLBLM_R_X49Y109_SLICE_X74Y109_AQ;
  assign CLBLL_L_X54Y103_SLICE_X82Y103_SR = CLBLM_R_X15Y122_SLICE_X20Y122_AO6;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_T1 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X83Y103_A1 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X83Y103_A2 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X83Y103_A3 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X83Y103_A4 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X83Y103_A5 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X83Y103_A6 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X83Y103_B1 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X83Y103_B2 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X83Y103_B3 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X83Y103_B4 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X83Y103_B5 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X83Y103_B6 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X83Y103_C1 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X83Y103_C2 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X83Y103_C3 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X83Y103_C4 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X83Y103_C5 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X83Y103_C6 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X83Y103_D1 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X83Y103_D2 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X83Y103_D3 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X83Y103_D4 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X83Y103_D5 = 1'b1;
  assign CLBLL_L_X54Y103_SLICE_X83Y103_D6 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_A1 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_A2 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_A3 = CLBLM_R_X63Y104_SLICE_X94Y104_AQ;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_A4 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_A5 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_A6 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_AX = CLBLM_L_X62Y105_SLICE_X92Y105_CQ;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_B1 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_B2 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_B3 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_B4 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_B5 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_B6 = CLBLM_L_X64Y105_SLICE_X96Y105_AQ;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_BX = 1'b0;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_C1 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_C2 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_C3 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_C4 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_C5 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_C6 = CLBLM_L_X64Y105_SLICE_X97Y105_AQ;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_D = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_CX = 1'b0;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_D1 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_D2 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_D3 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_D4 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_D5 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_D6 = CLBLM_R_X63Y104_SLICE_X94Y104_BQ;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_DX = 1'b0;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_A1 = CLBLM_L_X62Y105_SLICE_X92Y105_AO5;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_A2 = CLBLM_L_X62Y105_SLICE_X92Y105_CQ;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_A3 = CLBLM_R_X59Y101_SLICE_X89Y101_AQ;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_A4 = CLBLM_R_X59Y103_SLICE_X89Y103_A5Q;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_A5 = CLBLL_R_X57Y102_SLICE_X86Y102_AQ;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_A6 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_AX = CLBLM_L_X62Y105_SLICE_X92Y105_CQ;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_B1 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_B2 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_B3 = CLBLM_R_X63Y104_SLICE_X94Y104_AQ;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_B4 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_B5 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_B6 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_BX = CLBLM_R_X63Y104_SLICE_X94Y104_AQ;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_C1 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_C2 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_C3 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_C4 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_C5 = CLBLM_L_X64Y105_SLICE_X96Y105_AQ;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_C6 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_CE = CLBLM_L_X62Y100_SLICE_X92Y100_DO6;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_CX = CLBLM_L_X64Y105_SLICE_X96Y105_AQ;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_D1 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_D2 = CLBLM_L_X64Y105_SLICE_X97Y105_AQ;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_D3 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_D4 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_D5 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_D6 = 1'b1;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_DX = CLBLM_L_X64Y105_SLICE_X97Y105_AQ;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLL_L_X54Y104_SLICE_X82Y104_A1 = CLBLM_L_X56Y101_SLICE_X85Y101_BQ;
  assign CLBLL_L_X54Y104_SLICE_X82Y104_A2 = CLBLM_L_X56Y101_SLICE_X85Y101_CQ;
  assign CLBLL_L_X54Y104_SLICE_X82Y104_A3 = CLBLL_R_X57Y100_SLICE_X86Y100_CQ;
  assign CLBLL_L_X54Y104_SLICE_X82Y104_A4 = CLBLL_R_X57Y101_SLICE_X87Y101_AQ;
  assign CLBLL_L_X54Y104_SLICE_X82Y104_A5 = CLBLL_R_X57Y100_SLICE_X87Y100_AQ;
  assign CLBLL_L_X54Y104_SLICE_X82Y104_A6 = CLBLL_R_X57Y100_SLICE_X86Y100_DQ;
  assign CLBLL_L_X54Y104_SLICE_X82Y104_B1 = CLBLM_L_X56Y101_SLICE_X85Y101_BQ;
  assign CLBLL_L_X54Y104_SLICE_X82Y104_B2 = CLBLM_L_X56Y101_SLICE_X85Y101_CQ;
  assign CLBLL_L_X54Y104_SLICE_X82Y104_B3 = CLBLL_R_X57Y100_SLICE_X86Y100_CQ;
  assign CLBLL_L_X54Y104_SLICE_X82Y104_B4 = CLBLL_R_X57Y100_SLICE_X87Y100_BQ;
  assign CLBLL_L_X54Y104_SLICE_X82Y104_B5 = CLBLL_R_X57Y100_SLICE_X86Y100_DQ;
  assign CLBLL_L_X54Y104_SLICE_X82Y104_B6 = CLBLL_R_X57Y101_SLICE_X87Y101_AQ;
  assign LIOB33_X0Y129_IOB_X0Y129_O = CLBLM_R_X49Y109_SLICE_X74Y109_BQ;
  assign LIOB33_X0Y129_IOB_X0Y130_O = CLBLM_R_X49Y111_SLICE_X74Y111_CQ;
  assign CLBLL_L_X54Y104_SLICE_X82Y104_C1 = 1'b1;
  assign CLBLL_L_X54Y104_SLICE_X82Y104_C2 = 1'b1;
  assign CLBLL_L_X54Y104_SLICE_X82Y104_C3 = 1'b1;
  assign CLBLL_L_X54Y104_SLICE_X82Y104_C4 = 1'b1;
  assign CLBLL_L_X54Y104_SLICE_X82Y104_C5 = 1'b1;
  assign CLBLL_L_X54Y104_SLICE_X82Y104_C6 = 1'b1;
  assign CLBLL_L_X54Y104_SLICE_X82Y104_D1 = 1'b1;
  assign CLBLL_L_X54Y104_SLICE_X82Y104_D2 = 1'b1;
  assign CLBLL_L_X54Y104_SLICE_X82Y104_D3 = 1'b1;
  assign CLBLL_L_X54Y104_SLICE_X82Y104_D4 = 1'b1;
  assign CLBLL_L_X54Y104_SLICE_X82Y104_D5 = 1'b1;
  assign CLBLL_L_X54Y104_SLICE_X82Y104_D6 = 1'b1;
  assign CLBLL_L_X54Y104_SLICE_X83Y104_A1 = 1'b1;
  assign CLBLL_L_X54Y104_SLICE_X83Y104_A2 = 1'b1;
  assign CLBLL_L_X54Y104_SLICE_X83Y104_A3 = 1'b1;
  assign CLBLL_L_X54Y104_SLICE_X83Y104_A4 = 1'b1;
  assign CLBLL_L_X54Y104_SLICE_X83Y104_A5 = 1'b1;
  assign CLBLL_L_X54Y104_SLICE_X83Y104_A6 = 1'b1;
  assign CLBLL_L_X54Y104_SLICE_X83Y104_B1 = 1'b1;
  assign CLBLL_L_X54Y104_SLICE_X83Y104_B2 = 1'b1;
  assign CLBLL_L_X54Y104_SLICE_X83Y104_B3 = 1'b1;
  assign CLBLL_L_X54Y104_SLICE_X83Y104_B4 = 1'b1;
  assign CLBLL_L_X54Y104_SLICE_X83Y104_B5 = 1'b1;
  assign CLBLL_L_X54Y104_SLICE_X83Y104_B6 = 1'b1;
  assign CLBLL_L_X54Y104_SLICE_X83Y104_C1 = 1'b1;
  assign CLBLL_L_X54Y104_SLICE_X83Y104_C2 = 1'b1;
  assign CLBLL_L_X54Y104_SLICE_X83Y104_C3 = 1'b1;
  assign CLBLL_L_X54Y104_SLICE_X83Y104_C4 = 1'b1;
  assign CLBLL_L_X54Y104_SLICE_X83Y104_C5 = 1'b1;
  assign CLBLL_L_X54Y104_SLICE_X83Y104_C6 = 1'b1;
  assign CLBLL_L_X54Y104_SLICE_X83Y104_D1 = 1'b1;
  assign CLBLL_L_X54Y104_SLICE_X83Y104_D2 = 1'b1;
  assign CLBLL_L_X54Y104_SLICE_X83Y104_D3 = 1'b1;
  assign CLBLL_L_X54Y104_SLICE_X83Y104_D4 = 1'b1;
  assign CLBLL_L_X54Y104_SLICE_X83Y104_D5 = 1'b1;
  assign CLBLL_L_X54Y104_SLICE_X83Y104_D6 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_A1 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_A2 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_A3 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_A4 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_A5 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_A6 = CLBLM_L_X62Y105_SLICE_X93Y105_BQ;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_AX = 1'b0;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_B1 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_B2 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_B3 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_B4 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_B5 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_B6 = CLBLM_L_X64Y106_SLICE_X96Y106_AQ;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_BX = 1'b0;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_C1 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_C2 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_C3 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_C4 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_C5 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_C6 = CLBLM_L_X64Y106_SLICE_X96Y106_BQ;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_CIN = CLBLM_R_X63Y105_SLICE_X95Y105_COUT;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_CX = 1'b0;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_D1 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_D2 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_D3 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_D4 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_D5 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_D6 = CLBLM_L_X64Y107_SLICE_X97Y107_BQ;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_DX = 1'b0;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_A1 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_A2 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_A3 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_A4 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_A5 = CLBLM_R_X63Y104_SLICE_X94Y104_BQ;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_A6 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_AX = CLBLM_R_X63Y104_SLICE_X94Y104_BQ;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_B1 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_B2 = CLBLM_L_X62Y105_SLICE_X93Y105_BQ;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_B3 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_B4 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_B5 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_B6 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_BX = CLBLM_L_X62Y105_SLICE_X93Y105_BQ;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_C1 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_C2 = CLBLM_L_X64Y106_SLICE_X96Y106_AQ;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_C3 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_C4 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_C5 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_C6 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_CIN = CLBLM_R_X63Y105_SLICE_X94Y105_COUT;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_CX = CLBLM_L_X64Y106_SLICE_X96Y106_AQ;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_D1 = CLBLM_L_X64Y106_SLICE_X96Y106_BQ;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_D2 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_D3 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_D4 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_D5 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_D6 = 1'b1;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_DX = CLBLM_L_X64Y106_SLICE_X96Y106_BQ;
  assign LIOB33_X0Y131_IOB_X0Y132_O = CLBLM_R_X49Y109_SLICE_X74Y109_DQ;
  assign LIOB33_X0Y131_IOB_X0Y131_O = CLBLM_R_X49Y109_SLICE_X74Y109_CQ;
  assign CLBLM_L_X56Y105_SLICE_X84Y105_C1 = CLBLL_L_X54Y101_SLICE_X83Y101_BO6;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_A1 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_A2 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_A3 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_A4 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_A5 = CLBLM_R_X53Y103_SLICE_X81Y103_D_XOR;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_A6 = CLBLM_R_X53Y106_SLICE_X81Y106_A_XOR;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_AX = CLBLM_R_X53Y103_SLICE_X81Y103_D_XOR;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_B1 = CLBLM_R_X53Y106_SLICE_X81Y106_B_XOR;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_B2 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_B3 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_B4 = CLBLM_R_X53Y104_SLICE_X81Y104_A_XOR;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_B5 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_B6 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_BX = CLBLM_R_X53Y104_SLICE_X81Y104_A_XOR;
  assign CLBLM_L_X56Y105_SLICE_X84Y105_C2 = CLBLM_L_X56Y105_SLICE_X84Y105_CQ;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_C1 = CLBLM_R_X53Y104_SLICE_X81Y104_B_XOR;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_C2 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_C3 = CLBLM_R_X53Y106_SLICE_X81Y106_C_XOR;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_C4 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_C5 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_C6 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_CX = CLBLM_R_X53Y104_SLICE_X81Y104_B_XOR;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_D1 = CLBLM_R_X53Y104_SLICE_X81Y104_C_XOR;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_D2 = CLBLM_R_X53Y106_SLICE_X81Y106_D_XOR;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_D3 = CLBLL_R_X57Y100_SLICE_X86Y100_AQ;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_D4 = CLBLL_R_X57Y101_SLICE_X87Y101_DQ;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_D5 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_D6 = 1'b1;
  assign CLBLM_L_X56Y105_SLICE_X84Y105_C3 = CLBLM_L_X50Y107_SLICE_X76Y107_BQ;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_A1 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_A2 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_A3 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_A4 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_A5 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_A6 = 1'b1;
  assign CLBLM_L_X56Y105_SLICE_X84Y105_C4 = CLBLM_L_X60Y99_SLICE_X90Y99_AO5;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_B1 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_B2 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_B3 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_B4 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_B5 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_B6 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_C1 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_C2 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_C3 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_C4 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_C5 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_C6 = 1'b1;
  assign CLBLM_L_X56Y105_SLICE_X84Y105_C5 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_D1 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_D2 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_D3 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_D4 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_D5 = 1'b1;
  assign CLBLL_L_X54Y105_SLICE_X83Y105_D6 = 1'b1;
  assign CLBLM_L_X56Y105_SLICE_X84Y105_C6 = CLBLL_L_X54Y107_SLICE_X82Y107_D_XOR;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_D1 = CLBLM_L_X62Y103_SLICE_X92Y103_AQ;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_T1 = 1'b1;
  assign CLBLM_L_X56Y105_SLICE_X84Y105_CE = CLBLM_L_X56Y103_SLICE_X85Y103_CO6;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_D1 = CLBLM_L_X62Y104_SLICE_X93Y104_AQ;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_T1 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_A1 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_A2 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_A3 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_A4 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_A5 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_A6 = CLBLM_L_X64Y107_SLICE_X96Y107_AQ;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_AX = 1'b0;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_B1 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_B2 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_B3 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_B4 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_B5 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_B6 = CLBLM_L_X64Y107_SLICE_X96Y107_BQ;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_BX = 1'b0;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_C1 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_C2 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_C3 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_C4 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_C5 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_C6 = CLBLM_L_X64Y107_SLICE_X97Y107_AQ;
  assign CLBLM_L_X56Y105_SLICE_X84Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_CIN = CLBLM_R_X63Y106_SLICE_X95Y106_COUT;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_CX = 1'b0;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_D1 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_D2 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_D3 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_D4 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_D5 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_D6 = CLBLM_L_X64Y108_SLICE_X96Y108_AQ;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_DX = 1'b0;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_A1 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_A2 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_A3 = CLBLM_L_X64Y107_SLICE_X97Y107_BQ;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_A4 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_A5 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_A6 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_AX = CLBLM_L_X64Y107_SLICE_X97Y107_BQ;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_B1 = CLBLM_L_X64Y107_SLICE_X96Y107_AQ;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_B2 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_B3 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_B4 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_B5 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_B6 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_BX = CLBLM_L_X64Y107_SLICE_X96Y107_AQ;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_C1 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_C2 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_C3 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_C4 = CLBLM_L_X64Y107_SLICE_X96Y107_BQ;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_C5 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_C6 = 1'b1;
  assign LIOB33_X0Y133_IOB_X0Y133_O = CLBLM_R_X49Y107_SLICE_X74Y107_AQ;
  assign LIOB33_X0Y133_IOB_X0Y134_O = CLBLM_R_X49Y111_SLICE_X74Y111_AQ;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_CIN = CLBLM_R_X63Y106_SLICE_X94Y106_COUT;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_CX = CLBLM_L_X64Y107_SLICE_X96Y107_BQ;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_D1 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_D2 = CLBLM_L_X64Y107_SLICE_X97Y107_AQ;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_D3 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_D4 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_D5 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_D6 = 1'b1;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_DX = CLBLM_L_X64Y107_SLICE_X97Y107_AQ;
  assign CLBLL_L_X54Y106_SLICE_X82Y106_A1 = CLBLM_R_X53Y106_SLICE_X81Y106_D_XOR;
  assign CLBLL_L_X54Y106_SLICE_X82Y106_A2 = CLBLL_R_X57Y101_SLICE_X87Y101_DQ;
  assign CLBLL_L_X54Y106_SLICE_X82Y106_A3 = CLBLL_L_X54Y106_SLICE_X83Y106_CO6;
  assign CLBLL_L_X54Y106_SLICE_X82Y106_A4 = CLBLL_R_X57Y100_SLICE_X86Y100_BQ;
  assign CLBLL_L_X54Y106_SLICE_X82Y106_A5 = CLBLM_R_X53Y104_SLICE_X81Y104_C_XOR;
  assign CLBLL_L_X54Y106_SLICE_X82Y106_A6 = 1'b1;
  assign CLBLL_L_X54Y106_SLICE_X82Y106_AX = CLBLL_L_X54Y106_SLICE_X83Y106_CO6;
  assign CLBLL_L_X54Y106_SLICE_X82Y106_B1 = CLBLL_R_X57Y99_SLICE_X86Y99_BQ;
  assign CLBLL_L_X54Y106_SLICE_X82Y106_B2 = CLBLL_R_X57Y100_SLICE_X86Y100_AQ;
  assign CLBLL_L_X54Y106_SLICE_X82Y106_B3 = CLBLM_R_X53Y106_SLICE_X80Y106_BO6;
  assign CLBLL_L_X54Y106_SLICE_X82Y106_B4 = CLBLM_R_X53Y104_SLICE_X81Y104_D_XOR;
  assign CLBLL_L_X54Y106_SLICE_X82Y106_B5 = 1'b1;
  assign CLBLL_L_X54Y106_SLICE_X82Y106_B6 = CLBLM_R_X53Y107_SLICE_X81Y107_A_XOR;
  assign CLBLL_L_X54Y106_SLICE_X82Y106_BX = CLBLM_R_X53Y106_SLICE_X80Y106_BO6;
  assign CLBLL_L_X54Y106_SLICE_X82Y106_C1 = CLBLM_R_X53Y105_SLICE_X80Y105_AO6;
  assign CLBLL_L_X54Y106_SLICE_X82Y106_C2 = CLBLL_L_X54Y106_SLICE_X83Y106_AO6;
  assign CLBLL_L_X54Y106_SLICE_X82Y106_C3 = CLBLL_R_X57Y101_SLICE_X87Y101_DQ;
  assign CLBLL_L_X54Y106_SLICE_X82Y106_C4 = 1'b1;
  assign CLBLL_L_X54Y106_SLICE_X82Y106_C5 = CLBLL_R_X57Y100_SLICE_X87Y100_AQ;
  assign CLBLL_L_X54Y106_SLICE_X82Y106_C6 = CLBLM_R_X53Y106_SLICE_X80Y106_AO6;
  assign CLBLL_L_X54Y106_SLICE_X82Y106_CIN = CLBLL_L_X54Y105_SLICE_X82Y105_COUT;
  assign CLBLL_L_X54Y106_SLICE_X82Y106_CX = CLBLM_R_X53Y105_SLICE_X80Y105_AO6;
  assign CLBLL_L_X54Y106_SLICE_X82Y106_D1 = CLBLL_R_X57Y101_SLICE_X87Y101_AQ;
  assign CLBLL_L_X54Y106_SLICE_X82Y106_D2 = CLBLL_L_X54Y106_SLICE_X83Y106_AO5;
  assign CLBLL_L_X54Y106_SLICE_X82Y106_D3 = CLBLL_L_X54Y106_SLICE_X83Y106_BO6;
  assign CLBLL_L_X54Y106_SLICE_X82Y106_D4 = CLBLL_R_X57Y101_SLICE_X87Y101_DQ;
  assign CLBLL_L_X54Y106_SLICE_X82Y106_D5 = CLBLM_R_X53Y107_SLICE_X80Y107_BO5;
  assign CLBLL_L_X54Y106_SLICE_X82Y106_D6 = 1'b1;
  assign CLBLL_L_X54Y106_SLICE_X82Y106_DX = CLBLL_L_X54Y106_SLICE_X83Y106_BO6;
  assign CLBLL_L_X54Y106_SLICE_X83Y106_A1 = 1'b1;
  assign CLBLL_L_X54Y106_SLICE_X83Y106_A2 = CLBLM_L_X56Y101_SLICE_X85Y101_AQ;
  assign CLBLL_L_X54Y106_SLICE_X83Y106_A3 = CLBLM_R_X53Y107_SLICE_X81Y107_C_XOR;
  assign CLBLL_L_X54Y106_SLICE_X83Y106_A4 = CLBLM_R_X53Y105_SLICE_X81Y105_B_XOR;
  assign CLBLL_L_X54Y106_SLICE_X83Y106_A5 = CLBLL_R_X57Y99_SLICE_X86Y99_BQ;
  assign CLBLL_L_X54Y106_SLICE_X83Y106_A6 = 1'b1;
  assign CLBLL_L_X54Y106_SLICE_X83Y106_B1 = CLBLL_R_X57Y101_SLICE_X87Y101_DQ;
  assign CLBLL_L_X54Y106_SLICE_X83Y106_B2 = CLBLM_R_X53Y106_SLICE_X80Y106_AO6;
  assign CLBLL_L_X54Y106_SLICE_X83Y106_B3 = 1'b1;
  assign CLBLL_L_X54Y106_SLICE_X83Y106_B4 = CLBLL_R_X57Y100_SLICE_X87Y100_AQ;
  assign CLBLL_L_X54Y106_SLICE_X83Y106_B5 = CLBLL_L_X54Y106_SLICE_X83Y106_AO6;
  assign CLBLL_L_X54Y106_SLICE_X83Y106_B6 = 1'b1;
  assign CLBLL_L_X54Y106_SLICE_X83Y106_C1 = CLBLL_R_X57Y100_SLICE_X86Y100_AQ;
  assign CLBLL_L_X54Y106_SLICE_X83Y106_C2 = CLBLM_R_X53Y107_SLICE_X81Y107_A_XOR;
  assign CLBLL_L_X54Y106_SLICE_X83Y106_C3 = CLBLL_R_X57Y99_SLICE_X86Y99_BQ;
  assign CLBLL_L_X54Y106_SLICE_X83Y106_C4 = 1'b1;
  assign CLBLL_L_X54Y106_SLICE_X83Y106_C5 = 1'b1;
  assign CLBLL_L_X54Y106_SLICE_X83Y106_C6 = CLBLM_R_X53Y104_SLICE_X81Y104_D_XOR;
  assign CLBLL_L_X54Y106_SLICE_X83Y106_D1 = 1'b1;
  assign CLBLL_L_X54Y106_SLICE_X83Y106_D2 = CLBLL_R_X57Y101_SLICE_X87Y101_DQ;
  assign CLBLL_L_X54Y106_SLICE_X83Y106_D3 = CLBLM_R_X53Y107_SLICE_X80Y107_BO5;
  assign CLBLL_L_X54Y106_SLICE_X83Y106_D4 = CLBLL_L_X54Y106_SLICE_X83Y106_AO5;
  assign CLBLL_L_X54Y106_SLICE_X83Y106_D5 = CLBLL_R_X57Y101_SLICE_X87Y101_AQ;
  assign CLBLL_L_X54Y106_SLICE_X83Y106_D6 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X95Y108_A1 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X95Y108_A2 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X95Y108_A3 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X95Y108_A4 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X95Y108_A5 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X95Y108_A6 = CLBLM_L_X64Y108_SLICE_X97Y108_AQ;
  assign CLBLM_R_X63Y108_SLICE_X95Y108_AX = 1'b0;
  assign CLBLM_R_X63Y108_SLICE_X95Y108_B1 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X95Y108_B2 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X95Y108_B3 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X95Y108_B4 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X95Y108_B5 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X95Y108_B6 = CLBLM_R_X63Y110_SLICE_X94Y110_AQ;
  assign CLBLM_R_X63Y108_SLICE_X95Y108_BX = 1'b0;
  assign CLBLM_R_X63Y108_SLICE_X95Y108_C1 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X95Y108_C2 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X95Y108_C3 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X95Y108_C4 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X95Y108_C5 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X95Y108_C6 = CLBLM_L_X64Y108_SLICE_X96Y108_BQ;
  assign CLBLM_R_X63Y108_SLICE_X95Y108_CIN = CLBLM_R_X63Y107_SLICE_X95Y107_COUT;
  assign CLBLM_R_X63Y108_SLICE_X95Y108_CX = 1'b0;
  assign CLBLM_R_X63Y108_SLICE_X95Y108_D1 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X95Y108_D2 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X95Y108_D3 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X95Y108_D4 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X95Y108_D5 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X95Y108_D6 = CLBLM_L_X64Y109_SLICE_X96Y109_AQ;
  assign CLBLM_R_X63Y108_SLICE_X95Y108_DX = 1'b0;
  assign LIOB33_X0Y135_IOB_X0Y136_O = CLBLM_R_X49Y109_SLICE_X74Y109_AQ;
  assign LIOB33_X0Y135_IOB_X0Y135_O = CLBLM_R_X49Y111_SLICE_X74Y111_BQ;
  assign CLBLM_R_X63Y108_SLICE_X94Y108_A1 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X94Y108_A2 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X94Y108_A3 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X94Y108_A4 = CLBLM_L_X64Y108_SLICE_X96Y108_AQ;
  assign CLBLM_R_X63Y108_SLICE_X94Y108_A5 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X94Y108_A6 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X94Y108_AX = CLBLM_L_X64Y108_SLICE_X96Y108_AQ;
  assign CLBLM_R_X63Y108_SLICE_X94Y108_B1 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X94Y108_B2 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X94Y108_B3 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X94Y108_B4 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X94Y108_B5 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X94Y108_B6 = CLBLM_L_X64Y108_SLICE_X97Y108_AQ;
  assign CLBLM_R_X63Y108_SLICE_X94Y108_BX = CLBLM_L_X64Y108_SLICE_X97Y108_AQ;
  assign CLBLM_R_X63Y108_SLICE_X94Y108_C1 = CLBLM_R_X63Y110_SLICE_X94Y110_AQ;
  assign CLBLM_R_X63Y108_SLICE_X94Y108_C2 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X94Y108_C3 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X94Y108_C4 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X94Y108_C5 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X94Y108_C6 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X94Y108_CIN = CLBLM_R_X63Y107_SLICE_X94Y107_COUT;
  assign CLBLM_R_X63Y108_SLICE_X94Y108_CX = CLBLM_R_X63Y110_SLICE_X94Y110_AQ;
  assign CLBLM_R_X63Y108_SLICE_X94Y108_D1 = CLBLM_L_X64Y108_SLICE_X96Y108_BQ;
  assign CLBLM_R_X63Y108_SLICE_X94Y108_D2 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X94Y108_D3 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X94Y108_D4 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X94Y108_D5 = 1'b1;
  assign CLBLM_R_X63Y108_SLICE_X94Y108_D6 = 1'b1;
  assign CLBLM_R_X59Y99_SLICE_X89Y99_A3 = CLBLM_R_X59Y100_SLICE_X89Y100_DQ;
  assign CLBLM_R_X63Y108_SLICE_X94Y108_DX = CLBLM_L_X64Y108_SLICE_X96Y108_BQ;
  assign CLBLM_R_X59Y99_SLICE_X89Y99_A4 = CLBLM_L_X56Y99_SLICE_X84Y99_AQ;
  assign CLBLL_L_X54Y107_SLICE_X82Y107_A1 = CLBLL_L_X54Y106_SLICE_X83Y106_DO6;
  assign CLBLL_L_X54Y107_SLICE_X82Y107_A2 = CLBLM_L_X56Y101_SLICE_X85Y101_BQ;
  assign CLBLL_L_X54Y107_SLICE_X82Y107_A3 = 1'b1;
  assign CLBLL_L_X54Y107_SLICE_X82Y107_A4 = CLBLL_L_X54Y107_SLICE_X83Y107_AO5;
  assign CLBLL_L_X54Y107_SLICE_X82Y107_A5 = CLBLM_R_X53Y107_SLICE_X80Y107_BO6;
  assign CLBLL_L_X54Y107_SLICE_X82Y107_A6 = CLBLL_R_X57Y101_SLICE_X87Y101_DQ;
  assign CLBLM_R_X59Y99_SLICE_X89Y99_A6 = 1'b1;
  assign CLBLL_L_X54Y107_SLICE_X82Y107_AX = CLBLL_L_X54Y106_SLICE_X83Y106_DO6;
  assign CLBLL_L_X54Y107_SLICE_X82Y107_B1 = CLBLL_L_X54Y108_SLICE_X83Y108_AO5;
  assign CLBLL_L_X54Y107_SLICE_X82Y107_B2 = CLBLL_L_X54Y107_SLICE_X83Y107_DO6;
  assign CLBLL_L_X54Y107_SLICE_X82Y107_B3 = CLBLL_R_X57Y101_SLICE_X87Y101_AQ;
  assign CLBLL_L_X54Y107_SLICE_X82Y107_B4 = CLBLL_L_X52Y107_SLICE_X78Y107_BO6;
  assign CLBLL_L_X54Y107_SLICE_X82Y107_B5 = CLBLL_R_X57Y99_SLICE_X86Y99_BQ;
  assign CLBLL_L_X54Y107_SLICE_X82Y107_B6 = CLBLM_R_X53Y108_SLICE_X81Y108_A_XOR;
  assign CLBLL_L_X54Y107_SLICE_X82Y107_BX = CLBLL_L_X54Y107_SLICE_X83Y107_DO6;
  assign CLBLL_L_X54Y107_SLICE_X82Y107_C1 = CLBLL_L_X52Y106_SLICE_X78Y106_AO6;
  assign CLBLL_L_X54Y107_SLICE_X82Y107_C2 = CLBLL_L_X54Y107_SLICE_X83Y107_CO6;
  assign CLBLL_L_X54Y107_SLICE_X82Y107_C3 = CLBLM_R_X53Y108_SLICE_X81Y108_B_XOR;
  assign CLBLL_L_X54Y107_SLICE_X82Y107_C4 = CLBLL_R_X57Y99_SLICE_X86Y99_BQ;
  assign CLBLL_L_X54Y107_SLICE_X82Y107_C5 = CLBLM_L_X56Y101_SLICE_X85Y101_BQ;
  assign CLBLL_L_X54Y107_SLICE_X82Y107_C6 = CLBLL_L_X54Y108_SLICE_X83Y108_AO6;
  assign CLBLM_R_X59Y99_SLICE_X89Y99_B1 = 1'b1;
  assign CLBLL_L_X54Y107_SLICE_X82Y107_CIN = CLBLL_L_X54Y106_SLICE_X82Y106_COUT;
  assign CLBLM_R_X59Y99_SLICE_X89Y99_B2 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLL_L_X54Y107_SLICE_X82Y107_CX = CLBLL_L_X54Y107_SLICE_X83Y107_CO6;
  assign CLBLL_L_X54Y107_SLICE_X82Y107_D1 = CLBLL_R_X57Y101_SLICE_X87Y101_DQ;
  assign CLBLL_L_X54Y107_SLICE_X82Y107_D2 = CLBLL_R_X57Y99_SLICE_X86Y99_BQ;
  assign CLBLL_L_X54Y107_SLICE_X82Y107_D3 = CLBLL_L_X54Y107_SLICE_X83Y107_AO6;
  assign CLBLL_L_X54Y107_SLICE_X82Y107_D4 = CLBLL_R_X57Y100_SLICE_X87Y100_BQ;
  assign CLBLL_L_X54Y107_SLICE_X82Y107_D5 = CLBLL_R_X57Y99_SLICE_X86Y99_AQ;
  assign CLBLL_L_X54Y107_SLICE_X82Y107_D6 = CLBLM_R_X53Y108_SLICE_X81Y108_C_CY;
  assign CLBLM_R_X59Y99_SLICE_X89Y99_B3 = CLBLM_R_X59Y98_SLICE_X88Y98_BQ;
  assign CLBLM_R_X59Y99_SLICE_X89Y99_B4 = CLBLM_L_X56Y99_SLICE_X84Y99_AQ;
  assign CLBLL_L_X54Y107_SLICE_X82Y107_DX = CLBLL_L_X54Y107_SLICE_X83Y107_BO6;
  assign CLBLM_R_X59Y99_SLICE_X89Y99_B6 = CLBLM_L_X56Y99_SLICE_X84Y99_BQ;
  assign CLBLL_L_X54Y107_SLICE_X83Y107_A1 = CLBLM_R_X53Y108_SLICE_X81Y108_A_XOR;
  assign CLBLL_L_X54Y107_SLICE_X83Y107_A2 = CLBLL_R_X57Y101_SLICE_X87Y101_AQ;
  assign CLBLL_L_X54Y107_SLICE_X83Y107_A3 = CLBLL_R_X57Y99_SLICE_X86Y99_BQ;
  assign CLBLL_L_X54Y107_SLICE_X83Y107_A4 = CLBLM_L_X56Y101_SLICE_X85Y101_BQ;
  assign CLBLL_L_X54Y107_SLICE_X83Y107_A5 = CLBLM_R_X53Y108_SLICE_X81Y108_B_XOR;
  assign CLBLL_L_X54Y107_SLICE_X83Y107_A6 = 1'b1;
  assign CLBLL_L_X54Y107_SLICE_X83Y107_B1 = CLBLM_R_X53Y108_SLICE_X81Y108_B_XOR;
  assign CLBLL_L_X54Y107_SLICE_X83Y107_B2 = CLBLM_R_X53Y108_SLICE_X81Y108_C_CY;
  assign CLBLL_L_X54Y107_SLICE_X83Y107_B3 = CLBLL_L_X52Y106_SLICE_X78Y106_AO6;
  assign CLBLL_L_X54Y107_SLICE_X83Y107_B4 = CLBLL_R_X57Y99_SLICE_X86Y99_BQ;
  assign CLBLL_L_X54Y107_SLICE_X83Y107_B5 = CLBLM_L_X56Y101_SLICE_X85Y101_BQ;
  assign CLBLL_L_X54Y107_SLICE_X83Y107_B6 = CLBLL_R_X57Y100_SLICE_X87Y100_BQ;
  assign CLBLL_L_X54Y107_SLICE_X83Y107_C1 = CLBLM_R_X53Y108_SLICE_X81Y108_B_XOR;
  assign CLBLL_L_X54Y107_SLICE_X83Y107_C2 = CLBLL_R_X57Y101_SLICE_X87Y101_AQ;
  assign CLBLL_L_X54Y107_SLICE_X83Y107_C3 = CLBLM_L_X56Y101_SLICE_X85Y101_BQ;
  assign CLBLL_L_X54Y107_SLICE_X83Y107_C4 = CLBLL_R_X57Y99_SLICE_X86Y99_BQ;
  assign CLBLL_L_X54Y107_SLICE_X83Y107_C5 = CLBLM_R_X53Y108_SLICE_X81Y108_A_XOR;
  assign CLBLL_L_X54Y107_SLICE_X83Y107_C6 = CLBLL_L_X52Y107_SLICE_X78Y107_BO6;
  assign CLBLL_L_X54Y107_SLICE_X83Y107_D1 = CLBLL_R_X57Y101_SLICE_X87Y101_DQ;
  assign CLBLL_L_X54Y107_SLICE_X83Y107_D2 = CLBLL_R_X57Y101_SLICE_X87Y101_AQ;
  assign CLBLL_L_X54Y107_SLICE_X83Y107_D3 = CLBLM_L_X56Y101_SLICE_X85Y101_BQ;
  assign CLBLL_L_X54Y107_SLICE_X83Y107_D4 = CLBLM_R_X53Y107_SLICE_X80Y107_BO6;
  assign CLBLL_L_X54Y107_SLICE_X83Y107_D5 = CLBLM_R_X53Y108_SLICE_X81Y108_A_XOR;
  assign CLBLL_L_X54Y107_SLICE_X83Y107_D6 = CLBLL_R_X57Y99_SLICE_X86Y99_BQ;
  assign CLBLM_R_X59Y99_SLICE_X89Y99_CE = CLBLL_R_X57Y99_SLICE_X87Y99_BO6;
  assign CLBLM_R_X59Y99_SLICE_X89Y99_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X59Y99_SLICE_X89Y99_D6 = 1'b1;
  assign CLBLM_R_X59Y99_SLICE_X89Y99_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X63Y109_SLICE_X95Y109_A1 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X95Y109_A2 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X95Y109_A3 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X95Y109_A4 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X95Y109_A5 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X95Y109_A6 = CLBLM_L_X62Y103_SLICE_X93Y103_AQ;
  assign CLBLM_R_X63Y109_SLICE_X95Y109_AX = 1'b0;
  assign CLBLM_R_X63Y109_SLICE_X95Y109_B1 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X95Y109_B2 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X95Y109_B3 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X95Y109_B4 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X95Y109_B5 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X95Y109_B6 = CLBLM_R_X63Y105_SLICE_X94Y105_AQ;
  assign LIOB33_X0Y137_IOB_X0Y137_O = CLBLM_R_X49Y109_SLICE_X74Y109_BQ;
  assign LIOB33_X0Y137_IOB_X0Y138_O = CLBLM_R_X49Y111_SLICE_X74Y111_CQ;
  assign CLBLM_R_X63Y109_SLICE_X95Y109_BX = 1'b0;
  assign CLBLM_R_X63Y109_SLICE_X95Y109_C1 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X95Y109_C2 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X95Y109_C3 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X95Y109_C4 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X95Y109_C5 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X95Y109_C6 = CLBLM_L_X64Y109_SLICE_X96Y109_A5Q;
  assign CLBLM_R_X63Y109_SLICE_X95Y109_CIN = CLBLM_R_X63Y108_SLICE_X95Y108_COUT;
  assign CLBLM_R_X63Y109_SLICE_X95Y109_CX = 1'b0;
  assign CLBLM_R_X63Y109_SLICE_X95Y109_D1 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X95Y109_D2 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X95Y109_D3 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X95Y109_D4 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X95Y109_D5 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X95Y109_D6 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X95Y109_DX = 1'b0;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_D1 = CLBLM_L_X62Y110_SLICE_X92Y110_AQ;
  assign CLBLM_R_X63Y109_SLICE_X94Y109_A1 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X94Y109_A2 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X94Y109_A3 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X94Y109_A4 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X94Y109_A5 = CLBLM_L_X64Y109_SLICE_X96Y109_AQ;
  assign CLBLM_R_X63Y109_SLICE_X94Y109_A6 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X94Y109_AX = CLBLM_L_X64Y109_SLICE_X96Y109_AQ;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_T1 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X94Y109_B1 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X94Y109_B2 = CLBLM_L_X62Y103_SLICE_X93Y103_AQ;
  assign CLBLM_R_X63Y109_SLICE_X94Y109_B3 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X94Y109_B4 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X94Y109_B5 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X94Y109_B6 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X94Y109_BX = CLBLM_L_X62Y103_SLICE_X93Y103_AQ;
  assign CLBLM_R_X63Y109_SLICE_X94Y109_C1 = CLBLM_R_X63Y105_SLICE_X94Y105_AQ;
  assign CLBLM_R_X63Y109_SLICE_X94Y109_C2 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X94Y109_C3 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X94Y109_C4 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X94Y109_C5 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X94Y109_C6 = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_D1 = CLBLM_L_X62Y106_SLICE_X93Y106_AQ;
  assign CLBLM_R_X63Y109_SLICE_X94Y109_CIN = CLBLM_R_X63Y108_SLICE_X94Y108_COUT;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_T1 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X94Y109_CX = CLBLM_R_X63Y105_SLICE_X94Y105_AQ;
  assign CLBLM_R_X63Y109_SLICE_X94Y109_D1 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X94Y109_D2 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X94Y109_D3 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X94Y109_D4 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X94Y109_D5 = 1'b1;
  assign CLBLM_R_X63Y109_SLICE_X94Y109_D6 = CLBLM_L_X64Y109_SLICE_X96Y109_A5Q;
  assign CLBLM_R_X63Y109_SLICE_X94Y109_DX = 1'b0;
  assign CLBLL_L_X54Y108_SLICE_X82Y108_A1 = 1'b1;
  assign CLBLL_L_X54Y108_SLICE_X82Y108_A2 = 1'b1;
  assign CLBLL_L_X54Y108_SLICE_X82Y108_A3 = CLBLL_R_X57Y99_SLICE_X86Y99_AQ;
  assign CLBLL_L_X54Y108_SLICE_X82Y108_A4 = CLBLM_R_X53Y108_SLICE_X81Y108_C_CY;
  assign CLBLL_L_X54Y108_SLICE_X82Y108_A5 = CLBLL_R_X57Y99_SLICE_X86Y99_BQ;
  assign CLBLL_L_X54Y108_SLICE_X82Y108_A6 = CLBLL_R_X57Y100_SLICE_X87Y100_BQ;
  assign CLBLL_L_X54Y108_SLICE_X82Y108_AX = 1'b0;
  assign CLBLL_L_X54Y108_SLICE_X82Y108_B1 = 1'b1;
  assign CLBLL_L_X54Y108_SLICE_X82Y108_B2 = 1'b1;
  assign CLBLL_L_X54Y108_SLICE_X82Y108_B3 = 1'b1;
  assign CLBLL_L_X54Y108_SLICE_X82Y108_B4 = 1'b1;
  assign CLBLL_L_X54Y108_SLICE_X82Y108_B5 = 1'b1;
  assign CLBLL_L_X54Y108_SLICE_X82Y108_B6 = 1'b1;
  assign CLBLL_L_X54Y108_SLICE_X82Y108_BX = 1'b0;
  assign CLBLL_L_X54Y108_SLICE_X82Y108_C1 = 1'b1;
  assign CLBLL_L_X54Y108_SLICE_X82Y108_C2 = 1'b1;
  assign CLBLL_L_X54Y108_SLICE_X82Y108_C3 = 1'b1;
  assign CLBLL_L_X54Y108_SLICE_X82Y108_C4 = 1'b1;
  assign CLBLL_L_X54Y108_SLICE_X82Y108_C5 = 1'b1;
  assign CLBLL_L_X54Y108_SLICE_X82Y108_C6 = 1'b1;
  assign CLBLL_L_X54Y108_SLICE_X82Y108_CIN = CLBLL_L_X54Y107_SLICE_X82Y107_COUT;
  assign CLBLL_L_X54Y108_SLICE_X82Y108_CX = 1'b0;
  assign CLBLL_L_X54Y108_SLICE_X82Y108_D1 = 1'b1;
  assign CLBLL_L_X54Y108_SLICE_X82Y108_D2 = 1'b1;
  assign CLBLL_L_X54Y108_SLICE_X82Y108_D3 = 1'b1;
  assign CLBLL_L_X54Y108_SLICE_X82Y108_D4 = 1'b1;
  assign CLBLL_L_X54Y108_SLICE_X82Y108_D5 = 1'b1;
  assign CLBLL_L_X54Y108_SLICE_X82Y108_D6 = 1'b1;
  assign CLBLL_L_X54Y108_SLICE_X82Y108_DX = 1'b0;
  assign CLBLL_L_X54Y108_SLICE_X83Y108_A1 = CLBLL_R_X57Y99_SLICE_X86Y99_BQ;
  assign CLBLL_L_X54Y108_SLICE_X83Y108_A2 = CLBLM_R_X53Y108_SLICE_X81Y108_C_CY;
  assign CLBLL_L_X54Y108_SLICE_X83Y108_A3 = CLBLM_R_X53Y108_SLICE_X81Y108_B_XOR;
  assign CLBLL_L_X54Y108_SLICE_X83Y108_A4 = CLBLM_L_X56Y101_SLICE_X85Y101_BQ;
  assign CLBLL_L_X54Y108_SLICE_X83Y108_A5 = CLBLL_R_X57Y100_SLICE_X87Y100_BQ;
  assign CLBLL_L_X54Y108_SLICE_X83Y108_A6 = 1'b1;
  assign CLBLL_L_X54Y108_SLICE_X83Y108_B1 = 1'b1;
  assign CLBLL_L_X54Y108_SLICE_X83Y108_B2 = 1'b1;
  assign CLBLL_L_X54Y108_SLICE_X83Y108_B3 = 1'b1;
  assign CLBLL_L_X54Y108_SLICE_X83Y108_B4 = 1'b1;
  assign CLBLL_L_X54Y108_SLICE_X83Y108_B5 = 1'b1;
  assign CLBLL_L_X54Y108_SLICE_X83Y108_B6 = 1'b1;
  assign CLBLL_L_X54Y108_SLICE_X83Y108_C1 = 1'b1;
  assign CLBLL_L_X54Y108_SLICE_X83Y108_C2 = 1'b1;
  assign CLBLL_L_X54Y108_SLICE_X83Y108_C3 = 1'b1;
  assign CLBLL_L_X54Y108_SLICE_X83Y108_C4 = 1'b1;
  assign CLBLL_L_X54Y108_SLICE_X83Y108_C5 = 1'b1;
  assign CLBLL_L_X54Y108_SLICE_X83Y108_C6 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X95Y94_A2 = 1'b1;
  assign CLBLL_L_X54Y108_SLICE_X83Y108_D1 = 1'b1;
  assign CLBLL_L_X54Y108_SLICE_X83Y108_D2 = 1'b1;
  assign CLBLL_L_X54Y108_SLICE_X83Y108_D3 = 1'b1;
  assign CLBLL_L_X54Y108_SLICE_X83Y108_D4 = 1'b1;
  assign CLBLL_L_X54Y108_SLICE_X83Y108_D5 = 1'b1;
  assign CLBLL_L_X54Y108_SLICE_X83Y108_D6 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X95Y94_A6 = CLBLM_L_X64Y95_SLICE_X96Y95_AO5;
  assign CLBLM_R_X63Y94_SLICE_X95Y94_B1 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X95Y94_B2 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X95Y94_B3 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X95Y94_B4 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X95Y94_B5 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X95Y94_B6 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X95Y94_C1 = 1'b1;
  assign LIOB33_X0Y139_IOB_X0Y140_O = CLBLM_L_X50Y104_SLICE_X76Y104_AQ;
  assign LIOB33_X0Y139_IOB_X0Y139_O = CLBLM_R_X49Y109_SLICE_X74Y109_CQ;
  assign CLBLM_R_X63Y94_SLICE_X95Y94_C2 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X95Y94_C3 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X95Y94_C4 = 1'b1;
  assign CLBLM_R_X63Y110_SLICE_X95Y110_A1 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X95Y94_C5 = 1'b1;
  assign CLBLM_R_X63Y110_SLICE_X95Y110_A2 = 1'b1;
  assign CLBLM_R_X63Y110_SLICE_X95Y110_A3 = 1'b1;
  assign CLBLM_R_X63Y110_SLICE_X95Y110_A4 = 1'b1;
  assign CLBLM_R_X63Y110_SLICE_X95Y110_A5 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X95Y94_C6 = 1'b1;
  assign CLBLM_R_X63Y110_SLICE_X95Y110_A6 = 1'b1;
  assign CLBLM_R_X63Y110_SLICE_X95Y110_B1 = 1'b1;
  assign CLBLM_R_X63Y110_SLICE_X95Y110_B2 = 1'b1;
  assign CLBLM_R_X63Y110_SLICE_X95Y110_B3 = 1'b1;
  assign CLBLM_R_X63Y110_SLICE_X95Y110_B4 = 1'b1;
  assign CLBLM_R_X63Y110_SLICE_X95Y110_B5 = 1'b1;
  assign CLBLM_R_X63Y110_SLICE_X95Y110_B6 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X95Y94_CE = CLBLM_L_X62Y99_SLICE_X93Y99_CO6;
  assign CLBLM_R_X63Y110_SLICE_X95Y110_C1 = 1'b1;
  assign CLBLM_R_X63Y110_SLICE_X95Y110_C2 = 1'b1;
  assign CLBLM_R_X63Y110_SLICE_X95Y110_C3 = 1'b1;
  assign CLBLM_R_X63Y110_SLICE_X95Y110_C4 = 1'b1;
  assign CLBLM_R_X63Y110_SLICE_X95Y110_C5 = 1'b1;
  assign CLBLM_R_X63Y110_SLICE_X95Y110_C6 = 1'b1;
  assign CLBLM_R_X53Y98_SLICE_X81Y98_A1 = CLBLL_L_X52Y99_SLICE_X78Y99_AO6;
  assign CLBLM_R_X53Y98_SLICE_X81Y98_A2 = CLBLM_R_X53Y99_SLICE_X80Y99_AO5;
  assign CLBLM_R_X53Y98_SLICE_X81Y98_A3 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLM_R_X53Y98_SLICE_X81Y98_A4 = CLBLM_R_X53Y98_SLICE_X81Y98_BO6;
  assign CLBLM_R_X53Y98_SLICE_X81Y98_A5 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLM_R_X53Y98_SLICE_X81Y98_A6 = CLBLM_R_X53Y98_SLICE_X81Y98_CO6;
  assign CLBLM_R_X53Y98_SLICE_X81Y98_B1 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLM_R_X63Y110_SLICE_X95Y110_D1 = 1'b1;
  assign CLBLM_R_X63Y110_SLICE_X95Y110_D2 = 1'b1;
  assign CLBLM_R_X63Y110_SLICE_X95Y110_D3 = 1'b1;
  assign CLBLM_R_X63Y110_SLICE_X95Y110_D4 = 1'b1;
  assign CLBLM_R_X63Y110_SLICE_X95Y110_D5 = 1'b1;
  assign CLBLM_R_X63Y110_SLICE_X95Y110_D6 = 1'b1;
  assign CLBLM_R_X53Y98_SLICE_X81Y98_B2 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign CLBLM_R_X53Y98_SLICE_X81Y98_B3 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLM_R_X53Y98_SLICE_X81Y98_B4 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLM_R_X53Y98_SLICE_X81Y98_B5 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLM_R_X53Y98_SLICE_X81Y98_B6 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLM_R_X63Y110_SLICE_X94Y110_A1 = CLBLM_R_X63Y108_SLICE_X95Y108_B_XOR;
  assign CLBLM_R_X63Y110_SLICE_X94Y110_A2 = CLBLM_L_X62Y105_SLICE_X93Y105_AO6;
  assign CLBLM_R_X63Y110_SLICE_X94Y110_A3 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X63Y110_SLICE_X94Y110_A4 = CLBLM_R_X63Y110_SLICE_X94Y110_BO6;
  assign CLBLM_R_X63Y110_SLICE_X94Y110_A5 = CLBLM_R_X63Y108_SLICE_X94Y108_C_XOR;
  assign CLBLM_R_X63Y110_SLICE_X94Y110_A6 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X53Y98_SLICE_X81Y98_C2 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLM_R_X53Y98_SLICE_X81Y98_C3 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLM_R_X53Y98_SLICE_X81Y98_C4 = CLBLM_R_X53Y100_SLICE_X81Y100_AO5;
  assign CLBLM_R_X53Y98_SLICE_X81Y98_C6 = CLBLM_R_X49Y107_SLICE_X75Y107_DQ;
  assign CLBLM_R_X63Y110_SLICE_X94Y110_B1 = CLBLM_R_X63Y108_SLICE_X95Y108_B_XOR;
  assign CLBLM_R_X63Y110_SLICE_X94Y110_B2 = CLBLM_L_X50Y107_SLICE_X76Y107_BQ;
  assign CLBLM_R_X63Y110_SLICE_X94Y110_B3 = CLBLM_L_X62Y112_SLICE_X92Y112_AQ;
  assign CLBLM_R_X63Y110_SLICE_X94Y110_B4 = CLBLM_R_X63Y110_SLICE_X94Y110_AQ;
  assign CLBLM_R_X63Y110_SLICE_X94Y110_B5 = CLBLM_L_X62Y105_SLICE_X92Y105_BO5;
  assign CLBLM_R_X63Y110_SLICE_X94Y110_B6 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X53Y98_SLICE_X81Y98_D1 = 1'b1;
  assign CLBLM_R_X53Y98_SLICE_X81Y98_D2 = 1'b1;
  assign CLBLM_R_X53Y98_SLICE_X81Y98_D3 = 1'b1;
  assign CLBLM_R_X63Y110_SLICE_X94Y110_C1 = CLBLM_L_X62Y105_SLICE_X92Y105_BO5;
  assign CLBLM_R_X63Y110_SLICE_X94Y110_C2 = CLBLM_L_X62Y105_SLICE_X93Y105_AO6;
  assign CLBLM_R_X63Y110_SLICE_X94Y110_C3 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X63Y110_SLICE_X94Y110_C4 = CLBLM_R_X63Y109_SLICE_X95Y109_A_XOR;
  assign CLBLM_R_X63Y110_SLICE_X94Y110_C5 = CLBLM_R_X63Y109_SLICE_X94Y109_B_XOR;
  assign CLBLM_R_X63Y110_SLICE_X94Y110_C6 = CLBLM_L_X62Y103_SLICE_X93Y103_AQ;
  assign CLBLM_R_X63Y110_SLICE_X94Y110_CE = CLBLM_R_X63Y100_SLICE_X94Y100_CO6;
  assign CLBLM_R_X53Y98_SLICE_X80Y98_A1 = 1'b1;
  assign CLBLM_R_X53Y98_SLICE_X80Y98_A2 = 1'b1;
  assign CLBLM_R_X63Y110_SLICE_X94Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X53Y98_SLICE_X80Y98_A3 = 1'b1;
  assign CLBLM_R_X53Y98_SLICE_X80Y98_A4 = 1'b1;
  assign CLBLM_R_X53Y98_SLICE_X80Y98_A5 = 1'b1;
  assign CLBLM_R_X53Y98_SLICE_X80Y98_A6 = 1'b1;
  assign CLBLM_R_X63Y110_SLICE_X94Y110_D1 = 1'b1;
  assign CLBLM_R_X63Y110_SLICE_X94Y110_D2 = 1'b1;
  assign CLBLM_R_X63Y110_SLICE_X94Y110_D3 = 1'b1;
  assign CLBLM_R_X63Y110_SLICE_X94Y110_D4 = 1'b1;
  assign CLBLM_R_X63Y110_SLICE_X94Y110_D5 = 1'b1;
  assign CLBLM_R_X63Y110_SLICE_X94Y110_D6 = 1'b1;
  assign CLBLM_R_X53Y98_SLICE_X80Y98_B1 = 1'b1;
  assign CLBLM_R_X53Y98_SLICE_X80Y98_B2 = 1'b1;
  assign CLBLM_R_X53Y98_SLICE_X80Y98_B3 = 1'b1;
  assign CLBLM_R_X63Y110_SLICE_X94Y110_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X53Y98_SLICE_X80Y98_C3 = 1'b1;
  assign CLBLM_R_X53Y98_SLICE_X80Y98_C4 = 1'b1;
  assign CLBLM_R_X53Y98_SLICE_X80Y98_C5 = 1'b1;
  assign CLBLM_R_X53Y98_SLICE_X80Y98_C1 = 1'b1;
  assign CLBLM_R_X53Y98_SLICE_X80Y98_C2 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X82Y109_A1 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X82Y109_A2 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X82Y109_A3 = CLBLL_L_X54Y109_SLICE_X82Y109_AQ;
  assign CLBLL_L_X54Y109_SLICE_X82Y109_A4 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X82Y109_A5 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X82Y109_A6 = 1'b1;
  assign CLBLM_R_X53Y98_SLICE_X80Y98_D1 = 1'b1;
  assign CLBLM_R_X53Y98_SLICE_X80Y98_D2 = 1'b1;
  assign CLBLM_R_X53Y98_SLICE_X80Y98_D3 = 1'b1;
  assign CLBLM_R_X53Y98_SLICE_X80Y98_D4 = 1'b1;
  assign CLBLM_R_X53Y98_SLICE_X80Y98_D5 = 1'b1;
  assign CLBLM_R_X53Y98_SLICE_X80Y98_D6 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X82Y109_B1 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X82Y109_B2 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X82Y109_B3 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X82Y109_B4 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X82Y109_B5 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X82Y109_B6 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X82Y109_C1 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X82Y109_C2 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X82Y109_C3 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X82Y109_C4 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X82Y109_C5 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X82Y109_C6 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X82Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_T1 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X82Y109_D1 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X82Y109_D2 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X82Y109_D3 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X82Y109_D4 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X82Y109_D5 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X82Y109_D6 = 1'b1;
  assign CLBLM_R_X63Y94_SLICE_X94Y94_A4 = CLBLM_R_X63Y99_SLICE_X95Y99_A5Q;
  assign CLBLM_R_X63Y94_SLICE_X94Y94_A5 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X82Y109_SR = CLBLM_R_X15Y122_SLICE_X20Y122_AO6;
  assign CLBLL_L_X54Y109_SLICE_X83Y109_A1 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X83Y109_A2 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X83Y109_A3 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X83Y109_A4 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X83Y109_A5 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X83Y109_A6 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X83Y109_B1 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X83Y109_B2 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X83Y109_B3 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X83Y109_B4 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X83Y109_B5 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X83Y109_B6 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X83Y109_C1 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X83Y109_C2 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X83Y109_C3 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X83Y109_C4 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X83Y109_C5 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X83Y109_C6 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X83Y109_D1 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X83Y109_D2 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X83Y109_D3 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X83Y109_D4 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X83Y109_D5 = 1'b1;
  assign CLBLL_L_X54Y109_SLICE_X83Y109_D6 = 1'b1;
  assign LIOB33_X0Y141_IOB_X0Y142_O = CLBLM_R_X49Y105_SLICE_X75Y105_CQ;
  assign LIOB33_X0Y141_IOB_X0Y141_O = CLBLM_L_X50Y105_SLICE_X77Y105_AQ;
  assign CLBLM_R_X53Y99_SLICE_X81Y99_A1 = CLBLM_R_X53Y99_SLICE_X80Y99_AO5;
  assign CLBLM_R_X53Y99_SLICE_X81Y99_A2 = 1'b1;
  assign CLBLM_R_X53Y99_SLICE_X81Y99_A3 = CLBLM_R_X49Y107_SLICE_X75Y107_DQ;
  assign CLBLM_R_X53Y99_SLICE_X81Y99_A4 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLM_R_X53Y99_SLICE_X81Y99_A5 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLM_R_X53Y99_SLICE_X81Y99_A6 = 1'b1;
  assign CLBLM_R_X53Y99_SLICE_X81Y99_AX = CLBLM_R_X53Y99_SLICE_X81Y99_BQ;
  assign CLBLM_R_X53Y99_SLICE_X81Y99_B1 = CLBLM_R_X53Y99_SLICE_X80Y99_AO5;
  assign CLBLM_R_X53Y99_SLICE_X81Y99_B2 = CLBLL_L_X52Y99_SLICE_X79Y99_AO6;
  assign CLBLM_R_X53Y99_SLICE_X81Y99_B3 = CLBLM_R_X49Y107_SLICE_X75Y107_DQ;
  assign CLBLM_R_X53Y99_SLICE_X81Y99_B4 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLM_R_X53Y99_SLICE_X81Y99_B5 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLM_R_X53Y99_SLICE_X81Y99_B6 = CLBLL_L_X54Y100_SLICE_X82Y100_AO5;
  assign CLBLM_R_X53Y99_SLICE_X81Y99_C1 = CLBLM_R_X53Y99_SLICE_X81Y99_AO6;
  assign CLBLM_R_X53Y99_SLICE_X81Y99_C2 = CLBLL_L_X52Y99_SLICE_X78Y99_AO6;
  assign CLBLM_R_X53Y99_SLICE_X81Y99_C3 = CLBLM_R_X53Y99_SLICE_X80Y99_DO6;
  assign CLBLM_R_X53Y99_SLICE_X81Y99_C4 = CLBLM_R_X53Y99_SLICE_X81Y99_AO5;
  assign CLBLM_R_X53Y99_SLICE_X81Y99_C5 = CLBLM_R_X53Y99_SLICE_X81Y99_DO6;
  assign CLBLM_R_X53Y99_SLICE_X81Y99_C6 = CLBLM_R_X53Y99_SLICE_X80Y99_BO5;
  assign CLBLM_R_X53Y99_SLICE_X81Y99_CE = CLBLM_L_X60Y98_SLICE_X91Y98_DQ;
  assign CLBLM_R_X53Y99_SLICE_X81Y99_CLK = CLK_HROW_BOT_R_X139Y78_BUFHCE_X0Y20_O;
  assign CLBLM_R_X53Y99_SLICE_X81Y99_D1 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLM_R_X53Y99_SLICE_X81Y99_D2 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLM_R_X53Y99_SLICE_X81Y99_D3 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLM_R_X53Y99_SLICE_X81Y99_D4 = CLBLL_L_X54Y99_SLICE_X83Y99_BO5;
  assign CLBLM_R_X53Y99_SLICE_X81Y99_D5 = CLBLM_R_X49Y108_SLICE_X75Y108_DQ;
  assign CLBLM_R_X53Y99_SLICE_X81Y99_D6 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign CLBLM_R_X53Y99_SLICE_X81Y99_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X53Y99_SLICE_X80Y99_A1 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLM_R_X53Y99_SLICE_X80Y99_A2 = 1'b1;
  assign CLBLM_R_X53Y99_SLICE_X80Y99_A3 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLM_R_X53Y99_SLICE_X80Y99_A4 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign CLBLM_R_X53Y99_SLICE_X80Y99_A5 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLM_R_X53Y99_SLICE_X80Y99_A6 = 1'b1;
  assign CLBLM_R_X53Y99_SLICE_X80Y99_B1 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLM_R_X53Y99_SLICE_X80Y99_B2 = CLBLM_R_X49Y108_SLICE_X75Y108_DQ;
  assign CLBLM_R_X53Y99_SLICE_X80Y99_B3 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLM_R_X53Y99_SLICE_X80Y99_B4 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign CLBLM_R_X53Y99_SLICE_X80Y99_B5 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLM_R_X53Y99_SLICE_X80Y99_B6 = 1'b1;
  assign CLBLM_R_X53Y99_SLICE_X80Y99_C1 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLM_R_X53Y99_SLICE_X80Y99_C2 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLM_R_X53Y99_SLICE_X80Y99_C3 = CLBLM_R_X53Y100_SLICE_X81Y100_DO6;
  assign CLBLM_R_X53Y99_SLICE_X80Y99_C4 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLM_R_X53Y99_SLICE_X80Y99_C5 = CLBLM_L_X56Y97_SLICE_X84Y97_AO6;
  assign CLBLM_R_X53Y99_SLICE_X80Y99_C6 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign CLBLM_R_X53Y99_SLICE_X80Y99_D1 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLM_R_X53Y99_SLICE_X80Y99_D2 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLM_R_X53Y99_SLICE_X80Y99_D3 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLM_R_X53Y99_SLICE_X80Y99_D4 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLM_R_X53Y99_SLICE_X80Y99_D5 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLM_R_X53Y99_SLICE_X80Y99_D6 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_D1 = CLBLM_L_X60Y111_SLICE_X91Y111_BQ;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_T1 = 1'b1;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_D1 = CLBLM_L_X62Y108_SLICE_X93Y108_AQ;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_T1 = 1'b1;
  assign CLBLL_L_X52Y99_SLICE_X78Y99_A1 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLL_L_X52Y99_SLICE_X78Y99_A2 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLL_L_X52Y99_SLICE_X78Y99_A3 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign CLBLL_L_X52Y99_SLICE_X78Y99_A4 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLL_L_X52Y99_SLICE_X78Y99_A5 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLL_L_X52Y99_SLICE_X78Y99_A6 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLL_L_X52Y99_SLICE_X78Y99_B1 = 1'b1;
  assign CLBLL_L_X52Y99_SLICE_X78Y99_B2 = 1'b1;
  assign CLBLL_L_X52Y99_SLICE_X78Y99_B3 = 1'b1;
  assign CLBLL_L_X52Y99_SLICE_X78Y99_B4 = 1'b1;
  assign CLBLL_L_X52Y99_SLICE_X78Y99_B5 = 1'b1;
  assign CLBLL_L_X52Y99_SLICE_X78Y99_B6 = 1'b1;
  assign LIOB33_X0Y143_IOB_X0Y143_O = CLBLM_R_X49Y106_SLICE_X74Y106_AQ;
  assign CLBLL_L_X52Y99_SLICE_X78Y99_C1 = 1'b1;
  assign CLBLL_L_X52Y99_SLICE_X78Y99_C2 = 1'b1;
  assign CLBLL_L_X52Y99_SLICE_X78Y99_C3 = 1'b1;
  assign CLBLL_L_X52Y99_SLICE_X78Y99_C4 = 1'b1;
  assign CLBLL_L_X52Y99_SLICE_X78Y99_C5 = 1'b1;
  assign CLBLL_L_X52Y99_SLICE_X78Y99_C6 = 1'b1;
  assign CLBLL_L_X52Y99_SLICE_X78Y99_D1 = 1'b1;
  assign CLBLL_L_X52Y99_SLICE_X78Y99_D2 = 1'b1;
  assign CLBLL_L_X52Y99_SLICE_X78Y99_D3 = 1'b1;
  assign CLBLL_L_X52Y99_SLICE_X78Y99_D4 = 1'b1;
  assign CLBLL_L_X52Y99_SLICE_X78Y99_D5 = 1'b1;
  assign CLBLL_L_X52Y99_SLICE_X78Y99_D6 = 1'b1;
  assign CLBLL_L_X52Y99_SLICE_X79Y99_A1 = CLBLL_L_X52Y99_SLICE_X79Y99_DO6;
  assign CLBLL_L_X52Y99_SLICE_X79Y99_A2 = CLBLM_R_X53Y99_SLICE_X80Y99_AO5;
  assign CLBLL_L_X52Y99_SLICE_X79Y99_A3 = CLBLM_L_X56Y97_SLICE_X84Y97_AO6;
  assign CLBLL_L_X52Y99_SLICE_X79Y99_A4 = CLBLL_L_X52Y99_SLICE_X79Y99_BO6;
  assign CLBLL_L_X52Y99_SLICE_X79Y99_A5 = CLBLL_L_X52Y101_SLICE_X79Y101_AO6;
  assign CLBLL_L_X52Y99_SLICE_X79Y99_A6 = CLBLL_L_X52Y99_SLICE_X79Y99_CO6;
  assign CLBLL_L_X52Y99_SLICE_X79Y99_B1 = CLBLM_R_X49Y108_SLICE_X75Y108_DQ;
  assign CLBLL_L_X52Y99_SLICE_X79Y99_B2 = CLBLM_R_X53Y99_SLICE_X80Y99_AO6;
  assign CLBLL_L_X52Y99_SLICE_X79Y99_B3 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLL_L_X52Y99_SLICE_X79Y99_B4 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLL_L_X52Y99_SLICE_X79Y99_B5 = CLBLM_R_X49Y107_SLICE_X75Y107_DQ;
  assign CLBLL_L_X52Y99_SLICE_X79Y99_B6 = CLBLM_L_X56Y97_SLICE_X84Y97_CO5;
  assign CLBLL_L_X52Y99_SLICE_X79Y99_C1 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLL_L_X52Y99_SLICE_X79Y99_C2 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLL_L_X52Y99_SLICE_X79Y99_C3 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLL_L_X52Y99_SLICE_X79Y99_C4 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLL_L_X52Y99_SLICE_X79Y99_C5 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign CLBLL_L_X52Y99_SLICE_X79Y99_C6 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLL_L_X52Y99_SLICE_X79Y99_D1 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLL_L_X52Y99_SLICE_X79Y99_D2 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLL_L_X52Y99_SLICE_X79Y99_D3 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLL_L_X52Y99_SLICE_X79Y99_D4 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign CLBLL_L_X52Y99_SLICE_X79Y99_D5 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLL_L_X52Y99_SLICE_X79Y99_D6 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLM_R_X53Y100_SLICE_X81Y100_A1 = CLBLL_L_X54Y100_SLICE_X82Y100_AO5;
  assign CLBLM_R_X53Y100_SLICE_X81Y100_A2 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLM_R_X53Y100_SLICE_X81Y100_A3 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLM_R_X53Y100_SLICE_X81Y100_A4 = CLBLM_R_X53Y100_SLICE_X81Y100_BO6;
  assign CLBLM_R_X53Y100_SLICE_X81Y100_A5 = CLBLL_L_X54Y99_SLICE_X82Y99_BO6;
  assign CLBLM_R_X53Y100_SLICE_X81Y100_A6 = 1'b1;
  assign CLBLM_R_X53Y100_SLICE_X81Y100_B1 = CLBLM_R_X53Y100_SLICE_X81Y100_AO5;
  assign CLBLM_R_X53Y100_SLICE_X81Y100_B2 = CLBLM_R_X53Y99_SLICE_X80Y99_BO6;
  assign CLBLM_R_X53Y100_SLICE_X81Y100_B3 = CLBLM_R_X49Y107_SLICE_X75Y107_DQ;
  assign CLBLM_R_X53Y100_SLICE_X81Y100_B4 = CLBLL_R_X57Y102_SLICE_X86Y102_AO6;
  assign CLBLM_R_X53Y100_SLICE_X81Y100_B5 = CLBLM_L_X56Y99_SLICE_X84Y99_CO6;
  assign CLBLM_R_X53Y100_SLICE_X81Y100_B6 = CLBLM_R_X53Y100_SLICE_X81Y100_CO6;
  assign CLBLM_R_X53Y100_SLICE_X81Y100_C1 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLM_R_X53Y100_SLICE_X81Y100_C2 = CLBLM_R_X49Y107_SLICE_X75Y107_DQ;
  assign CLBLM_R_X53Y100_SLICE_X81Y100_C3 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLM_R_X53Y100_SLICE_X81Y100_C4 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLM_R_X53Y100_SLICE_X81Y100_C5 = CLBLL_L_X54Y99_SLICE_X83Y99_BO5;
  assign CLBLM_R_X53Y100_SLICE_X81Y100_C6 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign CLBLM_R_X53Y100_SLICE_X81Y100_CE = CLBLM_L_X60Y98_SLICE_X91Y98_DQ;
  assign CLBLM_R_X53Y100_SLICE_X81Y100_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X53Y100_SLICE_X81Y100_D1 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLM_R_X53Y100_SLICE_X81Y100_D2 = CLBLM_L_X56Y100_SLICE_X85Y100_AO5;
  assign CLBLM_R_X53Y100_SLICE_X81Y100_D3 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLM_R_X53Y100_SLICE_X81Y100_D4 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLM_R_X53Y100_SLICE_X81Y100_D5 = CLBLM_R_X53Y99_SLICE_X81Y99_AO5;
  assign CLBLM_R_X53Y100_SLICE_X81Y100_D6 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign CLBLM_R_X53Y100_SLICE_X81Y100_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X53Y100_SLICE_X80Y100_A1 = CLBLM_R_X53Y100_SLICE_X80Y100_DO6;
  assign CLBLM_R_X53Y100_SLICE_X80Y100_A2 = CLBLM_R_X53Y99_SLICE_X80Y99_CO6;
  assign CLBLM_R_X53Y100_SLICE_X80Y100_A3 = CLBLM_R_X49Y107_SLICE_X75Y107_DQ;
  assign CLBLM_R_X53Y100_SLICE_X80Y100_A4 = CLBLM_R_X53Y100_SLICE_X80Y100_BO6;
  assign CLBLM_R_X53Y100_SLICE_X80Y100_A5 = CLBLM_R_X53Y100_SLICE_X80Y100_CO6;
  assign CLBLM_R_X53Y100_SLICE_X80Y100_A6 = 1'b1;
  assign CLBLM_R_X53Y100_SLICE_X80Y100_B1 = CLBLM_R_X49Y108_SLICE_X75Y108_DQ;
  assign CLBLM_R_X53Y100_SLICE_X80Y100_B2 = CLBLM_R_X49Y107_SLICE_X75Y107_DQ;
  assign CLBLM_R_X53Y100_SLICE_X80Y100_B3 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLM_R_X53Y100_SLICE_X80Y100_B4 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLM_R_X53Y100_SLICE_X80Y100_B5 = CLBLM_L_X56Y97_SLICE_X84Y97_CO5;
  assign CLBLM_R_X53Y100_SLICE_X80Y100_B6 = 1'b1;
  assign CLBLM_R_X53Y100_SLICE_X80Y100_C1 = CLBLM_L_X56Y99_SLICE_X84Y99_CO6;
  assign CLBLM_R_X53Y100_SLICE_X80Y100_C2 = CLBLL_R_X57Y102_SLICE_X86Y102_AO6;
  assign CLBLM_R_X53Y100_SLICE_X80Y100_C3 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLM_R_X53Y100_SLICE_X80Y100_C4 = CLBLM_R_X53Y99_SLICE_X80Y99_BO6;
  assign CLBLM_R_X53Y100_SLICE_X80Y100_C5 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLM_R_X53Y100_SLICE_X80Y100_C6 = CLBLM_R_X49Y107_SLICE_X75Y107_DQ;
  assign CLBLM_R_X53Y100_SLICE_X80Y100_CE = CLBLM_L_X60Y98_SLICE_X91Y98_DQ;
  assign CLBLM_R_X53Y100_SLICE_X80Y100_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X53Y100_SLICE_X80Y100_D1 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLM_R_X53Y100_SLICE_X80Y100_D2 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLM_R_X53Y100_SLICE_X80Y100_D3 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign CLBLM_R_X53Y100_SLICE_X80Y100_D4 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLM_R_X53Y100_SLICE_X80Y100_D5 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLM_R_X53Y100_SLICE_X80Y100_D6 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLM_R_X53Y100_SLICE_X80Y100_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign LIOB33_X0Y145_IOB_X0Y146_O = CLBLM_L_X50Y107_SLICE_X76Y107_BQ;
  assign LIOB33_X0Y145_IOB_X0Y145_O = CLBLM_L_X50Y106_SLICE_X76Y106_CQ;
  assign CLBLM_R_X53Y101_SLICE_X81Y101_A1 = CLBLM_R_X53Y101_SLICE_X81Y101_BO6;
  assign CLBLM_R_X53Y101_SLICE_X81Y101_A2 = CLBLL_L_X52Y101_SLICE_X79Y101_AO6;
  assign CLBLM_R_X53Y101_SLICE_X81Y101_A3 = CLBLM_R_X53Y101_SLICE_X80Y101_AO6;
  assign CLBLM_R_X53Y101_SLICE_X81Y101_A4 = CLBLM_R_X53Y100_SLICE_X81Y100_BO6;
  assign CLBLM_R_X53Y101_SLICE_X81Y101_A5 = CLBLL_L_X54Y100_SLICE_X82Y100_DO6;
  assign CLBLM_R_X53Y101_SLICE_X81Y101_A6 = CLBLM_R_X53Y101_SLICE_X81Y101_CO6;
  assign CLBLM_R_X53Y101_SLICE_X81Y101_B1 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLM_R_X53Y101_SLICE_X81Y101_B2 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLM_R_X53Y101_SLICE_X81Y101_B3 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLM_R_X53Y101_SLICE_X81Y101_B4 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign CLBLM_R_X53Y101_SLICE_X81Y101_B5 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLM_R_X53Y101_SLICE_X81Y101_B6 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLM_R_X53Y101_SLICE_X81Y101_C1 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLM_R_X53Y101_SLICE_X81Y101_C2 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLM_R_X53Y101_SLICE_X81Y101_C3 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLM_R_X53Y101_SLICE_X81Y101_C4 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLM_R_X53Y101_SLICE_X81Y101_C5 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign CLBLM_R_X53Y101_SLICE_X81Y101_C6 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLM_R_X53Y101_SLICE_X81Y101_CE = CLBLM_L_X60Y98_SLICE_X91Y98_DQ;
  assign CLBLM_R_X53Y101_SLICE_X81Y101_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X53Y101_SLICE_X81Y101_D1 = 1'b1;
  assign CLBLM_R_X53Y101_SLICE_X81Y101_D2 = 1'b1;
  assign CLBLM_R_X53Y101_SLICE_X81Y101_D3 = 1'b1;
  assign CLBLM_R_X53Y101_SLICE_X81Y101_D4 = 1'b1;
  assign CLBLM_R_X53Y101_SLICE_X81Y101_D5 = 1'b1;
  assign CLBLM_R_X53Y101_SLICE_X81Y101_D6 = 1'b1;
  assign CLBLM_R_X53Y101_SLICE_X81Y101_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X53Y101_SLICE_X80Y101_A1 = CLBLM_R_X49Y107_SLICE_X75Y107_DQ;
  assign CLBLM_R_X53Y101_SLICE_X80Y101_A2 = CLBLM_R_X53Y99_SLICE_X80Y99_BO6;
  assign CLBLM_R_X53Y101_SLICE_X80Y101_A3 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLM_R_X53Y101_SLICE_X80Y101_A4 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLM_R_X53Y101_SLICE_X80Y101_A5 = CLBLM_R_X53Y99_SLICE_X80Y99_AO6;
  assign CLBLM_R_X53Y101_SLICE_X80Y101_A6 = 1'b1;
  assign CLBLM_R_X53Y101_SLICE_X80Y101_B1 = CLBLM_R_X53Y100_SLICE_X80Y100_BO5;
  assign CLBLM_R_X53Y101_SLICE_X80Y101_B2 = CLBLM_R_X53Y101_SLICE_X80Y101_DO6;
  assign CLBLM_R_X53Y101_SLICE_X80Y101_B3 = CLBLM_R_X53Y101_SLICE_X80Y101_CO6;
  assign CLBLM_R_X53Y101_SLICE_X80Y101_B4 = CLBLM_R_X53Y102_SLICE_X80Y102_AO6;
  assign CLBLM_R_X53Y101_SLICE_X80Y101_B5 = CLBLL_R_X57Y102_SLICE_X86Y102_AO6;
  assign CLBLM_R_X53Y101_SLICE_X80Y101_B6 = CLBLM_R_X53Y101_SLICE_X80Y101_AO5;
  assign CLBLM_R_X53Y101_SLICE_X80Y101_C1 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLM_R_X53Y101_SLICE_X80Y101_C2 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLM_R_X53Y101_SLICE_X80Y101_C3 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLM_R_X53Y101_SLICE_X80Y101_C4 = CLBLM_R_X53Y100_SLICE_X81Y100_AO5;
  assign CLBLM_R_X53Y101_SLICE_X80Y101_C5 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign CLBLM_R_X53Y101_SLICE_X80Y101_C6 = CLBLL_L_X54Y101_SLICE_X82Y101_AO5;
  assign CLBLM_R_X53Y101_SLICE_X80Y101_CE = CLBLM_L_X60Y98_SLICE_X91Y98_DQ;
  assign CLBLM_R_X53Y101_SLICE_X80Y101_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X53Y101_SLICE_X80Y101_D1 = CLBLM_R_X49Y108_SLICE_X75Y108_AQ;
  assign CLBLM_R_X53Y101_SLICE_X80Y101_D2 = CLBLM_R_X49Y106_SLICE_X75Y106_BQ;
  assign CLBLM_R_X53Y101_SLICE_X80Y101_D3 = CLBLM_R_X49Y104_SLICE_X74Y104_BQ;
  assign CLBLM_R_X53Y101_SLICE_X80Y101_D4 = CLBLM_R_X49Y108_SLICE_X75Y108_CQ;
  assign CLBLM_R_X53Y101_SLICE_X80Y101_D5 = CLBLM_R_X49Y107_SLICE_X75Y107_BQ;
  assign CLBLM_R_X53Y101_SLICE_X80Y101_D6 = CLBLM_R_X49Y108_SLICE_X75Y108_BQ;
  assign CLBLM_R_X53Y101_SLICE_X80Y101_SR = CLBLL_L_X54Y109_SLICE_X82Y109_AO6;
  assign CLBLM_R_X59Y100_SLICE_X89Y100_B1 = CLBLM_L_X60Y98_SLICE_X91Y98_A5Q;
  assign CLBLM_R_X59Y100_SLICE_X89Y100_B2 = CLBLM_L_X60Y99_SLICE_X91Y99_AO5;
  assign CLBLM_R_X59Y100_SLICE_X89Y100_B3 = CLBLM_L_X50Y106_SLICE_X76Y106_CQ;
  assign CLBLL_L_X54Y105_SLICE_X82Y105_COUT = CLBLL_L_X54Y105_SLICE_X82Y105_D_CY;
  assign CLBLL_L_X54Y106_SLICE_X82Y106_COUT = CLBLL_L_X54Y106_SLICE_X82Y106_D_CY;
  assign CLBLL_L_X54Y107_SLICE_X82Y107_COUT = CLBLL_L_X54Y107_SLICE_X82Y107_D_CY;
  assign CLBLL_R_X57Y105_SLICE_X87Y105_COUT = CLBLL_R_X57Y105_SLICE_X87Y105_D_CY;
  assign CLBLL_R_X57Y106_SLICE_X86Y106_COUT = CLBLL_R_X57Y106_SLICE_X86Y106_D_CY;
  assign CLBLL_R_X57Y106_SLICE_X87Y106_COUT = CLBLL_R_X57Y106_SLICE_X87Y106_D_CY;
  assign CLBLL_R_X57Y107_SLICE_X86Y107_COUT = CLBLL_R_X57Y107_SLICE_X86Y107_D_CY;
  assign CLBLL_R_X57Y109_SLICE_X87Y109_COUT = CLBLL_R_X57Y109_SLICE_X87Y109_D_CY;
  assign CLBLL_R_X57Y110_SLICE_X87Y110_COUT = CLBLL_R_X57Y110_SLICE_X87Y110_D_CY;
  assign CLBLM_L_X50Y108_SLICE_X76Y108_COUT = CLBLM_L_X50Y108_SLICE_X76Y108_D_CY;
  assign CLBLM_L_X50Y108_SLICE_X77Y108_COUT = CLBLM_L_X50Y108_SLICE_X77Y108_D_CY;
  assign CLBLM_L_X50Y109_SLICE_X76Y109_COUT = CLBLM_L_X50Y109_SLICE_X76Y109_D_CY;
  assign CLBLM_L_X50Y109_SLICE_X77Y109_COUT = CLBLM_L_X50Y109_SLICE_X77Y109_D_CY;
  assign CLBLM_L_X56Y100_SLICE_X84Y100_COUT = CLBLM_L_X56Y100_SLICE_X84Y100_D_CY;
  assign CLBLM_L_X56Y101_SLICE_X84Y101_COUT = CLBLM_L_X56Y101_SLICE_X84Y101_D_CY;
  assign CLBLM_L_X56Y102_SLICE_X84Y102_COUT = CLBLM_L_X56Y102_SLICE_X84Y102_D_CY;
  assign CLBLM_L_X56Y103_SLICE_X84Y103_COUT = CLBLM_L_X56Y103_SLICE_X84Y103_D_CY;
  assign CLBLM_L_X60Y102_SLICE_X91Y102_COUT = CLBLM_L_X60Y102_SLICE_X91Y102_D_CY;
  assign CLBLM_L_X60Y103_SLICE_X91Y103_COUT = CLBLM_L_X60Y103_SLICE_X91Y103_D_CY;
  assign CLBLM_L_X60Y105_SLICE_X90Y105_COUT = CLBLM_L_X60Y105_SLICE_X90Y105_D_CY;
  assign CLBLM_L_X60Y105_SLICE_X91Y105_COUT = CLBLM_L_X60Y105_SLICE_X91Y105_D_CY;
  assign CLBLM_L_X60Y106_SLICE_X90Y106_COUT = CLBLM_L_X60Y106_SLICE_X90Y106_D_CY;
  assign CLBLM_L_X60Y106_SLICE_X91Y106_COUT = CLBLM_L_X60Y106_SLICE_X91Y106_D_CY;
  assign CLBLM_L_X60Y108_SLICE_X90Y108_COUT = CLBLM_L_X60Y108_SLICE_X90Y108_D_CY;
  assign CLBLM_L_X60Y109_SLICE_X90Y109_COUT = CLBLM_L_X60Y109_SLICE_X90Y109_D_CY;
  assign CLBLM_L_X64Y100_SLICE_X96Y100_COUT = CLBLM_L_X64Y100_SLICE_X96Y100_D_CY;
  assign CLBLM_L_X64Y100_SLICE_X97Y100_COUT = CLBLM_L_X64Y100_SLICE_X97Y100_D_CY;
  assign CLBLM_L_X64Y101_SLICE_X96Y101_COUT = CLBLM_L_X64Y101_SLICE_X96Y101_D_CY;
  assign CLBLM_L_X64Y101_SLICE_X97Y101_COUT = CLBLM_L_X64Y101_SLICE_X97Y101_D_CY;
  assign CLBLM_L_X64Y102_SLICE_X96Y102_COUT = CLBLM_L_X64Y102_SLICE_X96Y102_D_CY;
  assign CLBLM_L_X64Y102_SLICE_X97Y102_COUT = CLBLM_L_X64Y102_SLICE_X97Y102_D_CY;
  assign CLBLM_L_X64Y103_SLICE_X96Y103_COUT = CLBLM_L_X64Y103_SLICE_X96Y103_D_CY;
  assign CLBLM_L_X64Y103_SLICE_X97Y103_COUT = CLBLM_L_X64Y103_SLICE_X97Y103_D_CY;
  assign CLBLM_R_X49Y108_SLICE_X75Y108_COUT = CLBLM_R_X49Y108_SLICE_X75Y108_D_CY;
  assign CLBLM_R_X49Y109_SLICE_X75Y109_COUT = CLBLM_R_X49Y109_SLICE_X75Y109_D_CY;
  assign CLBLM_R_X53Y103_SLICE_X81Y103_COUT = CLBLM_R_X53Y103_SLICE_X81Y103_D_CY;
  assign CLBLM_R_X53Y104_SLICE_X81Y104_COUT = CLBLM_R_X53Y104_SLICE_X81Y104_D_CY;
  assign CLBLM_R_X53Y106_SLICE_X81Y106_COUT = CLBLM_R_X53Y106_SLICE_X81Y106_D_CY;
  assign CLBLM_R_X53Y107_SLICE_X81Y107_COUT = CLBLM_R_X53Y107_SLICE_X81Y107_D_CY;
  assign CLBLM_R_X59Y107_SLICE_X89Y107_COUT = CLBLM_R_X59Y107_SLICE_X89Y107_D_CY;
  assign CLBLM_R_X59Y108_SLICE_X88Y108_COUT = CLBLM_R_X59Y108_SLICE_X88Y108_D_CY;
  assign CLBLM_R_X59Y108_SLICE_X89Y108_COUT = CLBLM_R_X59Y108_SLICE_X89Y108_D_CY;
  assign CLBLM_R_X59Y109_SLICE_X88Y109_COUT = CLBLM_R_X59Y109_SLICE_X88Y109_D_CY;
  assign CLBLM_R_X63Y105_SLICE_X94Y105_COUT = CLBLM_R_X63Y105_SLICE_X94Y105_D_CY;
  assign CLBLM_R_X63Y105_SLICE_X95Y105_COUT = CLBLM_R_X63Y105_SLICE_X95Y105_D_CY;
  assign CLBLM_R_X63Y106_SLICE_X94Y106_COUT = CLBLM_R_X63Y106_SLICE_X94Y106_D_CY;
  assign CLBLM_R_X63Y106_SLICE_X95Y106_COUT = CLBLM_R_X63Y106_SLICE_X95Y106_D_CY;
  assign CLBLM_R_X63Y107_SLICE_X94Y107_COUT = CLBLM_R_X63Y107_SLICE_X94Y107_D_CY;
  assign CLBLM_R_X63Y107_SLICE_X95Y107_COUT = CLBLM_R_X63Y107_SLICE_X95Y107_D_CY;
  assign CLBLM_R_X63Y108_SLICE_X94Y108_COUT = CLBLM_R_X63Y108_SLICE_X94Y108_D_CY;
  assign CLBLM_R_X63Y108_SLICE_X95Y108_COUT = CLBLM_R_X63Y108_SLICE_X95Y108_D_CY;
  assign CLBLM_R_X65Y100_SLICE_X98Y100_COUT = CLBLM_R_X65Y100_SLICE_X98Y100_D_CY;
  assign CLBLM_R_X65Y101_SLICE_X98Y101_COUT = CLBLM_R_X65Y101_SLICE_X98Y101_D_CY;
  assign CLBLM_R_X65Y102_SLICE_X98Y102_COUT = CLBLM_R_X65Y102_SLICE_X98Y102_D_CY;
  assign CLBLM_R_X65Y103_SLICE_X98Y103_COUT = CLBLM_R_X65Y103_SLICE_X98Y103_D_CY;
endmodule
